`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mu2X/E3B3Kf8F5vFsnTtbtujLQRmtyrPcImCKeBWrhYNXnFcLX/1AfMtJfrV4+lp
WotXpeHBqrcaQ2lC+/jWdQeA8irZzHKMnJezVZ4K8AOwUpCX6P6m0I/+N0IYXnnM
2OjLbFoWkwt1EtOkxVgCYcgm9zlF9bjQfQtYsubf7ejuZuYkOdeOa4ZSBcmXIR5c
dQSHtGbrT+satSPtrui7EdyxDDyNnRefM7Ni49RSPp/Yr4PKg1a8OYR6Bzlo5oKP
XM9OijuNxIDD6F0i0fYG3TvM6/KAgH5UQ5UKe7W1YdNV3Z6wXyyRy9lsXhsKtGXy
mljmwDRHI0P0vnV3Ne/mM8MZvnJdDOG22Ga3qXkKW9XzuTBjPn7f+WqsDnS8AxUk
dSPM9VVJVvJErhYdYOGl8AK1lSlrCjMfhtnLnKRrT+rCU4wzgEuivpxcI6ThOnpV
yjX1R/YF157BaJbID11D7YW5Hrg6nkwbWJTPkJiVCH3lLTlJU5AILItGO37ryhs0
b8PKIziwFWd3aIN/NNKMX6z1aD1yvvYojC/89KeGwAFHg1b8gmRQpjnAqBz15LM3
NFB6TX63anPzSgvqKNqDjZSl4j1+hsTJtbjLj9Rqg1pNcq5YROtM6jnQ+IodrrB3
4d8+Nk8T4y3GNJwfsoLu2VfyypZXjgsaTsE2CaVg6tKiS1JvxWXktkto9F8tqAbL
8rye2bi9mym2w93S6zuRt+oQZdfvhBWCiZhnFzmr65T9sPbiyB5AIVS0kD5a5AvS
ir/epWs6S7oKIEQ3kNo5/sbslNEGMaiAn5VpTpkadSYalLlgAzpqYyHT9BzbuBvP
L6Zc/GxwMG+Z5KdRQjs1GA==
`protect END_PROTECTED
