`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z5e6vqzSUXA/UCceJeVdYu/+i5Iu+wqcujoToaoFh9Q5hwrNm/xO5Tqn7JxWw0X1
njmBCVoVVJLG/AbjQohOpDu+XFN99EO0F6n8ar64qOxr3sT1X3I9DH6oL/xKTHwu
XczOjP5DF8Mvd2H9KuxoTBvjaEFRpKIuhdTkQiOGGhQzAbpJfetzAUoOMzAMh4se
iAFY/qEqxmmLpkrwRwwmjimV2loIN5xd+H8g2RFGqItiArxUlmzgG/Xq0fJ8PYDB
D/fDhUMr0n6yPadkphEuD+N4E9y6fEOn9BCm5KIx9+82ohrPD4iY1WvPKuW/fhkE
QcNf8WcxJGXPuhj0GFgd9Ynv28J+ABMzuBtodEXqndPUf+hWj3uYe1f5fj6yHtcg
sjViKOjHvn+w2brTko8mx9bUXV9+JEQRx+pdQQVBvl/6Eg4A02DpLuwTiPUQmG+h
6aXhTbs3wRgCVw13BgxHgyRTjCbI1Qol0T8S9FSbZ+UOVPEDoxGvKqHl/0BFvga/
bFw3VWG/yKohSz9eL3voCg3GUqiQj9RyeCipqjKdoIsHSs96OdengQRe1AnlUH1I
aGFCrqxviMaciqHRN9f3dXRMeEntL7xOebl3Q8h9E8tu3ECbavDQYnjuC/CIx+U6
bCEGGS4kw5DosZZ52EYqIFYLy+uXBNk+8KA0fSV2beMxvhEb+nbMlgpGz0tXePlL
Ka2p3ZJzfz/jfaJpCRHDeX/pgcEdbP9ZvSnwmGUFdVYflywP80MuwZyn6M1LUoa7
fDKh0+KPPtc9R0btEBneHhfddAAUeWOla5Bs17Bb6d8KgskkLAB9qH8ipC44u0fL
/8gl4K2FKAHQjcaMvG6CEXCfo+wfoFOSX06j+/8MRdivv3Tr2A9Ni6su2ybHg9Lq
2HUYmB0zLanrXbXQ3m6bhiSUCFlKCsGdnCh/I7DrZJfNROKRJvX7d6Dr78hETvrI
dOuRZuqPlyfITnYo9jykL9sXpmzdWXIAK9dFnkOioEhBWCZSHJwriNXCy1gESTcn
ei552azM4qutvApbhWu/OUxq7v9p2gO7du26bpViHqy9B1m5JOWbfB3QETibjRRb
twZXaf7X7OJar5nIKkQ7n4/BLu3Uvte+uLD0oWl101OTNGDtAPWLhEBMRhuX7odT
PwycoFLaglZVZsgEqT6dVMKaZBGxpRTd1v6pmtWYAV4soJs7jGF2NV5iLE7gSZ3/
trcE+pDkCzpwuUK24jGJ+e6L34Mb8fuaOSFRkQq2oPTzD6mXffkVcjb9QiOfEEWt
xGqggIXPmhrS1ODD2DOkLf0WqsvsA7VkOySMS5LFfRuRVz77vKywJEFjqY3YFW+I
weSW5mU+Xf7n476Ic+A012d3sbdQw2rs/XKxfa/h1m2Gla31skZ8EYDffAYOqvn0
UpmF1zg8+7D2tYzTdNhJs2refCJImx9RR5QJjeIOqaPv8VjK6eutK7+vQgc5iFCn
bpKmqDRC/ELHFgfnn5RhmLpbxwf9qAr/jAv474eS73Aal/iBis1+dTQFjdfVlKzd
zaY691sm/NknEADj25EB1+FyDtwzP3ednooX98kXYh3QrfehQaAkLBLlVqmsxYBA
iKLM4h5wuepvmp3ANRpnzJdI/gHFv0r8TCryWiTS4mT7Mm9HQf/3hGobEnN8NkeX
eiputBxkWaQkoheSSGma+VkS/CIoHcRf0g6zGaFXjj6vOJiwQn7SsMU0BG1bFoWz
0tl2UipqJefZnfldp57pC6mN/Q15bxCeoBiCmULNHQXExhiHsuT+FWd5COkaoi3a
b7PiQ+uFby0x0lWXp/EAKa44zwM8/EVqFFtzSGeh8sydhrrrxz3S74XI93K12Ksa
4qVhymm1zBK1N2qGpu8X9NO4A1+gUOdultO+vPcWd4ztDJ841aniKtpI0XIcziu9
D9XsAZtMyqbSeIZnXv4hIAl5fPmp3pBJq8qM1LystyZq+eYHLFPrd9+z8Y3/HME1
IQ5hF7Mk36CUj9y/wRavghhd630X/MTiDn00I8oR3rXs1HsvJ1Q26/QxQNveOBbL
2syS3DogoG78AkNvSTR5RnAv0TQVAweyxWYAnxXNw/b1ENuQHUtIefpu2KQsu0Bu
Gp5jRHzuCrAgw4VVgQ1t1a+4imnagSlfhFSmw8fFObNv7YLUMzVGtjbSl/jjqiZc
9NW5oH6kilSWTlIaWsOlxQ5YvoXSP7Sb15o3iYy1ElKpF/JqLV6RTi8rkf9TmXLd
B2T5zbnu42b7mCbsE+NstvcXCfBnbeJ6NIcTN1LyViuw+moYijlFDVPkO5Ee41tJ
lJkBWRmEVDXgNkB4cdn2Quzz/M7p1Gk4NkaqfM1VQyIKfbCVLGCNzPDghxVXhTau
F5bKqBihEU407Ccs/NqMNy/N7TDW1MyauR8GjEnhiw3Lq20877uG1LGwVLQ79JFT
yUAl0+Z+ORt2s7uNkilyHfreiFpb2REKF04WWYX1FcOHJDvV2EqbVEzV8jpgwJEY
UZ40/nTqj4njhKHs5qUndObV7FTw6uBWu5j5urrQpIqWLFWe+F+S8EgQiZmMqr4R
XocMvIYPuq8drOqrmmOcg2fbE/rHmq8of0bNzvXpOedqGzpQQTaFLRs7rNNHWnd0
aYz5hbO3VZtuctwz6mNDVOiwdQ3ZvK/W0S+XADL7mjqbjkjgWUN9/WiMh0sI7QPO
27YdI6wvcM/y06h0nql/s5Ap9ckvMesW/poRX46vaGl1i01dPNS+y2rxMkz3TliG
MGmqKUuUEfABh7LI6VUPhp1wO/Dx0+oV3F3HS84YTU9YTm6ciGOMoCwOPyyRv8G5
8hw3pwFfElryk7PzZPb9w99USybk2cMbA3WXyk0PGwqXiSASZH6oxSV7eoohoRDl
IeU/BxqwoU6cQpsBwO/GQhTM6ocFC0Zk4ZL9kwKi6znNuvRArShZs1tb7WG39KjY
Ni5xIcXTXmcC3xCbHDAT2sY9h82/H0sKMtWsNol3oteLe6NBw84hEvuMuctTfUA+
ZYOLl1/sU8xEFnwFWXyTVA+LdKp64AMu+btZx8TbcmOhFs4uc9lMCoTqDVOFmKla
qANftb76i/gjOobwE8YyW+W9VxxgYLFy7kmSFNxo9rqzPdE5kiXIiG62V/Ewj96v
u8R//sCnu7WIPUWKUKaJsOpECJ2Ijly3Au4ET/e1O6hnk66UEln4vloZAu5XZKJc
Pa1J6R1Tj4TNBHem3cBkF8e0UmMIR0sjydlpcQn88gR3uqWg9QJVb4wNWcFZPFkj
RGPIlfTqrdVNA+y4tnNf44BH2S7u3tLvlXYicdqjwjOfUnmPAiwR3Zwekz8wiGMh
9r8ucK8r5emOPoYk/LIjvps9AitOXoAtqk1flR6DIXTWnQNeQ2TYBnzKzmYYacmx
+wt5UR+Cfq+pMGRR9j7RerIC7Z+vR47PjJavDxYlVNZayKkS9Iv8Em/G/qHSdw4r
hU0JFo0+4JI0tKwgJnNP+ZPM8ydj/nPPBl9F1bHjN37zbhvYZvCxyKeC/PumpRcW
yqcjSHoC5Fr5XWRSa2pnK7NH9iNpdk5Yf5KTUcNBPGPsdi9E9dyWTLXO+j6kbGaK
JCBD791elfc7Nzog+KfLt4xojIlNSapzz5diU3ES1gmt6X8KgcytMWrV+YveAl45
r/rSaFf9NNGp90Sf5o0EcORhO/1dyAwLjJxGBSY0GG/RJxiDP4UAc9TBjdjxE4sE
yT6vAuQ+2NA+sd8YA2e/sDO/Np8vSZw22f7oUJN5y2i6jCAhFU3TSc9TSY+7uhHF
iB1i6K7PmqIZNovhd/GgqsfGJZk6+CGIEZvrt7kmOylwrmDD+sLECdh5NryGEybn
4aL57umybUYTVeMWZeWmFuM8e40Cdimd4Tx11eWuwc/N1XZUkwyFPnG9W+YyRWgw
xMiHCxR/NOnEHmtRphTrRmClHmENo2WR3ri7cQV3FLvyn6DF9HE9fiTc/tuSkUeJ
gSJu/hLt8D3pXbnxhL606xIhDffbEiiCnRlB1gr1Hbn+M+eb4aJD+y+SQhzHXbA7
6vA3kv+QvGhRt9bnBHecieqMk3vR/maS+yqv0P/92OLTrfU48x67pM7EZHew6bIn
OXep+gfDTcYANXzWXzei7FjtOfa2LQC7kGrWs3EZQ+eV39JrrbABfKF5Sd8Ypw7Z
ez3Iqb5NZdk74FBvBETe6QZLyw4VZYK1L3bHNeITWvgh/4lBmxR8W+8SrOozyPQa
M2teuavlP4q2s8CmtvzTWA7g+ZzQGU+G6PL305Yh6KORnK0nfI7ze8MdHehMiO4R
HTxsIYwmXG6e+++708vXNyi2y7gc5RthQZg2cl5TiEzSDcHP43FsDRqsfMEu8rRJ
saTrn4gr+clV6tYC1l+nXSz8CiMSt0S+P3uQH94eDT2DeYuJnFeZrWB/XT549qoM
JWslMCJp5J1+R5+6mCbmtIECc1LczadpjDyLMqbzdItM8aQ6+dWzHeNfF8OPLa2Z
SXZ/YYrDn8jk7+71MfDIoBHDyrA4QAEAqsy+Ahza4wL3jXFy4Mi5wA/Y4TbouozA
Biu0gxohSIkor6v9tMDlNEbtiC19KvqTDXn8eIA/ZFCeStkSa+ecMBuuligC4JeS
Es8TmQy/edsBZAETO5/N7b5lck9uJjsQ1cmZM5Jhv+8xytfm9tjh6GmE5E3mhWWC
8VorUVf43TXY/p/p5oiFz4+mwqLft9a/XR+Mi0nIL4hEYiXyxMTRUQ3Wiiao3bk7
ho+r6G/sEIIwh5KMWgFfoHX8UnGou/hZRbQwmZMQktMzbWjW7poPbox4S+uAIhWP
460rhzSXsmBKG04IH2q8YKUdxAhij/dyeOfiJIfhwO3O13KI+7vz1u+56+x+HZoA
Hf925u45Q8c9MRIcbwQceEHQJY08ZJXJ0iHXV4qlUXQ3CwPKCJL7YP72rDSQCU+I
QqB/Pesju+eIX5VdYbenSW9JBqJ2GkXMn/9bMcAYqwCUSOCTs5gOcjiIl9RyObxh
HB8MFYkJRWcQdW2R89fKi4V5eUqvMheFCZEGKK0Q7unCUdHM1Vo48KnporVXaeeL
Z9FD9AVYYCcMQCIYjKM1y+ZIdC7Qk1LcUTYeVH2iTZz1ArNw4OGwZj48RauQi5CK
lKJhGL5A1H+HOqUBA9pVtl4fggGcp68Ghe8HuzMREW480RaCgYlF6o+Uq8OaH6Gb
MdnvwuVO0BIu6nsrqiZvvD8I7v5W1D4AVNdZrFjrrtIF0Yerv01bV+nIhiHHx4nj
ArhRrcYCYFBTHPP/uIeNxj87kCVvVyw6eC6BMO5tFgYjQ/kqHN7LxEZJLq+I2spA
cYjd5DVehEoGo5/JLa1IF9YhnEzRnlkmTjWFPrqB9mIYtKNTBlWFhNegl6EODyDX
2J7LA+od7U3dcq8egpcKPST6304kWgilYKL+IYNmopL8TQVhs+V5ra6PQQ1Zq9/J
ivyiD0xqvYxujz4zw6uH5hMhTCOourpXobtLgFPjY9ZOy9B+zOCD0hgqrhd6hSWM
wAN5lgBLS6W1Ejt0bFdfegIxUJO6rPVBJQGQ3lxVkO1aZ9GFKLEQm8ZwtrSbj4qy
Cv7y3jPLNdnc6bk20J5uBTWAF9vx/abezUyOvwWyi/79ErOKeXt/0H5A3xoMjFkb
wm3eUtxC8ooRbSLQ1BPCXIMaHaNEaly6WATjDZ1ZVMtOBDhlZ7eAUR40FijMQVmS
aGMfzNCwguAbfz5XUbvQjJHFAHMaMFD3jHM7ebBIImJ5cnCO1L5+NrL6gAdErIF9
dzXs/FgfD3xsx6UcZYGAFciq+V3OxlWJ+7RKZb2mN0NOD86ROypD+znbTVDdjA/k
kVF0CftccX61/tTsFeSSL85+1up9kocz2GlgLpM015GVcTPJGUBcrUB7/VqUUNY6
yxO/9x8QciIgy9Sh/jPvSLrMjgg9XIa5G98hVnrlgoxOXNQgihzyewmSAsMu2OcO
tpdnPNyYTDlfcseiVyyyBJVD8Z+4p1+bj8j8HuVn4MTrUAGmHvXdUNrZV88Cr+Ho
aOz1H7Fv4f67ncVqv1CBdJn+k7AuWwuw6eH0/nbFioC9mvVQfF6BmsqMsj4LIDQ1
It22ePmjVYCSBCvgC2ORU2telZ97UEq9gpODxemPEOOmnXw+VII7cAfsALqV8Otf
fUA66OgNe5PN8SHDF5mGXEdBW1FdMuIEhBXjYyhPosM2/rFcB85mnz5yBzuyIs7e
nuzc4RdJI75TUrKpNQ+9W+WgActjhhgODdkbCShJw5p1HAphSkFbLhC7g4Q3xdu4
Lwqbq7Yb32P2pUpxgDno+zbPuwcBiIR0jZW6RsQugpzbvHGQ0xfIXD7vXqPX/Ffz
GyzA7BV0g2mtLSx+nnRZf9O8j5gVOcFOrsCrc40/HepktCl0BtHoySLeCmj3nKvs
wWC9+csWmJJLTFgDZ2F3N86wnTguRDvkQVQ3U6C418tSE4gMp6LNax3zGAahz3ZG
8g/aVOGyDv3JRnR7WbiLFU7qxSGkqJGJYfHDJ+pJHqNqGeFNBdJ0Ie/SlV8s2krO
JHWXo7EesSoELZQC3n3f7pk5t3FPcJmwOQljlEX0Gk28av4sdZBMvhgEOsmr40KZ
2CEM8QTP1+M2wy7a9JHAPmoxNmy0UlNKFbrNEapGSIQg8q0NjGMNuUe9ewWYTnbd
cqrZwFoZuUMgJ0vA+8QVojUj4S3CPy3I4+OIApvOYOeT8BowehoblqIuBlFi3Oo/
8OEvcO1eAfcVL+SFL3f6+4ytiFsCcU6L0KLwRT1UURFIQR1J59j1RZ7eYCAKz0mT
NeoBsAIl6wqpbwPNUH8DfbZdNG4NQvoTVtGrfBnaMGr51NlL9zOv+0w/e3vUwMeZ
5F8/QSuafRpMl4f5D3q/I2dNclB19R7Ut5o75bNP0wb6931js+eeeLTWp+hzmY+I
wJgWiM/d4QTYS3FrwEMlZo9KZ/pWq2JtkWwp7f7TGiDYHlN/rBZK4ykB1u2wnAgE
WV3lenTay51f7RIJfLk1nj2JRDIN79DFkOJHqp+cXua3qtlS2Jc+IPlQ9Qc7Illv
pv7wiSrxn7+fTw+togy/cW1T88cbk/g8IMRxp5UH19A+97lvtfXWMr0ZKGjdBYvr
O19eRaYH+bhYl1bh/EoniU68Tob8M/uM0jg15XawAdbRMagPFbUW0RiLbF2TBqUp
OrGsK+HAQMpLJ6M+Jiu5kpR9Z76xaCg/FVZ03Rdi9Zx8jiLMZUuHHnL8qWF9UzJ4
teDYvHWEr1zNACOneK1KIffFbaETLUYP77VGrY6WpyhZjMfgujnVWViQYOXqnFaB
8qUvBGnvNzIW98qnK/51j7OO8kPtf74FNPD7BrA9IEHasD3vIkjox+gRa6RE+R1s
5XWPngVo1+/2arBKfGWxIu1EHYXZyeCfsRUrcisbg7MpWMU/5tbhsZLhWnsBLoK6
3pvJgYx4BJk6eDRsLo6lzeVDJjZO9LXJNcNb4e7AK4NF7pUl1eZ88+iW3t9qFTfD
JQaHnrQuonlQuL+VV4qVHyROxwuscptFhbTGFJgACwR/lpRnmtg+Rzz0/rG9UGxx
F5INsGVewn9NDB8trkKkHYkUHuFv5EvY7x07t8ENMxrSTD1sCMcfZc5TUve1mZ9N
Ac2z3ZoWL2PmV9PUqhJN67bLBSNBLEjnCBjn7ioxgAI5a6o/avXzKZ9/8+BnpW0I
7e4eUvDMKmD+c8qqvjsNKU5W9rVQTeUSnxipeetHxMUMtr1XshkRr9aUP+ugsjlH
k+CFQY1H9CBT1j8PvZG1NSGDgpMZ9c/BGXZ9GRqzdVsJBVrSYViwjxLJdJ7R2em3
WjJfGhf4t//azA962dBCoJnaxsNDrF9oP4JfQb6lMyWF/uDPybY+jrQn9um0Iyrx
YmoMboLAg5vHkwpF8siK0HHwC3IxIlHMUtMK1j9IZZFrk/6MX9XjJZMwjAm5kpHy
ffMwNft3yJl5bOUQlle/O8l1WFfPRggO421drjf8cRT/L0qw/AR6ln6qw/Htz9wg
l53pcX3x7NFQQY24zpJa4czV1h3PtjYNvnD+txBh90R1VLI2tQFNHtNukVCxGfFQ
nTqLqqKgdbcEg4YZXF5PCiSQOTsOcmCuPOZzxKdw1wCtGzkU71/A2smmYyAxoBEZ
TiReTl2QQPJQDO1pWsHN8Y4ah6MeIOBTFab5rI8hsy5D2khoTEmAS7hrD13jKBAq
TVWCMdD796Q2BtywI57XfcGYN/ZNKXQpaqjs1MvgzrONKIdXG21An878fd1KiqXa
65wgJ5HhWRuAyNSDpjSkdcQ8Pgs0tuND1iU4EpeL6MGIEnR0wNXCFRcNKLlhR6d3
FIpT4BwWWXtUBl94BXv7YAMyI4L5dK/Us60utZTAulBTllpcAH54u9ML+km3Glpf
R3nvNKM9ois53wCzpSuVM2jAWwEkWWhK3Cjr4GXBI3wcR3hO8I0MipHWzYjBDcx2
TZl8evHQUbKDUgtVJqQi/bdt7TMji06E5fvRQIE4+x+ggLGDKZopKfWE2TTaY9qz
k1M3hAnmaQfJ4B0F/oure0I7dhPLGZ5LeMsUjMM2R0P+39FPP3Cl1PNolcwTvleo
f3BSHhzAAqC4xQ+HvSx+gZUsaB3UGwUiEDL5vtLWeQ1ZXIxWPNezpUhWnX+36dhH
gDgXeeTjNLMSoIiY9sXH7tClFmqh0+sc33F057ZtjCXnaBbkGblP85Ayq7rXzKPZ
l6tP9aJhS9f3Vp9822SLaIlbPTCGW7aCbUiCTz9EUlxUFUuv/fBg46ShQ08jMszP
SeUYQGl+xggLRWRvhPATctSKUBjHO9uvQQYkeR30BSvKk8XFJVdsz/PQNiepTSVD
Wkrji70YyqMGkH5Rjg/2VtFRwyAP7u7EmcqCdXKPDtaFbFBZX3F22LqOXCv8UN/T
IilyLP26sRfiK4wNDoapCHxyFnoUSYTPS05Lb3qpPiET9+rntN1KyI2LvD/cqlP5
dGmkVa17sd31iQFCnGctERid5YSBWgj+5gCepxOeC7PRao5frGWrGv8zECcGmSQU
4ZkPxew/+Dvu0d48CCaV5MClGwtCXqTThdXLAgRf9H0q/eZZKDc5MDCo5sg0XsTN
Ertc4RCvSQrOV0WhrP5w7jSRV/wlZ8vtdEL0388ffUEkFp46cxcnQMY2rLzPPrH/
PzlAxqhBjz+wsBGuFnIiXRzDY6eh2w1SCJFgi38qLl61VkAkCpbfrR0XWKryRE8B
zao42bA1WT/JMev2rx8XJ9YKYjrugVINiaovlhbbK1sgwVBJ341kTfZD4E0Crypg
o6fqVZsDzxZywDVtgajnykVqReIVFng+2wTZDTVzKFgUx8uHAJVnl5gLFrhXisTO
Dbalz+Qq5N+7haCRcnBkjPFWr23xYTRnwJqtf9j5AU39xBSETX6KId3HYqch9aDY
GzyuYIirDBB/O2CBickIDTpAN5+5IW/pjcGKgXXZmlI0gXHnIOrhmQKnHTRuxWj2
D/RrQqkgfa7+oG8L/NLxz2ANhNh0ZFtBFH891Wtw0y429Zi3+NbpsjC70X7YKI3s
8m3sRpK8ZimwlUQcWltj9n4Yuc/vqJ6QFF3dItxQpPs2xtvxzBkMRYxj9jK97AQ3
KkZH1OGn3Rsq5V9d81AYmHqxxqRNVUx/giDV6CrSLaicY5ycUxb+qkaf/fDHvfX1
piTEn57TF5yHOfsLeLuv5hrmS1U/QOKm7V631jCLLmmRxqmk3rby46mX9lb99l4a
W5oi7ldHhQTGovAT92feHLXxmXFC/+75iP2uIIoAJ0uSf4BKgLWpkilPfyDWzDi5
4HfjFWJpp1agNu5UzMsbWUnTGns0NawgD4V552jGs1iYxdlPGFCZDQmGMIpQBApQ
ekIzM3Hv3Sv0aLOpmddHQKoeTSV9U8SmEzRUR5kTOTh9VoZ/9ZxDtwgXq2iT1zwZ
oindpzEQvV6DsLUEc6kQ+EkzlqStRWGDOE2NrhO34iCYDjEycW1zUrDV+tfUfjov
hVJX3+7uquOv5mxWA1/mVkIqstzARdHSKabg0bHHynPuS3KjiHIzTwcbRiErooV2
3zrhh2s3d8M4V83Gs3WzCf5gDvKsU3282QxXfRhe0YQkHkP7B0jOQLgyVYLPtxiR
RzzUn67d5+4RMwugboxQAXf4M7aXixdDemwJlRXSpjXRDegUo95CvClgR+L6anpt
tsaFwc9z7JvYWuLDSXQs2xjXJf+4Mc+RIwbCKTj4zfw7/BXNa+AZr1HC0kdypj1E
aDhaJXHaK6bt7ErRO/ddxpxwLETJAJt+s2lYYU5S3JYAshTKTzfsgLmLylus1vnB
O92dWy5BUkdicI5rdB0fusV+6KkBivudKG9352VcqQQBG8zsi0VETYJ+95mRqTjL
tpx4Kx4vWE6REMk5TNJ+b3AYKyNRXdHHRgCKEkA/sHOCH3tSTCIMI86CHPhZg2rA
96WJmG/fL4LGVVOjQcmSllMaTkZxzDjjhxmdRlrtt9kK15+HZSGE6Eag12Si5UIs
njzvG2C6/mqK0tt11MRs1H1ZVcySo0c5iSH+4EZMS18PD4IJixXdR40upLJAJGGp
EsstA4eiowwTGSrvJrcCYE9QJ+wVFW/i02UpOiOB2Ee5ZNgrpjazEsakqbCKCSJg
O/0+U0rOjYIbuVPjvxTusWVE1RIoQ+5QeIAOobmAIkx+0sw54uHBPB2imRqOuljR
iEfWqK2YkMD6wVNTMSL2k3UokyNttrBdqTctcvyEp5OPJmzSxtJQ+PHEWyQuyRGo
TuE3dR3diIeME1rwF+AjMr86Dn6T0slERJowxc5GUzkYwCFi5LL/EaRhTzgiiq5E
MgnDf8RvDEVBgofhKzsB5ADlrX/ApJvMX1GwWg312D0Rg6RyFr3bYPrZfWiss38F
wBncunyjfYCcDn1MUitnfnbuE4gIaTUJCq2kuf1gRXJJWn+Zfa/ixbSmkEq/m/4t
FEe6Tgtc6gwePmNL8yml5XdEnwjtWafkJ2OuZ6T0mV1QYWLOXi0aeg2CXFnphDvv
6NDYOdL1ELl8Uy1GFI1NAsuwTzFwL1bYj7YrvzvIXnqXeF0Ryyg0Aeg9PZ6ixCnG
gwwwboj9ZX4RbGQ/OKOX6MUpz5A32sJ04VlxDcRUxV6byEa7c6a0x+la1j0wfF7/
aAe+3RUQ76z/hrfmfLQ7lBcAPILvL+O4kgZHB3TULdDsnpGwCsR3NMY6Sry2oTVc
pgXBxR5zvNZL5hPfoNpaO40qy+uonyYzK/urUKXQbYjlQ8vfOpLdt9Buv3v5vFxg
v8+9C5elb/6nldBWDT8LUf520rWhPpZLCCprjn9P46UyEeokGYGnQ11zMMIvAM5H
Wvwy4OpWl48fws4oPUoJu0WhpFzkeRhdxrMXQWLDnkyDLCrfpWrnjwE9v2Iy6/9T
2YEq5FoYuAXM84P3toxXmAJ2hwNxFggok2a5YwACix82DL/OR0uSn0BIIW+xV+4B
y2V4Kx7lGWjBGg+v2FSmdYl0KHOCzFefTzdJTtSMFOn8aqH+OU1N/SYUbI7Spj5Y
AkamV7J7f/1+oqfCU3myK/rHD1cbteQaQamSW7+iUqI1xZtEwfFAu50FsTwWnEkO
XxCW/qEUHv8DFHIEYG9lZd9HFDe1KkHzM78CoSt362IrKPyXaNhgb1s8jCj5cGmg
W7eQW+iPTpgJxu8t21bPhbkqaDqBWW3TtB9dJA6iGBu2qMtS3V8rlDkIcIy2qCTl
3BHtaqCabJeUlawGM0WY2pHd+U/XIRu8xe+kXF5HkDw+l+OJZ7ib3gcatNuzHNpt
PCI5mE6Mh6F6ZgXqyBNMPKorFHCVLb9ss6fK4sC+if73gfh4M/TbDSd3PSeVMm3f
Bsj9SiY12QzRBjLcXg074usBT9uEJxxs2G+KrjdFeh3jxbitFAt/FwG2YCPln1FQ
woS+reOMf7AWIGDuDY2S3H6XGW4o8KteN4UBsYsDxL1W8YQyX/3+/wA6pYxIajVB
vzN1btDfUXCBa+U1avsueTXwbP+sCEEGEJJnfPbv+FDzcRcn1c89Leuzc6Mn1RRW
vzoHcM17by/rg+SoeqKuljGm1OfreqWLureScVQ2Fj0Visx3Y49pXangpvKea0YE
TAejywP01/TSzzwlTebYd0Ak2E1uaFvPuCTi6Y6CYJ7rHdsmfSiBmy6VDbLfL96A
4ubIWXj+3d4hpFSvBAro+NgP0CCLVC2GQkWEaE7nwqAMnOffi6QKsUPC8uWNRe/f
vI7IeM+iS2KUHIyzq+0DPJqht/XesRg+PqhMBeUXv72X56N2kYm3NwFDeL0CgGDv
oy+DYrMPfhn0tiyAyZL3XWJ47RhN3DeWUxOxs8peXaHGkz8PeyIbR+iYJlK3R0Vh
cMaE/YapvT+tLxz0Ysh6RRdBkM7DctQVK/ARnD+l8EGB4iZCL5C8Ms6T7Im+5HRn
rTh5UHuZCCSBC2m6ypJeSKS3Ws1yX53/uBmhS9NAGWyu1THBMOLcGSNmWZoyAekg
HNlEnGiguSkEchFhp33ECq4jT7OCtVqk3RCxcalr3o8+pfLEHL0I6EelpZ3no4R/
ZLMHXN2QpiW1kX0e6EYn1OglohMWEPLGLNBrL6IVz97srrb1+yLvtd0T41YZzAeu
knPLhwc9QDG43Qyxdjj2UeZhVIvjRNIC9OxoLrJxz2XBqsumtgrOChUZj41VrU/5
gffszu4o71hOKfCIzOrdEEj/As3Ufk8qkFPNNu0M8JKXqr0BYA1HEnJ44G6/TGqV
krUP21NAaj5dNXD4UqMhC4kqwGq78Xuryo4sJ9arjeNQSuWdMfObd4A5MwyOPI9J
NpUuMmVYF0Uz8tVTKPMk6kVrZ6rpyu8kONftf4Wql1fcBkAyyxs507APubTgWRke
AtjTepgTzC4zyD6VYOuWdAwe/A+wOOE8ccPdNKHwXeqP7VBjVrBX5k2efj8rCwtu
BBToYIU1gKIJ12MvwelhR0JNsbs6Jz24SxhBZ8OoPFyBs2bRWnabMVTJ5ifdu9Lj
JszXFbuU15k6bgVBlByDMsG9dATEgsXpGq1nf8+9ZFdYmTXzSl8e6v1RMJPle9WC
jrfZTriLI1HtgxcyBQZR7uEwUP3E9asOgQeLvm8YrcyCY2pY2SXIG3kc8rb3IglU
Q3sxdGT0723/QOCqedSLMaAwdDB0P5pYKU3Fmy4NNn5XdqZ1Vm0PttNQDt74eVLE
PyLP71WWGdbbyBogqPpb87EtpqCMorcDY9d/Fk8V92ZpgCBLtOe5T2ZPMBxunVfn
mlOjYtb5hGlOH4qk6NEvPHGUj/D3YEtmcURJ37U0LH0EwVA5fkVEo5IitOMjsnd+
e3XnUamroEhX5fVZ9fndnDrQZHD0Lu54m+h+2ZeGjjag6G4KEI9ct1QRWdwuVUTE
q5wOlmG/Gid17+cJf8IYGVBxIagcyKCKYHSdmKexTTrNfAJ6Wpm5y9mPdrFDTFUV
1aAHoanyRokJRgeOZ9XiwZ08g0LaIB2E06yze5EU9f5jOcfp+iURO9gkFggA0UpS
zAno4/Y3pbAHQ6Rmua51t+WvA5Gx2Nplbg/2Q6PmLlU3dwK18Iy5DfvgNXyh1dX6
tQ/24dNXm2qG9Xo0+BKVZPHyzrG77oHaixMvTqkC7NRYUcLtULxvFDOAtR+eLcfT
zV6cCneP/+b/s2qfqNio4Q3y0UXASmzjm2fK0s8Hn4Ke/SE97bcz5ZrlfIRyBaPQ
yh85rCPPiPVAaJfHmG4ofi56pdGGAds/Ru/Qwxv01BRI5vIO6hlKX6savL5GMOXM
mJER0ZCXWoKUJCPr9SE3IxnPVgEeUBLaDSGQtM5K+6Zr3su01aVeVQZjW67x3tNT
rF7TsGEy62PRgiOym7SMrHz18iqLhazkHmEXroOPhE5ns1ighz8X5QgOkkCK58F5
elBaYMoGmEVQabgf+9kFdl6vOEqWarE7cT8Ev0oEKrnWXcGbUJVMFJSnyRdW6NRn
tAM6D8lXml3ro7ge19UHgrR69EZh+6Ug0mn2V9vYULjKsNsGWOEVlfcsoRAfzoB2
NBTpfGUVkW6oLDnbtZkPovUMXJhKAgoIt/TtzDKlt9f3s1IarxuUTu8Z09aMYNPo
4TOjYtCQMCLHpgj1ma0xxMDNQ54dWbFvsFoTwRDqnUIxb0FdnGUVBTcoOqAQhwWy
xSt1+jtA5E55UAREEx4lO043/Npf9rtgyV+g/HE3FKKka95BDIuA1K8a90/jOWh1
OtUDsH7cxCFb8ir+/Zx42BAKsMf/MuWFgaKjBKGOXLlEEcTggXzwbWRl5fNEG6tg
BDZotccvQ+74SPaVWQS1zcMvSnGBSamO0MU39t0DUsqkK45+lxomgpeLBnzHlPzS
QpZ+y4gRyKXBXrNBw+wKyA/fnV31ezpewG4yHYyz4Lxc6j4w6c6KSBfbEeYNngsY
re0ECWh8YC6QdeDLos7cEB84mTYFOPF4GM8iHmEMOKPGxDPRL0/ZEH2B10ldAp30
668ZVWPBNzH+sNyFPB/DP6jN5yDjIiHPcTbE8ORzk/9WS98TgdU2F5O1crGUKadc
rT8tGPJLN2c+FkiqNnLKlNqV9fPUSWJcpS9wiA+MJiB5aeA8sYrmUXjwBxGs4Ufk
b2ZRzHS6q3+ollSMy6iOyXiQzK/DI2UReUZow5OOCkxMEbCoyQNMDGS+yWLcXKyD
vjOx0A8eTgCS73ELL+M/iwHxOnOqiLJre084ACb2cgMRLUOv8ROK9ibjhy3j/ele
MQrFLiTdK/oZs3HV3W79miIpmkJ26RFv5e1bbcxebqOXAhsN/UtjXSa1iTKtC/Td
TVT65UrpyVVjK/CrtMUXbYgo9bCDp0cbPIR84ueUZ86bUVQVTJQlL3NSFLvaj3Ys
yZbyCjZ2q520GCnAg8nae8PFhVZXbogi+Be99d9cZNqoD8IigGxpEE+2LCu7jhiU
zbaJUUK3zkR3y+hv7jWHGh1h+isqiL07cgTxaIh3GecTp7Mwlh3ZEBsCQpdQ5E+9
uDXttvfhy385e8OsPbAIqwSZ0VZonYz3nVgJTP6P+m4IzlZ19bJd83AZ6IeFlHXI
HRRfjywfP8DnZZSy+R+0gJTOxBj2tJ21jhcBmyuSo5ZLgH4GiWE53EQ06DHIMmRs
uRIncOgGtwnb54PDdmf/2pIUkYbCYqYY7q6Fb1t87Gp+DwIWYPqk5o4Ye+0dxOzB
J0pM7KkDVCQZsxn+4V4wcYbsTaeGQMyGofUCiMc4yJJMwPRA26Je9FDDGjbgdB1w
cZTNsNosvwoVUoxc3piVALwsPCeciyx0s89rv64tutxrCOwgZRHikceUL/nGRJ7j
QlQ6uAkiALE/43gaSD1Au04K2KBHmZOm2ne7xRPNOMuZFoPxqN2s/iXFTqMfLiK6
qZVxW2S7wmtKKA8k5/C9T6KPowF2VfL5VfJEYksKeNXBYz6AElvHFL0NREAtvry+
10wjQ32QZizinO3LGUTLJNxdKA35/dqSIXyF++CVBliG3+BbJ6VS5FmZIK9XRNOv
9TxZrGfBDiAQ0lVQHEIg5q+ATQY6RXZf7rqI/sGVD7zf680482qmN416gVSZI1kQ
AEqfGZTweB6d63NY+98Bfrnd9E3ovUPIK3aEzJo5ZzPqazwwbCidtGMjNKsvYjY+
Cph/5hzLbZbYum04aR41eyVP7vyAs84BWd/9/DeGf+y9bgzVcDSOybWjy9GYT6o+
CTjf5alnuZp85F/Y8hJC/2wbaqpYNhAldnbt1h6cxxOWEIh1Zim6mtzF36hzFo6V
ujG7kpAbdecoHwuTjN4TWjDfCaH01kOYt1PPZfm6vWJRxo7KAhSlaaCC6C/Zx6/2
sIjfzSreiuEXY8tBtvEndD9fTweW2fZsBYaZ/X/S6CMY9mP6iDjaB2tGcyYB+BMv
eQY7/xB5S8qaRc9uj0fS8NVug0MLqlJ1dpoGOU7LGC1C8NjMTHNgtC2+e7+rRGlh
fU33HxN195DcQKJkTAcPAKjQcY2z5Ze1aINP82RG9h3/lQOYafsxvqrLsMkqnoQr
TBr3EOszdsAvnvBHE1NexlgBcNOIgvb+ADxWRT0W7RW5V7UQ/7gEbYIgSzo5s1kx
SgMHmXhftHaP0rLQPwzDEnxc5ubv5bpBBIiHxpgX0F5bpTnqh74CNzcjRLBFOtgQ
6JZjwo7d/LlPvYXCOkSYrC8WKGhEryaeR+y8IEjCdpZpjwEEDhbakFYfBJuOyFwY
HiWPT5l/SvCedVFsF2L4hpfD9LRDbGOYzTebmsxiSHSlqZ7wPjCVTujlVbmaUUBd
/guEBbfqOLPy2x/qdTp8wxy3eH66uBtDvYWm3eHbO3rxLAuZ8e/XCPk+FWTxyZe/
s2SNvPIb+YwMaWPnyFUs7ysenq7atcUrra44PLJlv0AJWLkM4eaZj7vjaxKVtYO7
pTMVckc55uxw3Lzm+qS2ZLhT93ig53mVi0ZaZ9ryKELVfDWhQYmj7UCzOX+WSaOP
c4NholYn6Xcd8X3miXa2OFz0Dh4+qHvLgarFPcL+MxMu1sCNNc09+YBk7FUANemr
/CfaYfMW9TWz9cxhU2tUMDmoG87/Hp3VJiBC+9dQBjeYfn+Hvf+9+DrMKmvEqbQd
Q6ikyb1Rd8ZgPWqg4c3oeanMjTMADJ/3F8pd/JsooUG+EBVjHUrZC2t8K4ZxT5yy
zXjUKRVkJ+sHIGTJyGXQOFzZa4zE8ANWZ/tZald2p2wBq9iaTdmndUn5oBp/dz8k
tcFTKFeUf0x2D/k+wwoIm8XyZfa/8vA/yAwqWnVJUw7Cdhdd9295xA1828p1SzK+
X5vzg93zvLWBv4MmA+vTVJwKRoc0YhAbghdyzHl1TfMHqkw+jnoCY5djq5VmAolP
mjo9YFzxgPUWI1YwEnFB05QEF0w5q2aPgAJqfM/Kxpa/wu9/vZvZ4MXpHXApu9kw
4Rh1oGma61YgonAYKJgYmOU1+ggR1UGKPPEUnunassPr2BJCNHHPeimHQ6THFjyj
QlIJei5r5LV//ylYKMtGkIDVkmfiWLKiXiJ80xUaDJ+33puvFoc2DTa0ca0wsgM+
5n/X62QAPDZxtJBYlnmrv8KzNlSpxSfWqJr8SsNh3v3rXvDwcJnVbnrJhujdCswl
H2R10nelT+XjJ0f/+y8fA9kqGhxr9p+ngEg7W1ii+z+6QAkZ/BzypZa0pp2rcjF1
OB0BtnRZ2gs/rGX4AxuaAj5a17BR9xYU8CVIgV+ELKsiin9pdYvIGVS1PisgEoBx
tJjUPUptMhufCHj2cwNvw3/g12Z73PvFvuU2pOUcOgzp4EvdZ5WaZD1M06wG+IwD
cByl/309UoElRIoSIfZXi/YpZfPl0SY2PA1sspktAIXMFk/EFYAfvRcL4blFcS5D
B8lII7t7lj44HlJliwLHpJhQiFP2SGHFoOMLZnt8rCtQjlggBUOCJYDVDXdlHaJv
7WqVVtBgGW0rwfH6lcGg3ICrLZlcUMNPCHSGuq3gb2pTyuCt23ye0jhS33jVH55l
PDP6/YdHFrg6fjp4whXvwRXU0wgl1Jb6RlgnNIekwHvAzUP3SV3lZMZQJgRmn7uk
4V81xMY9cdX0xHYdYn1XxscLr6V9s+uN5chEvHXP62acOIB5N7lz/ikC8aBocoaL
k/q+7iGCs0vbxe0gytlfDV89o7bGQROq9I++MTOb8h7OY7VVOzqf4hwok2Dtly5W
QOekQvAVL+7OuZk87XlkcoIYALECavTCOaHM4EXd25LydDSQSv9t0/V89lQyeSG0
oGElmWsFT1GSFBLPF7cxTfaf6loA+ZFN5prQaAHUzbuBjKpvRwjrX48BckVOBSA9
Bzt7ILMH3RmJKiUCgUULi00+CR1s2dyOnXSTWNOHtj69gi8VwYXzYfvejIyWZfDx
H3Ac3ZBndTM5AkBDycXbt9ag331skRoVidgwjfNyZkx28yjt1Hse4GpEg2EP2lXR
CD3c/HLsvHiswNNMx5ydIUZQ4SsatCRaYaec4L0Th18pACYHjQHdwMxD7cOUUZzo
A/GgHS6yThTsMBbOnpGUdmh6TJVI4dMedLuBABQaNkp4273CFQmM4q/Jtl1r0WR7
gaqIcS9GA/pt9vE/WY+OkLQzPHMVuVZH547YJUQc2gR0MMv9mM4M2uZGtl6DSDLy
LbP74ZT1CmMXUtM7VEkgN86+eUC6tCiB0M/JbWP1lVoVhsxJWIIar/9aNILNo+0/
frbSUyOJPh4R/llhMtRl2gCtcazjG4OyGRH/Tp1lha777o5rhJKDnYqv2mYqSdNu
zVz4Rk/UaTE6ZVdHRONUmNU3WeCinUMb6eyxe0ouVVIK53qciiiSfweklL1j4WNu
+T4shoYZGbDklXNZN8HYpQsh8CRnN4C3QOjPrS/o5fxlbbHfgsn32fPZLDb8DCmV
J2cByDM6mjZW0QUSyfS3LcJcPxzB0j0yHyZPSr4hxPXohEV0wi6qDBcDONx+euxn
1Q0VZlISNQyI9JKkZfe/xuGREQjhdSQakPtVIYPM2yndsK19DCn5Ifw71rJX+NF0
gRr2cRLtQDq+rFvwFp55mWYjyATx72gTluA2R1SGaAjLDcL6v9iHS8vz4Yh6wT7V
IaFI9WnMwOuHEtU3hYu6yTlQ2jCnZo+/cpKhbXLlb2uEpv9c8rzOS2YTfVoAhOjr
zuIR9WYEBCvhc0gsJU+ItZV+XpzJpoHRXyX9FVAer+BZGZbAZJaKE104KZZiTTTC
ZBouwP08896AT5Yr/zOT22xuG9a9JhJT0h3kT1MTXeuwU2+cI2kRSKrnpaXdg52o
4ojegVAfGCJQHDcFnkMNMkcpqYqDGulpK+C3kijA+sp2H8dVyMN0CfdLTvNC9ONn
DdCmvBUNfEkB1mzUoaLhbDkwAu9Ml5DaAViK8zILXBVHbnkdm10k/ZEfANwd9atI
IaBx4V/zISD20i9boX2/qOrBlHBzeYizxo+/pjiU27k9hG0c/Zz1hX3MUTIFdpaR
PqEkdwZ1y8NqoNOKKXSWSDZdfXoYeR0DtrDAZXMEyMGBeS4xYj0GzJiJ625a4oXo
3uTg59RLot7FV8rZ1PLtP9EidXp0EiZDIQgdh+8eqD06U/y9b4BD9T5WoqUoYMWR
ZSuxJ2HYJ4Xgikxott2TpfBgdJnNwkRyNNr5fIBHm/+vAfZEJhiU4PaZXXeKL+Nn
Nin7VKeisEVUBkH+Qc2SBL3EpgfXSAkZUBMXHSZijCxFPAwu8JBgNWruiLBtl8/G
trNtOsEOpaxuDuQQlFGPI2+OobYVdEWd6TtkV0O5gp2zXwFK6MnD2ljCy8H5hfzS
ggo4Kp2YvtrlW3/0d+rtZqRzt+/fwVxhi09OVznMvTuRNV08cVu9AokG1MdcHJIp
yl4f5Bpt88nomky8Mh0pU1+oAX6guxai2Qp+8FfkpXPbdRU9dw3tw/nQYz3NpJdm
V46+iyBDPe72i7r5C28N5y59o+PsJwytCpz0MNNO3IzbWcxyvbOBxetlIxM7+mbO
i8q5wIQ7BWMFOlwaDb6thYy0XvHGKf/yaIa0QHVpGi4NnIbvFhc1yy0MKuf07SWJ
gnm66S/248dYg/xYqfib+9oJy07KcgVbYs0K4PYtqO20+LPFLQXMzByKJ6/eLx8u
5VnJstknr4BInyjs+ETzA7GuRstl/7pCxXAQRsssNjSCmGPSiCAejI2qNlSlyc8K
HqS0U3RQ1Rz4J/4Fe6TrWLsH5x9Xx6aq/n2M9Ls2vkRZdsp2TzK1YYTZieSs7I55
sA7KP08uq2Wy98kTB9svPBLwLR2vZx9OMR1s1zzCBRmXvMHw2cmqS+f1oo2qdKuW
tahyKjGRf7TtCVrCSGl0CD5fe0EJzPd9PawP3LrbwH5ibsUVFxhNBAS3wsLbuIA5
59/JdGyRfFdk0fUqjWV41d9OHAuFPbOf05miTl9NwgY2XxFXNh0APClMza+PqoDq
z8RyyDEEIsKuvsxD1ilogpX3/omkHoQUsN8MiLBjhzgbdCJ6cuMLiBaoE9/ueDvh
jqqD1r5kct+YTx4ekTxhJY8EothHeTGoRif1zUGYoJYiCAApmZhFqxCl2Fs0I36b
QPZs+g9ycf7ZOZ0KuPOdVW+jL1NRVv6h8PUL2F9qREvUSUhEG/yTIZ8RlC4+WZDQ
8N7EmmYZ90EyDu4zGwOhX/OGpjkAZTrMzY/HPCF3aZWoKYt05+Si8n4BrHvd0PGM
NV65l+X4WAv4RvxMqJYVLXtz1+1a1IwLPkfZEQC4dsRyxL4ZSYuQG5zvbsQef1MP
T186WeAXgUJbii7x5MnD106ztWLtl/Tdgpwl8xETFY9cIJM5iUPju8ykL2cunRvD
2ryo407lWFSB0aa/qVzHfDmH+1Fuj+axBYg364bLZhLx87cltEvG79AXpmYL3Mp3
E49MVJoL3EfB1sMRXvvds1UhdPJAhmwC4kVWjVNubPRmZwK787BvlZiFym6ZHNcH
PHfmOh057Mccl18unhy4g4pyQYTJcJo8k0Akg+c5fBQu9SwmA9V2FCM34YfrsW1S
VAiua96nn631+QSJoMpFwGC0NdYwZv1sjmWGgddLtpbCbYdlISyObeIhKDXX4wsp
Qx4DcgtKqvD5cSdzj3NXUNEvfadP/KD1Lm/cUm2KaimmIuGox66p+5SPdbbZ0irD
3OVpp+XP17Dpe28BXXE5bP5zcAXivWKE4l9MKyW84cQMbS7zj+A9aunsR8Tl0Cfb
gl7M3uOUmXNAsDpP9hWX8EC1xZRFqOsoEqkHL+pw/GCXeikeQZNo8begKnXOetMp
/SghTwML8Vv22+oUQDJ4n24PQAVE/HAuqP6HtjNrx/sbS6RE8kntwrSebi5EbEhr
fUQux2kLKma4tFZCMucPQ7UhydcrLqs9mdMLPrYOApf8Tu9t0mIOO0GDVhneGzfg
6d5AofVAn9F/1oNnAztIJmowWmwG8Iy4kek/eZbvA4XcdFe6wkzZxA49jdNpr8at
su6JrquFbsg92jslt9l0WFTVdmRa3wB+PhhsYIBxyhYBZkSVM7pR91fTv5htgat3
Yv2xvWL0Pr1ozj0Y4yU0x4w3l65YIeJm5L7Uaw8Mfw/4X8CuKACJs3CutN41wS8y
XAde4i8KITukQM4ZhBYpoq/gK+G87SfLn8RKCTUpzJZnaIwIknGavisW9QbPRFv0
8JvmBm+LqixWJTGeR3httx4eToBXu+f7kHQZCdoylPXq67UxMv3157ZMTk3SFdDz
A3c7iOg1dKzc7DGqhFsaOEkujTDwiEQZfrZMyj1JhefNfJVyt5vpU3kBa5whzPN3
CqCwUq30b2v/SUubjVENQPvr+1Hs0Jaxpcw+EDzH3Zk8rNQzCbJFcrWAaRFstVm/
YDGvKW3vx9bB60wTLBj1apZCxpvtgE1T7/ksi73/93NVW74tdaJqJgkvpAXp+SNE
jQk52znSOLjGpOTWf4kATaLoa4dYhL7WyScDd8UKc0E8aJ6qpnXzr79iuWVG7xF2
1ngPiMFlXyqhmW+h1nuNd7JD7fRgbhi8rQ1EtfHZKmzGy1sOM/SVpD/uLtZxWfzL
CS7kl1dboiAPAjxk5JXQQ2LZxwKRI7m9YB1bZCz8q2oX9qw5Ek02amowfy4PTURw
HQwBQavukKf91dcdzPbQnWnpScckVu2TSOQjWeXP7gTviDAZ0wFqCrU4jEepC0jK
GoPDQFfyeiqJTaZFOJkD7+4vXGsWvj6O2x/Ty3ozO896fmXnpDllH34SszM20Bql
r0UUp1FcADdVud1UIpdItPcKGo79ekQu3GZRzt4SzTMnf/0D/fFdqrGiCkP2qkWU
cPwDTiF8mcYzkKY64FvnYyS5pXgZ7+UuC+RaHtKg7It7FP3vMKF3etoD/JDm3kyy
Ivy+XlQHlYVj1B2CYhDa0Uf8NZbBm4rBIrQINRHNxkWcaG0Ru4uePtgsyyL66j75
OkQpwnBC84h5IiYxWMHaEWbv13CSDKeztrDVjr4g5NvkZT9SEaFEZLUGNdAh2QQ5
6juuBOE/1ckEpu/2NZM6BLU73nkH8J/zR6omUfDyCpTTkkAbtmr/o84lX6aY3FcU
Xulu55KGBg1yEms2szDxZrXCt4ts3BfWQZqrp/v+LdiRAVPJLg0dydZZTiF1oH1+
Kpkv/KL9RFwpK9RN0fgS8g9RuNCp1MH9VuR7RWumLxnBi7GrufTkXXFNLLPGxg6J
XvxBbEgdw4g9Iw5gOgkpz4jBuoehKIwfef/3S6ZinAnQHGn27fi+TgzyHY6oSp3M
ukkSR6eZB+wOttpZwN95tU9g23hyZELHtUZVB4kJz0a3NX/pdEAmEKid5m3mGu/b
9rNVz9oaP9z2XfjT46et5OctdJsoCaIaQJqvvRXGCIOU5z5kpBmakLoVolt13D9h
XOP0mTQtjTrdwRVqNHeZZIb7y9v6qP0eGyzPS+zuD8O4sZsP709bZ3RDpLYMH+/S
VooEuThW5XZ5g65oesiaAJrzcDWqKTaJKUIybSTr6XZchCYxbHSWAtLCZgNt6YXb
6cYI2QrFlmy7OQa+/mCk/QGwJMiN+Y6vkoy9aVB+CHFVsdekLzqw25/UcoKnwf7x
ciC0gXOhUarJiztJxE/bim1WY5L2t5EfVX/EioMiMfvsyHcrPk0e0RjPmNB42iSn
IujJbwCiWALZ/8FtMXBciY71Cnu5fwE7XxecTc1QgrZBbGXPsJVyxci6JAaTz0/4
bP6G8Yo1gxAyV4xqFxRFx9fX26A4bdw9HrL9oABoM1TmkYo/3sjODj68IQZdgjGr
vEX81LWDW527xHejHZDMt0KXUUzPBEuXXTtrFdkteLqRuboJWyZx0z+W0NDjGbiF
IXccVw6Aq/uWxByeRrVs1GzaPtq6hgVOj6Puf9KzA5H5vRtYGtQBOxRuN/TiMIVT
Z/Q/H0out9dk8wLO0BgaMytaYZq/HJLuyXC8Z074fqm7d+jxJv06KbjbgO3Cu7zm
3nIzF+uobjcoG+phNJPvlI8SpbDXFFRB7TAeuvWV67T5APqnzEA0Eo6k8OL9AnZO
p6c+3mASzTBywg6fwJl9C70/hJVjlkZ9DP/GItFOnvB78VG+B7YwuQwsUoaFUG/o
rHwyMu1bPF7egoFZdVhjB73XkhKH258TnSRR4pQNBrB9R9nTk5goIbsXAjODi03q
KKcuKfDbBa6jiesXmpAdzdO8Dn34eAZbwuIx2f9LRGhDooK+WztcZyTNQpk7GH1M
Vz4d8kLsqL0pxgMtk0OfhtQHlPpR/HucARmDHVsIy4ozjkwuu6KoJtJHPxaFCgzb
9kjE3fjf0vYGC0U7IiwEiBZUuo3T+H14tkQHbnPPFpKm+GYpSH3IRCuGRTpw/emy
hLV42MmVxJho81iaBU7k5jZPIdQlozXe0WDs2LwIYa6MGEYZa8viBisU1gDwmevZ
yyKLzUtYyyvtIyNxbiiBhGow1ndNkUf00ZbVArgFk4OGRNsaiBXFFzIjHvZuZuTI
c21GjJ9DDvQG3MyYnaWhrV3ENWN/kqVjFGfwLDpwG0wpnsEB45shJVETXYZFnbUG
4eW+W+sBSN6DoUU4bN562lz64LcWS/RAcJ9u88KFvaHgw35xqdOIvpf9CPqcYz6x
GJbZgmgnwOLXUayA7PkF8jY1TOU07ZLGHRKoIqBq+Cks6AEA3KMnqnTDidhHJjbz
AivwJuq4ndKwYZxGsZ+3uvtVFa3n7bVm9iPcx0t7MQZPM2IXEDQZuZG0+ktMfQh1
V6wSZyF0bDIqn+RhOCse3/ueh1LCOfD9yOaolRnAGluU98tFfnFdAn3dgr8E5/Ma
PrXOfjpMLVQh4WdDgxvu9xQvBo2gf64UQ323kjfRUtnbrPxK3AiJPpNd8rJ83XIL
LWLIatBKWBgOlxRKYJgrPQgjPItMePpfn9LNFRS6LntOWv1nLBn1Ybrkkg0a12N4
N33r5VJdWzKxKOIhWOYi9GiiyxLDAD1i4puW37cnvs9b7LJSXwCNVBmvInZ3NwOp
Htf4mrDjmd5rpF3eMFOFjGq56vSqL0iw4EzQDH+qO/EbeTKkD5prxjeincQhhPw4
pUiKBWe68SuJPFhTwzFFlMSLHas62/pdeK+ZqCr1EvzGzrd3YifQwrhi/lhoMSC9
tosbatBLmxwWrPfgz7gdN+FhfhjczS2Eswg4ubFWS2iQjwJXI+zeAUgemzPxvIlr
1lKvVYu6XWwtpDrnGnnV96ryCU0PuyKw0qB/znKh0HiWy1xHl3KErYUDOCv8Vs8w
ixIxOV/Ntl4fIOdAyPSPwVlkjvEYsv4EKvbPk5Mod/NMk7TyR9mhOFdjAsKrTpv8
RUqt5WRzQA3i7dr/SQLhyq8WPaOHSI2Td4QmjRXU7EwJKpM58pBieEMmaIl7LCwC
FFer99t3APmqphjr6C2hYZo+Qv4pJ8kPPztijkaCcq5R6/0YGZUjryTHCcWXYt4d
637mF7mXNkMYPcT1xNGgNvNKnUkEjhJv8R+gp2hu5TlE8WNshr3ZWr1kXrH4wRBJ
z/l0KLYK473KLAngUOiLgLIEoIyYB8g3S/mwLjl0KuZ2O82knjdQz5bUhZOBvpcW
/op5bALZPNA/v9ZGxOqoNyASquvcjt9j48pQwmmLGKYdXm4rtch0OthgmTEZGKYG
6ORFFldIxbizpXs48EPv/FhXw58eN4Wm+qnCqvUv6gDRcbML+jsd7SOjCPQp4Kym
nF9Cyxexk/520Inq2muHIG45Fsr0U4o6SSFTJKIOjYXIfL742EorAPNtUMNJp2aa
wFF71cOvOgX/oTSOFwdLZchpGz7l5WuCU4BcoV/7Z7S/5bfaALXzMJU6B1YqLJZd
OWh4GcoRT+lRLUbPfELQhqtyV39fCFFScfFHwicxff8zUSAV3TfwKQGHnvl4+pCX
C/8MmK5jlk9hQZ9CA3tZs9ZtmwZbzyID65crDI3Yid0s3dFoy0b71YyEPzGsz+fQ
t6M/PCEdjiX8dwrn1Rj79bWpQ5FL63Tn3uTd++hJ84wvGh0NdcRBIvo91qMEZ/JC
ugy9qsRjRYv3QfegHABhQUT4HX4raVOBdzAucwV1pxCmI02VdaJdZXO0DF75gMEg
PrYQFUEIx//9AwXFfaWrjxHCqaD2gyAfu5JOY0nRLG4RRzAJz96DzWiePuYdSFtG
U4bSjuOEGlCwGSXODuK4chfhMLz1yv5wVtzdNjbOKiE3LgS3d1ml8ZHTnpzu4eQ1
JmelOdJuOYknGnqrJCCX/wVFvpxu/kt3aluN9nnUgNBqEykOZpnpctxCXpHKc1UX
TT4k/Dc/R3L5qvYtjs9PRkt8a4mwirmyJlCF44eTYW9eX6cYs6yYS0FQHkTf3OIT
KsqTrDURAmotKbkkyNbQ+HdRWA/dXl4xlBbgQ07AXJueQ2LilBuZ/uK0//jY8UCF
9AY7yomcKNYTijSKEQckbq2HwNL/sGXNA2pLt84JMosDLTDfEE3a4JJIlzYGN3Oz
jskOmwlu8bce6zTszVe8XpuhkylUtAglFRoCgzo6BRbrHMeaH2Mum1m0DghxgvuU
drPVnCy7/U8VenA1/lXNkK7ywI4JNrhQLXvpG8oSEZN9h2brurbBGcMbAsKXulU5
DiTIHzNUFk78Wl/XS1TJ6vtACCcTmpGgCfw9IO0LZG9SoncHQYaQzi3JIk2+QhzP
a1GjcawB2/Xf+08ERjROlIneygKAoGAh3P8RQJHvvsIliJGsq7IjTF6log2U8mJi
4qiS6iT8p4nWmLSWN/lQE3kL8NVB4kxn6udJRGfgYR7brsx+JGa71mZkB4kWHEXM
qgk0tK+1m/Jfsi9sjPVvXkBbzw9Tf5QH2G3B7BVMgyGLlxE0NjRThkOM+jyytCgm
SQoLrlqywF+y799UK6GCiRVrWGGr2A4db5FBq094tYzxabiHJVofwRJdXjd2Pa30
jt7sOyRBfPJzR0Jp2zsCE3Ck5omHPN41PnjHvm7Fhhkn/gGEkmA2MNeyZmnXYXL1
Y1wcqCF6wZh7w4Xb2M+L09MqRqBC92FycZpxbWgukEo4DZ9ytxqFFHDnOyJggs9D
MFT6FgtaBorjJFNyGHkGg+cvfur3XcWnXtnw4ml9ZVhGYX2Qp3Oc2lJOecd5SQDt
7rCfzutJy8BbdOUTm0N6EJQiM3GWKoO+H3PN09z2PdCB4CZv8i6otOshY0R0XGt8
o8YDAyIUQOAhqKPcDsTYn9dUKYGI9fqDseprxTbx/fq0VHaD4YcQMBet6HpsZHlW
LwyfrDfEUqrVhzhh0PqAooosCtp69LjSU/zmOcY1weWGfuBNyM2KFQVM3dWVNXou
oqSanSBFaQYjLY2zxi2OVmbZdPlPcprRPK1PtBDCXGjofeycJ7CHnAbDNA5DRDFy
qc8kaYqQ8k/Q1hiyRsMQxJ7vd2ETb6836cRt3NWMalLIDaag2/VVyFLEyBFhmq4+
CObkIk3vbR+JfN5/suz+E3/Fi97BeuZk25S4cDv3dthBMco6BFDPTjR3kdtWMGAZ
My6axjZlQvxhwgW8nRNaFkbxd4qATXsfh5zVS3Vq0ZVKKwlWff8FzZER05RvuLil
8V59mKSvp9lN/j/Jt6ZSpJCfDiSSDip+aElYAHv8TN5ruVZR7D527sZC0ptIb6IZ
wX4jr7A5k9LMwBam1bEpRm45vCkwq/LcZL86KBj9/oopp95AoCAHS/fqjgNcheGM
cS5J8r5vPlRWjulguBO8Rq4deyMFJImJkkusnjpUJDbaFejlwEatpznW9AMzosld
R5zG9/vIW+O9syw48amGrUAtOLQS3HKWj3sgtqb6QBL3r4FVhRgys+sbDD7oCcRg
wHW5qZUD1JCP8Sd6gjrEbuMLn9Zyf+9EZ/vGwq8YDzVTap9X8tOaUGQbuA4tJQal
QmNk+nFa2lQXHblzyKNOuMfVfibbmoKMNshyF1vOFyw1Sh4GMumDKCzCJuzvao7/
+ppc6WUvu0wSbtSy/kcHVmy5TGzBehCK7fC+FLutCtStFg5+daOlxvgOhrE/Dw5f
7fRlE1hFfLlxixuZ52ZXHrHdIw+jBJa+uzvCVkBatwDFsH+RNU0ixYz25B6qVjjW
l8QiAQbQvYF33JS2IRVMkG+InBEu1wIKCpDADRXgIFCVLIVwTEmHO5NBdjLHq3+9
FFgswz5hoOcrvPdubg/I3WicDE4F4bPUUBrSMgpnH4Ty7IjtSdT9GIREGaqFCTN5
94QQVehxe7k2WvjryYfXSft3dY5H1ytEGJDaL/LPJKpqm9dC6bKYSUTVOA9AmVAZ
h1wcXwd8Tswpc7bk0XIBBLjR13j5hBCOPlp1vSBJfPEyZmBgCrAF7hbEgUwE4VWo
zemTHkV42KljIhTFRbqgQ782cxhADbMcAJ6fg+FmwcXOVttSubdINKIbVlyslqwT
UngOLVl/xrGa9vVBVfRGDoKs4IGbTRY0eLQauaOH0DkyyHLn4CSuZ9MXC2IzzzKq
pFfB7IviWaURpwwtqPjJ47/RtWRl07cHpQGbuO2e6QRONuDH/Z8ARfInKK/fL1l9
4Up8YJNhcSMYnxzFSOILIPaWIfwquUJ15u11rLIkkmFfoRG8Z2Ys9L8wqhZemYiV
FIwk20U/mjvwctQcI+umF27jPR6eSSZuELn4dedy/Yp29OrI5j6dUS53tc8SzAAK
WoP4yNKSOj9950c1le4Zqg62/QsASMm0N5MW/AXe7gFSA57F2BR2QitR8U5qjHFJ
urpoyMzABDzuLnO0RSlM/ICVQBfEzF8dlmf9j/+/zni10QC377lt+BeBhI3Sj9b1
s2R7DNFtJsc6QTJnC/Vk4JSif6rpqSmjXDb9J6tcouxvskQ5a7TjCW2A+ks0cVBE
IUuuT5cPfygNsQSsKkoKAK847kpWYcV0h5fAwnwWL/LW8bwPMQAg+U/kzld8eq2H
5YCUq401unfd87pdy/5RyZ8Ph91l6mh1Wa3QTVVCpPPLrpBwdKAEEV6G/Hy1VjXI
Cx2GxPDn/XZk0ljhbXGnVY2y8yDKnzQPLdSnm2oODro7rMfC3B5r0jdi5fYDRNVS
HNlSlOQxraFYqNA5HZHd1KGP4CHEh7wi3voP1zzx6M0ikWFFGFv+kogBD++47Kxw
L3SvTJxynmhTeKpX16Mh0XDpHSnyAqiNQjN7u+WXEWFHkfLi6UJhtfS4P40I/OYk
KEe6fNn59kAUhPbQ020/dbthp6lKfhH53CGi66wrZLVsPslXcSFrWggxO0EU+bRF
ZYdJY+yO+Tn5X+FBPAGaQD3JYOrqCAwJvK7tZklbiACinjTcvu2XtORXEunZhuWj
tnvrNuBNGoWs0VPngx9Scv1+e22cELSF3WRYDC9meKvU3naKa1rC+b3hJE7bsj+e
kxdQ98MkLUBpVoYl6eudXflZDlGDDhj/Sjnl9gUE6ToHMA6bqBRs87ug1d3XTnqn
IOeHTazLLRJ/FArsIZtcKAJc5R3RxW1OSAkGsdLlEFidYzk8ybLihnus+jT5ebpX
bojmz5sPVKbImaeEi67C8HJbKn1DRxVXgppa26Iq/HibpoZGO8+P6BUE5cwosPcX
zVdBiZ6nFvCs/natJcinqQXHOUY7ib1M9pp2imea7x6BiI5YJl5a6C1acLfVPWLa
AmIc0IFBfVYyQehs8t6lOZNDLBMN3qW0n52NFVvE+AKmItX4WSmA4VXXMHHjIyEx
fowIxB+/vyYlC+Kn2czSAb87WN1aufSKonQ0X2mwtGg0Ddu9hX+5VcV0eSWENrJ8
FDGi12nvrmnXpfRj35HLxGldjr8vxtaMa7Dlu1ebQ7Wy91By79uibpUTKnl3/rYj
15glagk8Xlhx+203II+YRdDLw0rPqRRgkd7SzeaxRYpcqUhZ9AVWZp60h92HptQq
2Kz/R4kQgj6sBmHVzlozz2jz9LtVG63q92W6JEh92stCSSbiEdawey1hGI4KpXPH
O9uWvCcVIvgbRcoirZXbyagDO3OrgxOw7roI05BwkPOgSgpSIOCgc/3Glob/Q1sx
AdFFcMDzx6GxecH7TqHEOboH9hZArq6S7JmYQt/FcXZltZcyBRYebxmCJZKzw7bQ
kcihCqUeG08M9x3RaGwROSbb4B7yqCN3BLHKebyjIw7rTBXyOb3f77fzLh6WrDhc
EHtATDkd4O0UNBcs6C7fh8NEiQERTyIX9NLTI8+ye5KScw15g67Fzh7p5bE3/fML
TTYoe6+uAf9u0NLyg2kn3exDrLzLYN5AI3fzZrK8ZWQyjwuyg6r0JxpfMuct2n53
R6MHYfAyDWi42UYaaAbWJPl9rKGM8UFNgwCEhzgkpAeJ9UsjKcwkNvoM/ZMRhfpj
MHsoM7E4JP1WcY5wBukkKskJdreH0efxLgmStLdUuIkanK0wSsl00MQloGBcHMPS
PvdchRwpUrENFGVYJCbWsMiOjo0plk2EAZEDadJ1Ggw3UYcj5ZjimFqiTo/KVLd2
Vyw1i4mvb9ZJXh1WYdLIKEICabhU7yF8aHsAiRlQYbSu+LQnwILQ50qGH2+0WT9T
RH8FAYnd9xUYCOzxJ5q5dz4eKQB8BrffBFYoNlHY3bZV4l6jJfGJqA2MNduihYRX
80WEoIX7Y75D2E+Netdal7bWrU6WqdKQ8wNBv4q2L7p54eV243PHgcw8kEgPtBoZ
72ZkkwxjuycLLJs68d9ovsVBAWBNXk09G4gevXnuG/XvmJn+7icVnKf5ZG1wZfdy
p/miuQ/IILlkdUtW4iyIAigQn89WcthTdztlLELQlpnTG2qoNpRnZiUQeEBslIVk
/6lP1gwbgMiFSO2i8TmojhDnHUhXXCiF9lJ7YNwqmMlid6ugoejnVJFhY391ETau
6Vp3xck05kFtdKqQZlpmT92c02lzk4lcvyvADe2R8aLMvWQTpZhPB2aEh6gklHv/
JPs7pZ4OOmxKcBgZn26DgP0SilpAMtf65bzxo8nLefjRM/c0P6DkRfqH+79hz3i+
ygFygY79NRElNMrMykFlOropMsCXgf+KmmhiDc69talDzRZ7GwKnjhwTY16m/7gD
fWGhfMx+WcTNQQIDsuiYElSy82vsoc2kUTTHHN/Mmm5NOA0i/+isAyJbfW5Qag9j
RzFZ9LHMjN79Zk5xsgJuG6NBC3m1wL8BIPBzQTzgc7bvhXwOoMGmQVVTBUMjRqks
/SsHMYsly6QWAioCMiT6uxTlwjR1rlxnQnrZjcm+uO4smE70oUFVYVncfCYWIlOx
rwU3CGJlYO+0mDYfS1WuLFNv8D3cbWzVEMITfjppojspHheNvEI11WtJpJ8QWOST
AnnAO3mneZiIzqKavJUCCZ2BnDInotpOpDpeCv1rNUZd+N5aCinQVwda7PNmraub
96RaRWQWDtMA4Xb+Cc1f2hckLWkF4w87o3Wt6hB1kDCrF4KubHk22pO1LNCWqoMZ
mNtb6lR9nmXDA5t+QA/6zKz7wkcrHR6oOGQ8FKcMmM99hLIy38ANwdMwUVimz7nb
7sbKMq/DkGRXK1BexGs5pXFP9yK2PgDlex6gwSB7XIjoNnE1pC+1Vc12jFysVmSZ
+6p2oCUby/Iz4e3cSS7VXLea0yLHyO1B+mvYGSXEBvS+UCmXIU8+AmxSCqFXu13j
zRQieYRD/UPM71r+ydKo9jiLNali05sXjwZc3JQ8Wht2WbDuMBApi0VpMO7tK1sZ
h7/aWURTt/fP8hAq0T/4+X78GfJgLDl7DvXqkuzmPL2d+jU4JY7KlEgpdZKjm58X
4jbdeIeYwxNO2z42UkCT/wB8T6Lqu7mTI2bX9KTYzxCvK7z0wysOCDUkkwcWU2cq
EnkkFncTZh+cufTbyxgWLajmBWqgIT7BigLjBQx+RgYopGzauBRV6tVZ4sef89oV
HU5nku2HzQj+neTRklyZ17qFAW3vioVukFuwPNoRDD5l2ugAhudfZ8gFxXsO3GG7
HTP7S1vPLFwoxUzE/NKg7SRa01fFRjEHavy7836m5FZjz8JEmGSLAcJoALkCtysj
5dnVGvfOWhxHo+tI0dfVtB4kEWFwYB6NmT7p5JKGYdWXvwZJeWnNPZRNRhzC6DW5
kQ7xdfIAEY10Upfg4v9gVN75PIFItegk/qHcdxSxqP0n/ylJAKnPlHLguMJEwY1u
zsKCwyrsZHX/W5wlZW+52hC7r5rVK9w2aSXhwj9I+DPtjL/qMEj/oaxNfkw4NLGm
d7cUIXVnyMIl59/KgdpZlsIg+nk+q4OMqlGJPM0ycvY1NAH1dPtchkIDCdXgtK8a
BM4wN1DmL1x1rfGvxVC4FbASy7TeIS5AjNx/nXS6LdGWkXYg8hkdq1mMLT7o/cXm
focc60yIbeNZaPouZEZGJCWBxtIvIwnVH9UuEDGO9xC3Sry332C74QguMBIhqka+
fqDjusR1y8BkV1U84Bx1a0viAxYyCbwydJOuQPLdWHG5Wo6VQcopnruGONkqUfOh
2M4eiULm4uM7GH5JPW+Jvx7B3VcLeo4Hbx6dCjCUSEw5FMBgRbC7LtPSKl01uWCl
mzyz0GuTQOMpcxe3NzTYClHrefh0fy0B531XT72FUVrNs0WjgXJOiUaMkqh9Y/fg
ZetQ0zmohC191tJ0FV76XXAiJ8GY+kXgBQyqKVyIwu8OjZF32Ueova3yWQGMXYKe
jmv4XwIxbDuDNxT7gplifs0Qxi8qRe/BJLIHxP0aE2F/3Gj7js+yuMinhPWU7b6l
nqssnv27225S+gQjlTDeB+It1jte4e+YPQN2+xjnmK1WMC7lghlLKfn3x48oT28V
X/DyNKx4cjQAoqhKbu2NyYfbN9XlI7kxKNCVJ2igOOAvxtAT91NL+WB1KtXR4fuV
F6WJooXGRaqQTht4bjrQTOhyCvv/xEV+jYmqjrq9WWxtMjBXtszmbqNlvhR3kmS4
d9vsSJrtW7YJGfICBFJkD1GnhZtKjLyHHLko21YkWlgPJjGKus1h8fmh4qubMKXc
o3jlRV4S7vE4IJTypKv+emmBu8O1UhKhK8NB6vEl7MYhIyHt3sD8kNIhETtWMZBB
zLwxVvS3NqlGej5SYwtXrKtvcio7apmmUbrmrKDJkA+P4NURF3ymks7kmeGYkw04
ciIMfz6USqsyf5niU7wE6JhFY2wlpFC0JHYDHf0VfIQkFdO9vg0CQxZgwjCMzrjw
HcRaYL4n8Yk16lwn2jAvFGcSwxM3hiWDqNNew/uW2r0/VySkzwQLjg3FdUugogev
d8hanB61BzXSPCJSnVIRr2HzqN2x9gLrP9M4zlgNrS38Wn1xqUX7H6ayyhAR8dOF
o2ktnoPNYpdgHn6nj+op8YnJZjmseqB4M5cjGcQL0msfITXxAZEWQjjg2UlLy8GT
SqX2DCSFALWYR1KzEZUqASYAsc/UO/ARQjEoC2FM+y35NP8aOgqKlBaZgChSKvZE
0ISKfIg/GMnQHmaGujS5Z4f7UaIfyFUxlEZI8fhrS9Kc1Q0Eojv+WhVaNklR91BI
rPjSu8btydgxNnhhK5L4JgqmHwtNYjDq/z3F6yHSZDvAW2AXEziHygkuGc82I2uO
JLq2KkJZiuKnbXxY3SxmGe2usxVPiwP8uPTbvJAonIGn8HbfUQid6W5kJc1LA3gb
yH0YNCB/fKM2k1PBxj2o6AQzzaXtS9xoFldDUkkaVSxOBgqcSxcYmtr5jGRc6AC/
0e+kfg66T8J0RFR5gAVosmUrhXYRfbCap2m4bPz+9GsWh18NL9NZm/fJNBec9Xtd
cW2zQiH/8fiJsDVX55naoQV11v0m/hRClWE2Ih7fXT3BKbo1UCMql9NDsL0ZfALU
yzEx3YBkKPVDSf7OQejtcEvxjHy4N6HUGOY6EUcXaanvYqzXNlsY2x0GXdTJ6YyG
ZXxrRpfDSS3k3ukxeTN157I8iOVRXQ9bZp1cqNIvhKa+/fVtlvGLgrznToQ2FEQQ
uE/NNE8ouGhOysmrN6SjSA5odvWvhitNL8c/9/J3ZhjpEb7HIpzSzRpSUtMseEkf
KJK3CnureZkMBkWVUbOFDYBoYj6W3v6jVK5gPJjtsJMmXoTfusbp3aFTTUFHzIMl
94ZFldXK8NIxlZABILhSd1qilavxwB9YvRqk/KgzrJuUsd4O+Dgj2OtiY6D/TnpG
paFbVc+ac+pyQdVThyeS2wdbz3rq6LjaZJoRK+im0BeqFb5jxVp1BZHCxUb926yI
+e2QiHda83D786MqOD2Zo2jFMtFsKo3IULg7khqj7E6GxZfQbaODzVlo0Wzsmbku
N0N0ocj9b89L+4o3nNdD1lRyPA71gjoZ8FFRZwWLG5gGUH7UOeV/ggquSWHcimh6
faldqDzFR/Ty6MhVaMmUuhFgWLJ2EpwMiv81Bd87BPb/Kf2G2bKKoLFscJqiW9Q/
9xiSxKkTA3014NTaqDZpBqeEOg4zZ6RF7CdslMc99dAXb2YDlrypH97wZSr502em
Cs7EYS7LG05OKP8eoYRkLkAmD15RPxPh81hj07BJlfTOWcOhhLggmpfKyp5w2CbR
FXSgqkAWoxs6NAS7RgcY25Fp0aPxgo7g/+/s6Aj3neubCL5WtzajnvCtaSRedaGj
YgJcOZhnTQL6oql9YoE6NsIOCKNFw7hoQnrNaAKgKQya/e3y8C7Z2MFourMY5Ni3
3sq+BXwoWW6mP+iyRYsXhgny2j090BF3Inqey3eaoExbR4eGHSkFQ+p9Cp8S39h9
/SDYF4XuWbWREmPRBmDjl+Y4mf3FYaSeb0Ri2GhLbH/7csZ5KKWDZO3v1MjgphVJ
RPPe6IGdO0GZ6rB0KUefjCcXw7mKcNdjWSGECt4OTbxZtvIwhLzfAcu/Jxb8g1TM
/QNAiaWiD3Q9859L/UyfcoNOlngtJJC9koPGs41xxMQtmSYDf5QcIARqN3Rxk4Tz
Ooe3vwe4i+m2r+6Im9DB4Foto/p6lzPVLsqi4D04AvTWvVDHXSoQNWzTGEUrmeJq
S6a5mENmAzczP5qFMsJPJ0t6VRAmJKYCf26WDke8QQi/4M0XQ8ZecUgS1KDRT88q
ob6FLfMaTd52474qTD7QDOqPINocy1XPhWTI8oZjyrWOfmmlRnHTt1M52VSO4ntc
UuRPgKYjZ7HNjZ7k/No/ocrEFCa7/Zbu/7zNFSf2TZlACvacZnlFQJVX8LVW1Kj4
UQjRPVIwHXmRyhVoMJCRAQL5U4vt+1Mg4cxpbCXVA9+AyWAdZ8b27DjpqJhgksYG
Q++pP/9KoYVl9SzR4zeYxN9JvJBLB9ZAzbveg64NyX5CWwXziLHnpi6laS+aJDRA
7oJgvGC+25ZXN9zje9v0IIpFvJRFXUFbKogNevhyPKLitBm+URZ6KNO+aj7b3f3e
wwnUrR7UQBs4UJgz8O84RaUbmlB9b+6tYi0xVpJnNULJT19uZ2kvc54tPLQSHBBH
rAkAfmnrGMdCnkMiA6LDyUPVaG1NvaM3bFLI8wuNC31pJNy1CjTqf2Z+22pwppre
DEioG8vQdYzMtsC97aFHYyrTMitpMyqRTbWn9DG8Al3zLlurq5kP2hu003zX5vhA
hnb7w6zvCBm9yoiZ0+21yO5+gcgw7SQKdTHr5mNHqVLOTWkWfd6dOryPepoRUXKU
k4h9FXGZ+9F+cI0J1Q1a6ejR33TkhDtmb8QR1CwgNLZV86XVsHFFBGTrGY3XDFWt
vJA5psoFgCF6Vx+mt+GPOVf/9nZq7B2BhVramw9gXkfi6CBAeWMuutbpINZ+PHNA
fGYGAodpdC3pS840WqjS6XVCN+VkumQaWriPzewU9OvU3vFEYiqxcL8yQeA7Dn2e
4QnUBmDWtuwgOKsTSAHv0iijOGZ5ZrJLDKNCbsNXjEdSoiG6W6BqUCiD8aQSh79i
RgIrJjK5qvklD05nDTViB6NnAGatFg2i9Y274r+Y27de81DyA/kGTdH0tDYNYID5
DsWj23ASTQlOVJLKyvGziijN+TzumxylRWLykFdAui6Ks4I2l7/GpifTjDiKJZr8
M78eWv1QwfI7t6wVMubpqOq6Q4+H2u9VloasNADo3ZBjhSWv7+a2QrSJyALyuNDc
cvOMACIv3r5xMDSZ9Gp7AXI25QoKxbuZuQzm75P8nIdyZK18Cn6Y5F4UD3z7GLEi
Tso/OtVo3T7dqR0MSNIGOMhifFL0jXOjdx/DIMTI7fxONwFBDtbqRconISAuo/oN
SsZ17PSqf1CiKJyW4mp71O3Fyc90APb9fCu8Ed6Ov7hvtuijziGTeapkDZRtwucD
ksr4Nl0WNg5knOCV/VWkPwAA/nNrdWiRHRlmrujD8N7ZHAajg6aTVcJS//rH6XPl
gc/R6ssNY/i/XcI21JqwVyIDQyldUnb9tJnzUZSyuARRJBphoWNnGwllRaKQz7Zb
NWenhKFn8/yFnE/ns6H4c8s8phdyD7XnP78pBgK3GFseqJ0X/AAJT4xQQKIHIACP
MaVLakMP8Pv+YvrV8+hs8wNGnTOm+Iyqrprvbw0+9n5NWEs2Z+XKU1riuk41YZpQ
AzvMYW7ar3WhyfwzucQ3cMw7OE6TmOyvN4we4oEiJLBAIQlw5TQ3OjAZ0sl578Gc
qBSFu+XZiSmNve7grVrjjtw0m7/Yj/J/kQt0R0k3/vaRFIe1Iw5pGCc4TvvlmDeL
4dGaTkeBiWrNGwrDJmzKPq9LKDe7VQaz4PbCTUGqSqmCzs3XMF8FX6q1j7Ng4LfJ
lk3pXhxG6nrfhXRUfYeBFUDcr2k1/7GQfZwtMykb+dV3yE5Cgos/0eqRXA5Lsr8D
D9TZy11p624JCS7atk1EMYS3Lv/FuQowEkh6TCPYFmATvoGjA3q6qbD8G705CoeN
weito0xAX44z8nkBSi1mxXCVj6oVNbB5q5YbHaC8J1jLb+8i+KqY4jSJZS/umS3u
OAS2IhF+xcI2AgyGLEAUlo5hebFnMS2XDv8nVZmk9DlZZJwk6V08bTS1wzDKRpXX
WJpeJptUX8ekoNVCINBb3uIFeXpg9IO8oeB3OB9ublHHNFVLBuXNm2E/JioPmTBL
Ga9xAaWqZQXvIjCiWD9l0RFPSCQ+oLJPSx5WlM/FlZPIsZ+T4oIpCZpe4vJjG/Wi
uPm0wDC4Ed7wxzOpHlaPOnjkxv/kqrv2bf6K6iHZfPEuxt5FilnP2Q7lONl34T7o
zng33tqw3VS7PvQc6Bxe6+bIL00cIqy8djb2rsLQNNqXPBGGGg7Uc+LRLVxNoT3n
ovKhO0G8D+jXiIogRydjkwurWpY/fybaUN9RuaUcvuxev11nMNYDTCcMOfgvGtqh
Eg+XUKO3kG9Fd411M4ln45v5Tq/pHgv+6lSCYE1S012QvEd+AV6inuj6J0zd4RBU
BE4bSaHpq6JO+UOVcrWF13H29DDlFdyLch5A7kq98nHP8bjCYkebMJ0cSPnpP+lB
WfLz9OZAP8M6DxwtKILqBO2kiAsNNoqcuZ0FIxi7aX3nRfwA9Fdwb/jNiEX8WN2Q
xaSyrKWo8obm0UmMOfqvhg+4+WsrQMpMdHuEqTnmVFZUnR0Xu5hEX/r9a7Qekm53
jJUktYnG5ZWKEAvQvPE3+ErMHMAwJkVvMareBADOk0eORpeaYCy7O2JIRllRwHJU
QVTPdqYkPGx+3i/z03+Q0fef3ij1QYWNk0pTmNt0aKlmF32aP1yzf1x/lH8/SCMW
iWiPLDpCWKOKfeEGWLlVL7Idzv0n7Y0TSnaxlPExwSfUQHDF53L3ZPaCJA/VLnPL
PASSymgI0ENFH1ZBguYRzIwa7XXm10vbHgS+svvRRCPISLyw/g+tmSCMoNlzBm0R
bJ1EENpLNmRnIC6e1C/yB51pdSoHnjKTD4O0ZVUTDScukXPyLCxc+YuBAzkPUEMb
ARKVJYaoBIGZPfqyS7ulbqep2rm4t6WXLiwCQjDkuUdGH4dgD0xxCOq9Szx45Y8n
WHbDYNp7zSQ1S5IScPiUkjl3XQi6/VaYulcVdY8chwaRH1PHNbkaBGinVMs+MtBp
ytlHVr6VJSfvvLD+tMxMhzbF0nslKPhmBZjWbpm7GOi2WlttXXCCTZTcTMU8jFry
iJAzrFCJQ15XSvTxrVAIq9/sjV7Vq762OSih45Ohw54yLfRp1U4j8OgP5PBaoiLD
mZZ2r6zylOKeijZQqigD1W+roB5OTpX+iFQ78W6BCXXYZOFAM9ye2WUcYl50xsmP
ACCrwV2Gr5Te9Y3O8AOnFYUNCiB0veqrcxe9yHODahRDgA5vr6T/MTDOJFrcNcQ+
AaR7OlfTPOaF1r6zrBfu2fVO4iBs+0wxKJT8Twd7Rp7IgD8vs1jw8N4vI/eSzXkM
unJnp0Yn4I1lY3AWjU84LoYGKe+awiAQ7YS7XjL3MO1GQ2PqR1HSdWV8SjYwWgaS
LjdMarkQCFJI1WM7njLpQSaxO3FrMzvldTCXXhCVxou8akHCeXOqrqz4OSAt4FOT
WnnSGHX0cnCzhRoTk1CLv6JtydnF4rO4adl1YESEPjBrcvaLt0pYQsy61+1XooqC
1GCsYo4zqGBv4vvjVxpo0HtqQUA8sbcEQDMDogaLCBCLgdZJn/eJe6Gqz6lPN9AF
2tz1Dm0vBuqnc5QAB21tjX8gVFlIz4a1Lj0qpmVY12wpFTiVTYOuFuJb6HXrc1du
/GidoDRIQ0E8cGGuiOjER1IkAAlpOj0qGzepX7u8ekTA/SpB56LHa4njf1MaSLjS
FwE7opTKt9nUVmfQ++0tsa/04xSav9wHjZ3UlQ3PRqWPoXI6ZZq2pA9C1al0oYb3
xBbHkwfOveho3qzBc7m2Wu/PVsf89O+cu6udn2tBDhrij14RbAQcM/kB67ytyVWP
8utYu1AQ925PGM21eRkS05VKQi8Sdxy06Jg8PSgZxZIB8oAyNzalA/jHQbubaW5u
Ch+OxVM6583bRMCpIDnUH3vWBezfrwpWv+z3m1R6p6ejvIdGv8xAahkpG74peqN/
PMIcHiDtmjqr3DlOXK2be6wABlvG5zBYLPlAEG5PNoN/cmRKp8/aIYo4gm9NEmIU
TfJlOWlgsVVGADQKfJ+7dofHV8CunbMjHdR10y+4Jr2dK9c5HRCSinhW4qFD+9n/
zu0jAHEScNyz6+rGvD6d66jCEo/wac89BFh7N1LwjElSZ/s+BhmWQ5nYvw7oWww0
aQWBonFbRdeTKFxSZrlhA8c71XrIvfcPEvIOnb5CNNxV8lTFREQNpbdWfbhU7eGs
QuZj6uajvg06ewhZUVNxn6IafC6E9UccFzwXZH5CytRZrv2vOtVk/jYCIv3yKZ4v
s11zeSTCHEqHK6N1jtUBVnJIt8eO7NGuUHWpU3QQUX9NvIOmmCi5vd6V+MRMA0j0
bYrioWrxH6f4r+oT0/vH8AHaeUfMJ7p0JbVLmbbX7SGp2YdqIC5KI1c8Jgy4Bz9M
2IJ8YGiOGbY0oNORVGLZ+TtaDN/k955bQ92ZpnTFyqFcp/nhh9yoj7Qs/e59gKS3
ayYHSEIruNhKY0tH508fxRloH99HmVQP2D/sZrc6lKhsQKcWpuZFTZd44n2czoo0
GLlgN5HUSMSRe9lm+WUdzPtNUhSpwI0Nzb7leUKU6omcdB8KLZQpRMedDV17mxQP
afgfQ0CCO/PXxKzflz9rHcH3hFF7B0HKq9d/KESzGKnpIWSnJtU2uaR3OXm3uHz0
4kiXcNQCyMQb83rW93YdrQe359ICD00YqQJWqC0PK43EQKbTi/IDkKp+PW5rD1kk
HRhGQAeIISucA+1gx9bvpblnWd+ZaRxGeT7G8jfZcqZZt46HVc+pFeYdhQEA/kT3
EvnzY95mEm9eMdnZJEYdlbgyvywYv52NrsKlvPlmgtopnqhWIIyfYm4QbQJXonAG
zPYOJ4Owa2F76q0EpN53GYGb29O7pw+l7jeIiwDSusWAz3ijNV8Bva7xMIShA1Au
+ZmKQPVK3u2eEGkIXrR9Ttm43sk/oLrIDgM+8o6/qC/03eaWzY7d/YQqE7Y6+rq+
6Jg+j+kkm90E6N+uwUZ2TRUlf7brt/Fo/9mePMS3G8Ki04vf8LdJvr/0d1qh6fR+
SZYCiZv9Nk137QvWJxd/S/gNf4uCHWGDM1WekNboowc0IkiRquZ1vnR+1439odZY
BiN3O6l39MFV+q3A+qNr4YxHVzmzK5KkqV+w0VYsOxwATKzjnbsb24vvusPDW3IK
6HTPQvEnkC2mjziszgeFUOv//XAPOVGOJ+LFDaU8RsXEj/OE8K4S1GQYkcqw4YR8
KjKbiC7aK34vFAlpWNP+0xq4RF0JBx+7eERGf1jq00cPnc9hZU43hvhPSQLMVnT0
nu/EaQBuluvFuaVSTD3TZsFhj7euVLxLH0rRh+YSx6f21hUZfOjYKmdBW9FFOWaa
eY/rwBtxq+ChKc0TW0Ff+qHIv4gINz9obCC3xdg/rhKDBAUko8my75kAwej78Z1/
XmRzHReWezirqFzPqtSLhrgcqBzrtI3BF9pd7oqvxNE9JyrtcSXqEpoB+nuhehX1
dnHUUB/9LjuXBSE1GpCnXjMxSMGQ7RdKfVyfxex3s/+sLgpgk2JVEgi06v2xnxEO
uOfq1/5KVPRoGDaBOps1Qfy57CyCwDfnQCI0Cy95500jg42CsGEVpLZ5jnb89mWJ
vnxoHcvJmjUemVcZVm+ddWeXsjkFNjqyxOAj0NMNuRSXQFx2sslPi0jiMFxrZ6Rx
gPz5mrz085CN5yNXN0vjzfyEJQIFi6WelLCVh800mtKwd/6KIm9WVBtjtz3FwxO5
mwVfYAja3DeBtQMxpA6w1BWRWECO7BIYt9gtsEn9K6lxaBocpdtsr5582+nlSw4r
Z1uldVikRkV2+LEofVcuqahnJtPqiBEkHa+0lSd63iQP9F9/vhXmniwR9Arf7yLg
ySTYxV5x9Z6J/9jhQalNK/ppS1fHJAn0xfHi7WnfGTE+ArP6uxeTtNUEe11Rk5LR
yP8WUJxIexux3WUJCcgdy7i0tCBMdpDrLhXlfcxEqkcPOHI8ugjcnomyL4fhU0J4
f2tRtd3uu1fkKDSYx7RRj+WWp86HSyqrU8irAK0Y418SsdoCp0G+RCjejvuivtNq
X4ubCtZJLtKqMIcUgqiXSn5hf3DIKTG2cdvFl4BAzknq5PNswnFANN4Tp3x7nubJ
RrJgVkDK3MIGSIvFAuzlISIrzyyHFvMBGcEscyNt9m1XWkG6uMaSQ1NwQGcRrxvr
Nn0qlkHjum7DDjwbQyPk+G6FWvB55RsxMf5gN/+iqSqfgWnwxfuxnzP7lRXrcxIu
iRqG7Kv+2sNhmnFk4LDI1fMqe6djdiSyShAfzm8z71Gl17tKQs7LCpH7gFR+5tRr
nPCEEqn2Gk+DBxA/5mV/tyavpRMbDD5l/cCMdf1nbVE+4tKW3v4kB7KCbo3dVIVm
FpaqpIMxM3ukI5WpLZS3W7Gf+wu8LDaLvpxycWFh4Y8LB5lZvLCJY1VXyAziHiNZ
eTIUJCLB3pXF82OK0vz6usqZpdkdjX7oQm8vTtu4YQErafQdTlZgfZ8C6OT106lK
DQfogCmADE16524OJK4iNJxedndrKiIq7PnyGJLxnelInrTp1s+naPInnkOd0F8Y
AwzE66LGvNHokVCNu55KVAhjZRZIvGkRWJZBuzMS53ISY1DGnpkDkmzTOUGkcJIv
Cik9poiqC8T6QM/6BTpWSD+oKTY3i0Z5Gx8cgLxxUuvY6WB1CvVLrXw373HNUAZx
88bzxiUDPLVAHVhX0iTr12dW4mbq1IitVEOYfE7HaeO/PSDm+xGvSS0sROTs2GD/
KR9+tohXzFBIEw3/I+0zB5nJhrLKQQFI8LwDPgh4pwUzTAIDRIABymp0v7zA0PRP
AW+qqbm96b6TN4+dkd6TYylPKhUtIrflHrmS0TSltoq9rWnDtnz10B3p9jgr25SK
G9/YWyyDXCeQMG0FJPVQSNlgsp/NGc9YGg3r31vvzU/FDjPXmzzBfr4pLxGaVOEA
91CNS7vPnKOPUkECaTfbqC+m6t5mA2GLAgt46fHJczuEBmxWcFWn3FnPuduGQbih
CU0dHMCa0+rGoyL0eR+pvvqaDD31XRmEyzF3cGrWWelxUEK+5Z4y1crKySd3j/Bg
dBE4vGtxarzlq6g9WmgA9FJL6/OURp2wKXueRiyNuQwTWI+NUFJZr6SHHIiy9PgD
oGzkWpOUN2BFxwrUmufiJx7Kk4CjRiVft9phxAzTrEXghdMcsTEtlF4DGOkLMdmq
ErN3pMQUWkFY0jF7CMz1LqAVAqmbUUih+VKt299xf/SGAzLEHgjz+xemIhYdDiRK
wK/j0m6kfHg+X+hGUAaZspvBX5jI3PHOpgeX47NzlvgJPSxQJYyfedDDGWa/8s34
Ev6m/q88BDtlbP/mw8/AO4tVU/mKxW6iLFGQCc5ezTA4bZI7WALFevFwDOT4U2CC
IrQ+uuwtA55nVfDGaFMpCNnBgTyBA31SZByIOs14XP0UztuBuY/gNisfo5z4kE9K
qW9jk4sFAk2ZZGn+huO/V+M9oAJZBFBsRMGEVsECYpdb6jGKUZpFmSRNlZPUDLIz
YODLkh/ruBdz6jLINZ0J3LZGIKT+7EOKcMF0Lauynxl4idEbHDR9FxfNMuue/+HG
93i3FNVcsDTjxbcmEIzuTk+o2ImMD17O2yKVuxdTjjeEtULUdhQGF9BxPEGIdPv7
CfN6IgdCuk6wn3dekGwzR9AeeXuQYHA9L3awFqgYqfAbolBh7ZxRz6pmG2rrPWeQ
g6H0/phFhlofdgKU9PnIukxl6LrmH2wwyjo4RrpgAiH1sVylpUfOEmE6ssGxfVPo
bPIP0D7Zd8xGj5lM1NG2+fVK72K/ggmNzsYfP1wj3sfm49s+RbVmYu1Fa8pCMUsz
ftGs2vl84pE+4CHcxEJwrfFsIZPUIGgyk38PLOXb/79nxr67z2hsh/XoW+BgqtOo
dVCAatyDQ4pQZE2RazY/1FnKlo6Opt5R4UZ+lNLTWKStM2J0P4fsS5o4MRuhUWAR
o4qbii90aR05Fh+CPt7HSXnX0oOmwigDx1JtYoLSXZSK6hPBJAAqPFnl9TtTnnMI
9Rj5+5zNCKSjXv7Mdgb/xzAIkRNxoNHUJHAV9w9U8LSJlUiHU6/M/HwvXLqyVg00
arxqtBI5f8CYSSXqR8CYku3qujb1fCKYjKniKYmD4CRQMsYK4ZMJhf1iqMufbtUv
a/dqdEWFFc2wvLmzbcN4CuJZi0DL+Ca+FnXYE75ePQqGj+vxD7gyxEsiFp1SkZaH
iHEVvzk2VwOKzNpeW1PaoAGTfv7BIOITP0Z4cTo0Xb7yYSLoUWOO0qYQEyLBH1Ly
79ofx68zn9SFH9PiLaXD/1yvrPsuGhXgLNG3OMZCLIxnaIUD9zTLu4EqYRIjjwVS
YB1aULK8A+nqUcpbLjVJ4t6uhfr12g0WNAXeZRm6FeEfIXYw9tbGNCWx0QgvuDLX
SnZLnmXd1M1USD8nJCiFAQsEA3bFseBY6aGBSFfvo+O+5PFdC0b6/XPLrLLqKWe6
8/3Qop5Pg30nEEolPFLwVPeNsPz6UeEH79GZBz/lV6wNMmjXBlhshurHb5cbD6cG
Vt7EyDh4lOO6LRAIN8VAgoR7V80vftIvUuRA2yZXkyimRVEgZ4qrBCdSEsxL+EDp
l1kP6kwtg+Ia1DkasG2omB+GWyGRVCi5QK3x77RwH1aXRSOsuLED677/SqGLi+uz
jJyHS2bX36pBpHz8qRZqMeaIvm/vZqHTM+nW4K2meBpcuxchnsGjtbWFtjqbC+lY
hD9ynYBUNZ+aW+geSE40mBZzH26uqkf9u2VJlLLSCw6TjulMhdcNvKyTCf4tmP9i
glNlngSqz7dz+8OPP4y+al9jw1Zbc8VdV32dRk0PCgAyMSby01dMKzfkVjsKfip2
Kg2HGGB6UpllGau9O1AL0FbwiUU2bed6yl0qBuBAO+C6yEaHtP5NX7A4vD4YXYn4
lc3msmJPsvvBySGfTabvNLB3bjvcaNAxVMcYVvcxJzH9suVjA2eYcMw9WQOKBVDM
Mu8OQwt/ow7E4eKeUtcGCaH98vlHdEHUmc5AF98XeU4E2So06ujhHvdTVkGJ82iz
gfFbmchY9r8kpY4Qvwj7Qhy+6OQis+AXDPLBiRo/EbsHtDVhj9GqV7PyB3cFb35X
gWZDzIPerBCpc81TeRIlTOkaNMpPVXMww4l7cPDMfKoDWBoxT0/dOYOTMN4kPEYC
EyJ5DhQL1ma/lCI5+7+Dko4dh5OIeQXKQHPP3oLd8r7ZpHBfHAoLckVaox4ErXmp
PbNd9NBPkuqzF5ygBAz/3AtpwF3oA35DPav8xhXkS/G4M99ht1Spcpy/2xjArJqI
aTg+8d6eifYjnAwgpXnkN/Atulgmk9ZFufmxcLyiH4sdYAQKK8B5Qj/hqLSb6gUg
PS9+T0L1o6rZ+AjmKq7X2KNuujnNyP2Ymhx1MjIm1fNvM1yBFmDS7fAScFGn7xrc
AhH09XPAeEfdQmbHBNySf4yBQASquXohD9ZVo0FquvXvRnx1siXS3LEEwsgZAGMW
fA3s62KsYWsiawXo2qAO9pq1Sp3G9aIHlx3OlW2xunydUk2iUF3ovwzy1MO//guF
OKDSL/0ExkryOpZIlTqzbwI5R9IkSsiy2QGUBmOHFKy0oaTiLxYcGs9dPRbUf1qU
gdVP8X5ogzWHITHnA4aQP4fSDf3E24NrCO4OmzB4beEcUX16Ml4FjUiW+V7QDyGh
2KaH7x2ylBZvyd6Cexa5vha0BxpHIIUoiKIAqKXIgtjR5Fz/adhI3JuCJUd8qrDT
XKwvKibOAHb5+SP0Q4Gs2FEW4t1GhFs2JlvR4qVF6KmnThHN8xkt4v8lHVnXRO5c
5QvxIQpIzubYIPa7Im1vFmGjNip5JWe42zC/kxlEEmmT+Bt3/NebBesSBUTWFFJK
SCY/X/92Tki1jRZT9t51x6Ib2m6lg7Nq3S/RAcD6ONIhw5+tYoUCN+R8xuHOS2Zx
9GZw1gPQk9Z0fkfpAmddj/7+RLbIDQ+mQXrdWnxTHPq/mLPY2+EoXlLsYdJA7IsM
qOweAe6GzSrpaO8T7CCNpV/l9Od1ShsNrcGM09yzhtmvb+2F+T2iocAgSiQ1gp9Q
eVX4HaRamkQFRndGhNEAlJGD9wNyQsDjifTHUdqxGm2f+O55v6eyB3zChiTJFJHd
Xe3ykmiqoSEEuid793pYqJzcH1ns/YX5A2XqGbwmu8uAUc4iHz+fcVXBe/I/D+Jp
qf6MpbVxAzUAlsYpvUgwdQjTga4s9vpyy8xROEMsesAbtjSZ0xypa1q6okc3qWq0
0FbIr4K/yT9SoLpiB68RTrQ2bcjCt4mt2wFyuSrQ5r/75n6vAudAEwZHI/I+KJeb
wBbpCXvslvzZ+/3DwdrcGeI6YAwJGyVExmL15d0BfN0pX16YG5T7WpVyk1TXTeqP
kr7pJ1ewq6UrVtIegVAiFARWIl/UCvNbK9Th8vzx6Pbu7a389hhNRRH0c/qxrlM2
EO0yAeCT0EXfqSpgBDyH7qA7ym23+iEaS1VNhs8ex7RB0NvIk9Qykp4qwAgjmPJG
Vy+IJKiKtlrdznU5PWJYJcb4yZ48efTSRmFnVNNZPJZtcEEZow2MinZUZJgfb/sJ
DXmE3iCxtdcInYGLTuB9kc1V0eq8YPnj66uFWQc6EElbag+AA1kLpmHqWalaeqgH
bhRfC2kBWYqoG3JPNcxFMSAbJAuQjE3n12QN41XlK5+UsDJ/s/7K6uwgzI//rCQ1
v+gpFKe/9gWoKE95PHHaDUNV6GjfDsjgpYMxc/Tnn/T7+pM/ssAI0Ls2tKr+dSIc
0qJ7Jnmf+fCBX3MqgVu11BGH121agVS/3Z5lUG6hx5JSPVKW68GebL6Cz4haswVR
EPNgA4IibQwiTE9MEYO1eoVZvasBI4f+W/8GFpWk/pOR+W0xkdGUBG7qU75dc5v1
ouL1ZWLmmGYqZdFpqmkT85TpTjZoi30e5elyY3VP1Zh2v8k3i4EVi8BzTgQLWnlA
WIdNSDX1i+Vd+vDsO5zl3Un6DJYsLDjrTt+usrwwRno8XfLiy6HlXvcklCB+JZy1
GDuhBbDsFQ153FmeBczzzlY1gvA6dUHlXDwFfiBdGCuCkUfe/XbGwW0WvrQFud7a
R/PbELPkvfRJrN9RGCyR6YK8hoBPRzFI0AFupVQydSS7Z6J5Rpieif9EHsPp3B+c
PUWLZIUqU0K0Bwu6Gu9Fp3ufsJT9cQ/OcWvzlVIAswxY8J7GL2rsR+ddz4LIaKrr
k9Vm2bQ1ynmykPPd1Lz2iTgRRk5fWHPpdPIV+LKZ6FMEz1v5tLR94eYaLkc+ZxkH
WFOCRQT5OpaYTwC8bLEh9xNTUpgh51VWZBNnA+LuGDW1FBCff3xLP53aYAhaPAVp
UQtl5M4EBrn9yfnFtZY+gpTW7buQAlz5qVp22AA08NuaeR7t/T26PJPyX3K6waC+
FiBzlo5MNTl0O4amOPFUwaWh/V0ylouf4sZN8eVWxJW+DpAYCUfPYgX3QE7nVRbb
MmEiKVcyqsWITYSUrSRDIwX6r8PMQrLIzk/kOVHwEXsa14og/fyEPZBTx7xcTj80
aaAh6R+QAJN1E0TUpOFrndFOJaYSIG65M+YxQiazyALRx9RTitNQuay2QepZLUET
DJLCbCoeixX7thKhYiBBPqBBgSq7BGY+wqLD3l/GjRVZ49xpl2eCwYt7Ypa8CW3D
J/+rEpUPy+h3uz9zUcLq3wi2dkvimbx5lFedcHeykXjfH5RrZZ9zQoLw5boTFUcH
3uj1KYh8iQqXtS9gsBK6W0U6QvX9w6FV9rMsC6I9ruc+3rhehHQ3uv+ZWrr6sZaL
MrLk5juELgK1n+adXOVYvdagq5byf7VwhQS94uyfiifhIklxKfKQN6L0EG1M93Gs
tj3ggq849J8JjLrnafGMwJ849LibH63PCeAbqjFliDxiye/IITxpIoaXCH5oFPuR
I9mmI54M2o0rVSPkHNrLz3oES+wV0C8zR0NCVyXKjhWcuLwOhC/6dvpTfDGabFix
JDK2VGDTtb43jdIHEMgUryPGERScgfLs7LYh1JgiBwwIbJYx7zhuYLRbBS9IGAj/
Z4vyEPK5SxRUS7v/ET+youFOCW3J+/xwbFxbYPolvoMYDNj6p4m7iOaJcT7RqEDi
WNh+KaJ3bykgAFL86ROjudKBg8YDyAL5wIpf92ykU3mXfehrl/1VYA3G9E2F3HUo
bGC7iSY4smkcVJTl9wKfeYzTv9sZuqmOaf0z1Q2LhRNYppO1blkmgK4Y/6ob/wOU
grwJjo5dG4F1fj3kp6Gv7qQAch6PPSrsniJ6GSMHKEYegV/EnCGcm3918ytvwEja
X1tg7yzoW1uAT4rhQtB8MdbzIvXaI/9lHNP4yyg7wB2/f6TIQVixHYId2HEjNiKj
4af/LurZrDVThmvKD3gr0dDWrmOKz+JsqabOacmIX7gdYTPseilhA54jKen8QoZt
EC6ZN/Kx2LRQGjZQbhdThlgZJk8tlOgCWRAZ67jW2DmNYWhGrOEC69G+QGc9VCTw
RGAFX0EvEBISkPZCw9I3ymbJg3KWEC+bj632e3fkVtaI6xZT2VGHPs2idDFydUQ1
czEquNjE3me7+DQAVcf3uaPvg8/ZI+HtB/kUaj3nyI3wAiMvMXMQkTNP88e0Eki8
JtJtb3NgMmHowM+He7vUMd/kwyzS+irUuWIPB0C8cU5Z4SNH2KVrRsKK2sUYAm1W
Z7yLqJUoMrPpXoYiRDbm8mzKZsNwoiRdYvYP14Mr4m/A3fOmSZcSPV6vhr2L90Tt
I4WIDdQdiVPMkllkf18cBNcU3p12BTbeMRsYY43+Nm+BEhNtar4wbmDgiP19xFVa
g6cI+tLUbO++KaTDeSktFN7n8oPC9Y4PSBst6lLE8DoEG8YGEx1MgKBs9/LccEf4
yQHOFWI/9f4GvI4eHNotMmt1rEZ0Z3rCGw7Ijxnkm1ruEEoQkKWnBL6a1apASFJu
T6NHDiAzEiSe1B8+G/oIXAD5cfntBxGD7v6dT+mrTm8hmp74PJEhj4wkAB9K51A1
IucbzfyoiPoeoeoxSQN8FqVVIwl2f5Wy1uaOIff2SnjMsc9fiFW2s3SmUzcEapzm
mLWBHpxuujeCE88gyIHwNY6fflS2IBpZrpYw9IePQysnAkTJ2cDWfiCs0rXMZXF3
u9kan/R4elMpmpjyRwUyKZ9onV3xb7Rj9KqHmJhyodCJk7LKBmafAUThCPYrebjl
+EWQW928zAA96ziNzxcwLCXHXKlE/a1eTva1/V6233Mur9+j71708JmVzZCOdUBB
CQxRtBem8On7lL6e5MXbqz0bnoauNmCEzm9vGikzq2HEgHNpmgX5/oGcB05mLVFm
HX43csBPlKi356LyYGyNGSFS++1LY2Xp5ADdqiXF2/qSwLs4TZy6w9POBP8sKSyO
pzpcrvXQx4BXwbhj7rhF6hzlVGQ02/wMFruBViEbvPqaEwPgMVbK+bj/KJNMmWRS
VXXcvbbeNnkQLOXRwlXVo+46T1ulzjplEx0x58pFQNQD5MfjhCWaE9KAYfog8enn
3NwtqOtbeOv7YW3tOOtC9oThGUNd44d/nMbR/pJ6cqQtDdASK6W/yCYoH9dwXKcH
sb0RrhZMakEj1Jjb2ZSZ50bRCTasvWDx21ZzxNK5UoGF5lzNFvIpYxtNpvK3QPgx
PO0XPApL0JTfwojvns7kcbdks2MIgLVmp29aIYi1CILBQ73/ZINK2GKtjp6vUIhJ
r7HcnFcqY/TzuFpNs+0D0hg/2yL1rWaRVG5HcWi4TiEoL75e1stdt2Mg8EhreSLf
DFUE9V/a0c5bq0OB+kwOB7B1dDE6W7IhQXKfaJ2TIORoYhbtFK4Ugibyu8lsRjbs
LoX8Asz4VIskX2YIo5JbwPqP5it7mEVrg5JjV6A6ltSe0GbZP/AH1dZwr9L6Xs1N
ilbHKn5KMSzSK/GS/ysrWm+SU02FpArgT/Y+NAktrLkDc05Md9Tbo7vit2N0OPoa
0hwcvlFQ284c77+LJeXJ6khF4nxrAeUE7i/29rL8w3gLrnIpa6FVmvIRxfcyL1Yw
hZEHYDmQQ4U3suRDlWS6XK6IQ5lMmWwc9douqDkSk7iHrybCcC8c78aJMWY9RoSV
UI7xu3Uax3RNN7ECkeH5xumj8Wbpo/yE9lxWSbpcLd1ILmPJE7gvBjDQd8dX+ir7
a+TE2aZY92QYE+nTpO8Dof+LQ3ncLPbIFJ+g/2+/FGC4J3/Ps9G7zZ0OWRNiK6Xu
VAuF6pyfnEgjAOWJCJYxzrATnLspMB3G+x7Mw8jPdPVOV9LC2X+WMbAB6IHrtZaA
3JIiBIM/OnSMO5cI9FzckRdBpRn1DP9pvUQTraXIhdAGNrEsZ3TTRaBaWzd5Nwn1
5LwqReJ4k1I0Fl4id8LSsh38jQ7LS8nAKiYwOA8D2LK9RG8C+vkoR0tfug7phvnk
8wPpRTcdOw6iPVtm1JtBsxXzKoi16kYu0IKPynhm8T8P5j7AFK0Sm/xYzyIB98qb
+Zwq4JMuzCPdXthtamgUd25ZvTkCUWVDPh5XwVOs6+cCwZ2uL+IUbmxCGne5Ymmx
96OVQh0CPS9zq1e57/lEy4GC95UqEs/2/pgTNs0Jido8bU1hx1pL59GMRf6/zrxs
ELb1zHpxTJT2Nfendd2kEnef9ZUiBB6Yquvvf+XKUjGLCOvF69fqLlygaaE4URFl
n2f4lbwoYr/FNreOtj5l1ls7Lg/3ixwQ5pXZooA6/8cqJSRVlOsl5YzjvFbTv+4/
M3MLOpI71rJcUovTCJwHxHSI62CATnLNYrxK7yYfYBFHwP2jBVjlkb/b82citSN0
K2lFLh4eSvLNwqjN39nr14F/qrir6P75p5DueWgBg8UOG9qpxcq45x6J+TS231xH
gGVSSTh21R7TeNdoHplQc+PHD9INniwpqVUYs0+pxUiIm2AxhtW6goTyd7EDY0h0
2DW7LISUU11rFAmpCDyRsRE157Gxr27ZL7qNB8Yi/iIgZGlF+6YjUF/PGhTtgd36
tJUfxoIU4N+swq5wZkI9nj4gI2liFn/hDlgQ8tlBFe9E4tRkAs1qFjW/OgpQ4AuB
dWpmVq6qUC7851p+HJ0ZAQoGEhVrg4lGlUYltC/dN9fVdn7JeKVfJ+TbGLceibka
/CtXBpdvzDdIDj3+p786SmSV7aSuyjHEJXgX+UeQkVl+5gk29Vo3e+4qEi2r7Xr9
1ZmfkwuoThemai4lm+WdB/SSLHbXTSVBeC+U0yIXo2OqDY1iOJ/kY7RCXkfqnpMn
cL/JHcK/8mfLOCNyvS53ku+8bPEjS4T6sRk3D3LkW15XYdzoM5Fr8bqaAZ+NXyuP
Wv6pHXycz8Lf4Zkjpzi7oapHMfM6684yXnn7ibzzCQCrXcoyRqkJG9S/aVyd+f9D
HImRkdPN71hJCYo8zlDR5q175jrtxBLbbwyafB+0Guoakxh87Us3WYBHc8dLrsbI
ayTNoYpuisqTGtRZCPbL5uYvmu4ajHT28M1uP9uApNpwBwv+2L6Aghq23CSEWct0
8mJJ04UQ34qA5cSCsp07snVAHxCmmD+MB3uxGuMZX27KBwoQg0A3XsuVdmuhIsaR
dl5ljOCgalljISFdZeLWHsftWyPFaqSDXAjjvUDiQEmfT7FDJVT8ekNTPw0gjXIJ
0s4ha9OQzmvGLdsT9CfVJ9ToZxxfOJAQPeY6vs163GSGz+OQGknugPyFb8i7/eOt
iHnPnKjzzqRVHSGdVylFW+BP1OUrzxSXYPYDVGG2hMgkscPMguAvXcvRjiKdD2wn
vKh6vKvduy1L4gGrbLabjnl86nQRDH8ov+gbNjAjrmAJhP/z41zre5eM1H/GZHRJ
rJXqztK84kbr5BU3FZnjTE++gQhhCVu97FXLmiA50dkTj3JCd0/SfviHGM2UA1AC
caIcxW3U9AMlC8j12HbFVVbFY7r2dvXYhotfmwCj1R3H+/LeKmEaFLGxij7+RpMr
aI+tRinJi6SxuBcg3v6VvPik2j8lMRAmoSsjoMi7UT4yF9GhOecO4ZSZJ50OxUjK
lTUteE+CFuPvCxrLn/H+GAoTBIZqsQDXtXEBIZ9FqVP1NJeZewoayLupTujsEjaQ
taN/dHwjg/JGbVIMxex18u5XMVa24rZEvaQyC93GLO93Yt1wjsYfXRKUCCSyA8K8
lAludsvtsYid8KvJBMG0boHzX85iTZreje1DxmHfOwL+U8eGx/kXSN2bbpMLd8mG
NQxb7QxDok58ghnEA146sS8dzT7X36/5cEW/htEeZuJs2Nta2rJ4QGwK824RENP9
wn5Igf26vMeZxv7KyLzadH3p4DjDyXlFqN4zi+QVfgCuF+et1wMeFruHGlGSXldS
adDIWxUx+bgxDqnnYYj0GfJe+DizGJnFU/btmNXWhFQWHnnJojsPcOuER+DwzQNo
`protect END_PROTECTED
