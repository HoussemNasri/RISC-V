`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5LtaGc+x601QU1YJ3fk4YDjVwtcUu6Qv7W/Rq8HHGZCHRnksm/QcAL77Fn+BTmTO
ECcFxSe79AYwbYZLk/Jabvm98fG5BQ+U83REy6EERU/CokHyqcHM1gJwVQ/jiVlE
agtFL0OCtMDNgnMGhjTze0ZfFtoYnAWadtCGt9PLJ3A6GVPjFUW6sN/Hef/Yj+4N
MpgRCrwmXp/dVN7ngNQAyRrDBiBBRcGVuA4xDdz6ttr1QprlNWaOm8+4imsWODiA
vAX6VtRf6Bbow2W/Vi6PvbeB0Hg/DjHbDiULCHYsFNhA+d8FWI/dgecr49m2VxAa
sEw+RREbwr70xayYCUm5HiwXC5NuzuCu6rq6O2zQ+j1f8WbLNLIFo5L5aXUroCo2
1FAJxFfX4ccq3WezB1du0hwOO7B2CbrDMIgOZIplWyeR/hfz69uM7Dh5nGUix6WQ
4tXcLiQxSUcpBQZzuzhxJ9excAlr2VBL0vFFxdwG6oyJhqV3nAjHeeU7JYViQyEj
Qfd2Vg+UMf2y0Fr/gc9PJ8k1MxJzjeFJzicJ4MTjilXsSUkXmEXlfGsOzbVPYpaH
j3pae0tGF4PYRzHintdcuX20V2xR3NvFfIm85cjkUUSJz6IwC56lFyhcuoQk4VTt
mn94rvlZQFL2xWiEmlNrKeLjdnu80cV7zue7cYLDWrUHqFxC3tP7W7RD/3NnRUw3
x1m6NXdaarb7sngfEtL/JYBMVuGcYjSub9rot1Z/tee7ZazRp1DcHElUAa0CTMWX
Hx5mN7LONlTw8zxi38zG0OUELa0m3nKfnbnNUmEl4+Z59rWzF6XHuSmAsMFbhuaT
PQOsORkAKsi4uiiKN6772XpCHG7TCjexBGiWOSMOePGPpsTlibq883tTA6+K4RXf
4y6bINLf2AnahuCOJcNfzfzrQlhyvQlE7QI9VLarW3AqYB13afxb8iDzDgD9lJYX
1bkEeV9Q0KV4z6MnqKAroHh3m1BYQ2glCPC5lwVWCQ3ivFQDfp4pql88hjMXLKuM
kM+85vDkG6gxgVoLCj+Zdo1glhq+qy//Vy6CaanHYNd07j5VJVipxc7/M5aVOS4e
MBLg75HwHOSefEE8/cnNTaYWtu48+DXFzU9wPYKIK43u1v+axETO0lU25DMkgfL5
QS9kApQ+6hS4X8yEag17uep2jCDCj/w5GERAZVL2LYBbR8zKN4TBtdCXUhuSDeWy
UtO3mGfF9xXkwWCKerAOjboEAY+9ZPRNmTyAZBZcsonn7fTsZCRwBFrH+ao3OSDd
Khj16wmUJcPysgGetvjBTwd1C4T8F/p98LyqlZD8BAlYOUggQxjCGXvkHp/ZYsgV
Zowk/RvqbsubLZ62Lj/FUNAcQJJoIPf9KGz4ryW9TtYKcJqT0EL4YpsA2+HyRMc8
3nAzPRwvdrNgSkwu2wkFF0nM3BxmDWzykO5pAyA+Tf+mISLUA9zI1shsDyoYZ7yc
v40ixSrfgmwHNXp6szaYQ4EtsMEB7UDv8HgC+htZejftgbyompEjrR7Y/naMODeK
3HBihNkrwhEnp8iTArxNBOscbCNcZ0EGpCXd+RAlxgN0JMBo7/4v3rIBSA+9+zXz
MrmHlIFZ6nMRaDZKytO6W85KpzATnsezowdQQtOdWa95+oGeU1Sj97KYI/4EwUvh
QV5GTDtpM2bSNfeZST9VTk2iTY6aJ+Zx+TgPpFqqRX7H5UO2AEYnHnVk7BfQ7qJj
yFkKWB8LkJ3vt4nEQo1XUGcutd9EdD3K4aVM8VDoyv7sXJRMZR910zT7pP/ISeB0
VqYXHU8RjBPiJA3lWVx9knNS0Rh/FisUY+TlV/YbsNtb8BkzD7DX2IwNAU0lCz0T
35D6HoaV3x5EalPNi34eGM8LRdZpiy/l42hOCLG6x8c/4enH/DGmJccm/l/uVV+H
ZxVIfFZucLOIKen50Jibcc4lRLfAfVPg8dWR3/WtXIsu4BVLHXaVBPb//LJvh/PB
1l90AScIlB0QSIQa02fYkLk6WGiSXC68HkgNB1Phqs4xv/CF6E8V5cQzr9ReOikx
VI4lC4wn5MzGZhlZlrq2Jwi2e0DEh3tcgWKZ3xI7kA2WPQdR7qPGIp7TFUIRsH2n
2SOYFL33GdxC8WLTWrxOH/rwclg3L+z00AuB78PfzZ19jf7WGWE3YoJYK4wbcudv
MkDk8nCQ9kptkvvgfccdOpZdcczdjhZ3ZnhJj8hrM8ZN9de32JMmrHyLgYsHOHnq
4AS6XUr4R4PrwTtzE2O/8635Hl/kP+DY25YGtDnBQJ4bST03miHXlPvPUKlcdo29
XI9blgS6oFLVOdd2NAQmuahTiFYsdPg0ZXcRinGgzF3aqx1XVFteUGsmKePkBEsn
jWXwjYlXxlkjsO5Q7mEHgEmJtobg/mPiLfHoJAc4RsPSI4jLTPzp0CCIsIxZOP7x
glRyvERpFktWQiGv1lK6OmkpkRsfCaiSsKVPiEE1Kn2C4kcXC4wbZtb4FXVJ1Q2x
C/qrw8xUmYCGB07SeUvyPraqgpkjO9ljE0Z3WGNvhUXWRF/xCPI9HQ3NUKTl2sfs
vP+G5Oz0D18drfo9uags7BSnDHZheHm7MWnIlhSSYKbOzIIOgW2TXxcQeypeSLDC
LEmDE1riKkCC3d7r7KnYy01KfQscp9AnLcwevnEuJmg0mKhoxf1yr5LRPwn/UteQ
B3M5ZnimAvtjHg1rXPQiakq3Y2jvL0qKQZhiKKIunwfuZCY23q62gkgjndXJKQg7
MBv1hUifgFgaStJ9ynu8qQJ1pDSYjuBg5mwfHtGx3C9A7pz3MZPXho+5SnyesvZN
cdex6mu9CAvfAvEdAlahDJkhX1eH1TZC4eNajyIJiIXp+fM90QA9E+ezz41ppbWb
Af5wb4+wEH0En6cZCLV8Ee1pJvizaeausGf97EOBoDc=
`protect END_PROTECTED
