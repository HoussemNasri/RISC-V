`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KehjJ8w/PVhLYy96PLQkzvMWXwyzisLtJyWdqVUOFF0473btovPXGAKy4lFjiP7Q
IZLaZ+pgSCMRGrAH42giUEjn40tS8I1Fw4bL9wNbgiFS7x8S5uLBT4wVxLmdCoOs
dPraTwKcRJNxbkLtmMyOOqfuLQJTMiKpwf0wC0JBfMRSrIHFaksavnmSmd8+GvCT
GwB9Ux4+bygUxjs/RzlIiGnPfFtLihqgaDATFeRvlfTDZb8NxZxD1XZOcKefWW4P
wgO4lJY3W1pFrGejswelpMn9UvtuAkq87/8pXPr8eBQeDW0LMVCPMrmgaLen/9mC
CKFkAxs2Vx/36i/EksWu0Bh4sPNXcING6TXuuF1gr1XayAxwt62ArAvQExagR01L
v/Blpm41QedyX0+YbulaCrGPcPAaWD7dMw1uhuyoFMp/ZnE4vvWHLtT/VZIfvLHS
LaBGnIWOZpd4di8yV8XhALKHHX/bD45UDuES3s2YJkU0qgdTmXQyMDzHBiM40ngR
ARcH84yG7sDC/IavOu7JCAtqOUdBdQoXyzuVNPvHkN2HUxprmueJY4UjIrftQGGr
nWjXXlSPETdBavTAtBXEdgqVqHCKpdmWa897CONo3OT14xU5pNjEgPw8S7UpHXpl
uwI5/5LSV0pqVNduKaz1nWfCMy3VY1Bu/4VoZV0ngi9Y6vw5Uq2uR0lF0jahDYdG
7NF1FeI3WLm2mbXBkUJNkvBV/Nnsio3U2UGnuAjqfTbNlm/tcG8Sw2zfbBT0RQFO
JfLICnx+J/Hf2wMHICMRTrsXzfSLRkq0HvqtH/1Eq5aDmmfbaxGQbU/vqvqKQ7JG
Qu5BwTnz+7qdC/xN6nDPEMeNhZF1bTtT0stTd+QeGCP7WTMkMd+hTDmXYAOFIZID
fj0Ieu51vjtVLSDZTWju173ZHg4sNvYANsRjrY2wjhQl5J8N03WGC6KvvLZElSPb
jmZKovcCHcNNVZUFRo2qOOvOnVNWHxMw6oZlgg1vtmu+KkTZqwNmCzcGicE2IMKh
VKTxJvzVGUCv7FsVUtlTd/f+gZB4hrcgGBUPqsJHC7I+K3EEvN7FrTLPhHrLSmrV
VMro7OoI+GQXeuQgHq3+yy9/fbyxjpA3Z0BMq0jK46GaIIdtf2mZ0duZSZIXmi8q
eXBsSpZVUEfAOnqIa9SfD/oBtMsl1A2buSbvOrRIPgYXrMyKOWD2tQcGn+WadiML
2C87tGy9w2Ww1q6FNhJ7FikS3YWxsHAdEgiYZS/TPa14JIoFCCqD9N6o7gZ4f8Fm
QlABdusyC5bCANNW0Gajby0QgbDrCn7An5ORcrR6fLQpbBlYSwpsomdAR8RMNCMD
9xfi8vt3XB/FDi5j5Q7nsPO3JSTcIrp+kKWED8ttuMUUuqaQo1YKnpy9UoYx46Gu
/Vqsh8zS79kOUEXV/1yOXPXjLZqATeQA98rEaviufCOWNkPcN0bm/2WRXmv7ruUV
1vk31ss8S6oiI90/5HXVM1R3GApjBCWVGNPKnx1wvpGIlslpQB4DXkj9C10Cr5cA
jpVoqNDKxy1SrbWsJNRKnt6SbqmvaknM0qDSNHPxOOcaT24zloS2KQ0q/SWsvM99
hUx2Qkkh/xjFncVsMltCum8WNRfkyh8a4RcLGshJcD/YVXEDsT1g0QbhszHvzfxr
7aKbcYyjSiFmMMtsUwGzKQHIEIBvIf3dOa+TaM7K1S04FrEshBgLGHa5WTlNTqsz
US6Y0IJZexmzMmUlQ3aAFNn283m4qLQkMvd41JctXbXvV0PlcI6yi8+eOwrEIXUd
wkU2AxmKCvvU02Yr6sl7xqHJzLx53VMu6iS0tUWm4QqI7abB5YB1/G+k31mNBKtR
S1WXf98zxj1mm/NF+nW+4RthSOZkISeTF3piS5MfdTent2WePEegk4yG1Kg0YokT
Bcw/dh1A148dPYsrfm8oB5gnDOP8Nlkc3JveXk0zTKUVtyUAnlm7aAd+v9u15L//
e0awHD2sdaWJNZ26xCPADwqG/55PQWmPtxBrP8lDSnvrgfqL2ESNG9g3vprROTcl
e8b6ksY/BYRmcwywp/VtLdeupx/VUY7FUBI3QSgOhGmTpV+GanBqUxmzOGNdeYka
eJWYv0Kj1C2WFIVUtAsMJzzhJ2bEDafxnofDqtmQ9tOax5mPutOGjHujiS54lJFB
uaK73ZUOwA/PnghS+MSxliEXJDxcpLAc3RNE4edB1tn4r8FfAf+CGnJV16H1BSFV
Q3HAqspJOIOy2yN86Iq91HiEUmEeTy85wY8lJ8/xt8MYXfO9F1DdjI+E/UVirxgf
8qIrotkx7Mck87mksb6bgzjnLBHosHrwHSmQfcptAQgwzL5Qe0czNzl5gxGt7Ioi
0xlQJYlaa/zxs8MI7BjGnEizPwjkTSRM0BzzPamTm9UcceCDuUdLNkzQnUBfZe/k
QwoBCwSzuzDQjDY5/rHV5ONE8co87Ir9WWGn/o2081r+eXLoC5zvqDqzK93D7Bfa
DaQgJUbnJBaGEVanA1cvsYCufhSqvGuWhcEFiN3I99HZJ7VgMQYMb/dkyTaahaKM
wOsMTrNQaDDPHLG3ZkWFC4f4uMhU99+An5rh2KFGJ00ZzB2n0NJwciOJSgBwdgV4
1m54GgCpnouZ/MX4ru20wDpM094DG3LQyiJ3KjyP47IejmtemaeKKN9ni2PNmw9c
epw660COofWFyXwdezDoUb8gI/93wmHkxq3Im3EzVu3mL/Ki0Joldc6n0/w7IRs3
Zcleo16PyosHXctkL3X2dcdJIMREDlZaPCNBZv9a9GCFCjctKJvHN3j5s2RPWs12
IYqUYqV0X9VeqIW4e77wAnTKMi/FVPnxyRtRw4D8IaH9Pi3rvy8A7hl2G53UAhhR
iKQ9eZYM6HEsYkfsuLmD8JYmX1ggVUC3AaS8BBMOvnpr7XlSfLOfUcOa8SXuj+Cv
tSF2o7Pf/iYkbUobwQIlNjpwYckWLQotI+DdK5GxzX/OneGW057nSS9TcVdUPDfU
lPuGRQ5pz9cuB24aYnSuHWn33KO4hh8AGeKA/SThWnk+xUh66cTWb903dbsTv0aY
h7u5httTmp3o1qLFZd5lyNQKcPuL+ybMO+4VWTc7CpPpX/H7LQqKoIeSe8eNdDFg
j2vsqiWm+xDZnBIB4KlknBamjQFslEH//oB+v8bzNYDBRUTmUyjoweFXmM/G5i8/
gHyq8kUTuJtfDESRKXs7zJxlJz5fiQFQoOnMMGTEoJFruVQHZxzLH3rko8+ud9mb
14ed4Mdsn+65Ov8/elg4N3rJyShmpgefGWcJp88hTa3fTumluABHqe1PhQ7P97Az
/2RC96rVw20zRWuZxi2IkNjOuazqBjFSwj49DV/I8UuwOQvHKJurFMtD0SnvJlfE
fLOml5KdHMcDknJ8ieklsrKJ2CjpWWUGp7aORO17QKb3xisAujfWEGIUhymkI9mG
4HYYrPE0eI6Oj8mYUX58D3pB7XHPByWPvdgS2Xk2bXw3n9oh0N7SMNVdXhDVOis/
06mnj5tEmHkEm+A6mbrbkQ4eNiJ4ofkcsixnfFfj6vnRxP3HG9frJEfV2/6z2YFW
t1lY/bUAGQJhItHDY4/AIwa4ORCE/KSAqLgvHWfTeeroBGG2VqjvdmnO5dSY6vFs
x6ydv2ret5GL5U2m2A8/UsDjqZG/A5+ADsq69E82FWj7b/zkbtMy9Rl+PNEO7S48
GAAWXdPxlS5/fckOzR5qRncjSQmXpCSVSZAIY0ADC+EO7cvT9dMbU+rr2oCxmt55
EDxgw2YVBwLHpeGeAQXSuDvt4I1EDYE/XfOKdjrKjoeawSAhNcWYIEYJ0e3RU25i
AnYToyVjYyydL+xTGf/drdn1byNKW5aBEZKhWIGPTlKr+tVmFJocpd2sX7ZDniVO
b5ksC9zOeuwYQoJo0sqfbH10nIa1v3kpfI26Tyr9KzscQfeVuj6NA/YNqPIsmW9y
5Fmk/famM1sfUxEsdiBNWKM9+WvO/hC7Iz368m4HbFafyRA8enWskjs3EoMG7eH/
knipRv3TnEVQlljU712Dw7BoE5dK0J/Hib1cxXdu5ir59PEVRZ4VU+ThOt4OkG23
aA2qa0hFIac23HR5JITnYzORzxwLPM0l+1/vClZDr/mIW/gLih68cC6vGgCxZkee
EEtLmogD0I0O1O+nagxy0krXE7UHN6G5DcunJbS+mDVPl9hXDA6VDaB2PWFvnmyi
VdyHRtl0vHU2uJ5wWKLier36BnYitLRLVj/4lO+6bCgFVDVoGpUYqboKUQ8PEb6g
yzk0dtfpTReaWRxZ//m2WDP8sH5uVgx6rFU4hOBteu1W1wUVUFuKbOv5eRVSMmOo
mNattguvGWU38w383CTwZDv4AUtIvo7zoBH0E7V+0XhikCQg0jvWGgV34Oai0KJz
MHnNbq/peo65sT7easvyjEOJoPTkxqlRdpmChbnqtNibs5rFc1nJZg4xSBi/Qywa
tCHU8KxKiU0xucW8whHx74zPrZ2HGrHKmrl3L0Z14jmntlSVUBpYCh/OZyIVrAQR
MK6Fr28G4lMScy1qRqHd9gFFKXKFb0Eo08+DawS76BmMSr0y/G3e3id8LfcujPGI
nwie07wJeaIHJOUCalowzlSnKg07YQ/ycT3KX8N+CycmhyS8usNrckw9tp815zVF
FIVa8oaQ5JYUMJ2ARVqAfY4F8YepmFTabGVUzpYxKG0/65Ti61MKmgMtH0yuDG4B
ci0/gaYqhB8s9Xf9yXq7mwYkPRfjXzRCoBe+NMR9Yk7LVTTB1IrLg0fVY9PDFDGo
YuADecdJxLByZs/tObh+C9qQiAWExn4XjWgAcGZUU8eMoZ1aKXa9IXwgAp4HwpK7
+vUyFEgb3LYDjbN20hSI8RdqvGMe3nJ1OqbGHhMbou2Llh4+i6iIzoB9PUbQ8zuY
6Rmprn7sCKf8X5iA19YWUHFlrT/oMk6uThlGFfNYZltKqa9ta8cPy4qfBI4rt24p
QqvKPp5owicqCSBXRmq3CPM1OU1T62/dUaPKtElpj5oEjtLlwfyIfiiZ4BnjGDcb
rW/Y4K2r5r9PFyEklvCxNY/kw0pzXYRz+OhmqQ31vbrGWx5xsCdVfQcZNI5lAdB4
3p9pS9/1Bhb3R8vH8vQhWbVBTnHzRhjasezlTlwWU+p5drQ2iBBXRNA+RUJi+r28
NXhTcXr0mVTI/66U8eToH9JcKfEGHRXOn+sflqqk3JCu8Lx9OsKz2e1yYKKSOOuw
R1qU5xnIQZjNLJrZ1ztHRPzGh4lPye6lEUMbWLjQxjEkrj4K6OY5HQ5M/1QZ7vOF
ofpPzssJ0ACuYLlw7Mimdx5G6VG6rfPoBm4B2m6qgkNrx9g31z0plC7bLgZt6wgY
X68zaSp3LejByB6OW6gznidZ/b9wjvqhqqGCnYvbCxlIF5OoVX3atnIxl+TiZnEn
LmOfVIkj++P+KEtdgdiI1qwJyWNsqE4quG14VDo4Vs5guhBmwXkxK9XHRaEFOXgB
Qn+Msl42+ZPwD/U7qLlEHBKtnkA1/HY+8MnY64V8XoJrlGogPv+UVfXI7PaYr1Hq
MZ4b/BO9aGml89Zdd7pSjjvr2+VhvMBteLYotfNrxo0PPCQG9P3dmMF7g5ScWXMd
zkxIWR2a/7LsfOiaoxFq0r3gXJ3m6khMoOi5lDJ8z73JOnJpy22t7yG5+n1Nx+Xt
5+jfbzt4wtbk5jXr0rpW8Sve87wfCYKxuczeCdoVYXBV7BPTHsopGcpFyG2/n7B0
mt2hapoOvXBaBS+4BqdE9Ka3Ae2L/BDKA+1g9mC6s7AKG4hr+m/P4OURo6LJ7yrG
KppR2w9Tk+UeFMnt5OiuGUoIFxgMAgQhmR/lrH/ssLplbFWW8FP9vZM5SMbTTLTB
Yo/YvAUlJRjHcUf/XWRzf26jiD+76vo+nIFlo2UVzIpwh/LL4RpdCLqXGE627EWz
rUYuWdnHuLUTm43SqIu4h2f2Useq4lysPZ/BTy2AXGq5ll1/PlKur5aoPZl16zDd
P9E36SAgrVMozHVMlX04VD1vAAQvEkEgdEb39IRBhDU978aT7HrNreNgK/cOFgvF
S3ozjDI0CphOON8l/IVWDjnsjx/jqhVG8c3BPHXCmrluOt/288q0ecZNRf3IqfYy
ER59rF8bu+j8+a4C2M8QHSf3xKoZOexkqWa0ubHsPHkcZLUHpD7pWxlogXqQDufw
T4FjulO920xTx3alIecTHcM2s7p1UB2SdbAc39SGj1LlXBv8tto9csAwx4hm7voa
jyBTBKVUED59H0cSBVMMbIxLgKhe3e4ZjI/+HscBTxUEsC1qZOPJUeoMqBl9x1V1
ou2fPHtrxCb3IuuGHiTRbNBgG9iJeDzq6eiELupLdky+OIiIWalzuTXTAnwBkWdC
1MZR6o+AYnsmEUDFiLfKV9Zk+Qplh1L8UvOstQWd9D/3gv2VZVwXkT5CADOcJaNH
n99DX9io2nVRVxhAgkL1H/dppwTJTUWvcyQ+pccw8If/JGWxh6uWFem5G7vd/1Jv
SaeNVIX/f9xLUxaXvg9MQ8dX8yrmngKRpaSqXZ5Ho0x636WY2Z09SKJqOdhe4PGF
ncjWmGFxHyQJWqeHIwnItcNSQ6PprcmtUZc8CZyX0UQ4evd7lgWSphfS4C2ZF/gv
DSnUxtxeP8FfcaU3l5jYhhnKWJEo37GgHTiMQPaOxcq+/+jqSZpqtEh4lW4tI9qR
RrXi+ucUoK6DgqcS2atSXUVBxz2C/i8OAzMuSl05l2DEgZOSHh8EZS8Sprmyh0Z0
wb5Xiv1LS4nannfInJW92YPn805ujVGy4AvSI8iG+x1KfP8wMV3VBen/Taz1NQnZ
C19rCSzahaDYi7t8n8ZvNA7D2wrcY3WzTPufbFALXNlV0ktta78IXAG/7H9Hauqm
YucGRMfxx6+9K1up1znn2qVLr4ZEijeR13BrJjHd3x19SYHVdqElJ9/BKVsbqvlx
YVvtAr2FlnbOcEAfbV3gzWWjmazgtwooSxSHhcZ899+DOxH+tw9gfwY2hQYBpA7x
GGPgkufevWdb7/8WIynZe4q4FJHPHv83cvcizCmRJlhmwyCH4nviKnxoevVTWjRS
Cre4JIdURRUta+UzZDOESGgGVZY5J4LE5qQwfVsQp7rZTiSvNrT9TXHguHNPcc+E
nu6BX8WU6/ed+TF8HTWQqJKzwiMnICf0aKhk4GMT9wLU3kCNIfbm10Agz9PBfs/t
63g4H6ESiJyENnz3/fBJfxNntyfvl0uy6/uPjHHFKqTsD/s6cODel3rAH/jUBKsa
KFUBq86636BKnTIm7b3S8gbXsrXXkrh3cLilxn51C7XgBAA0MFwVxVQs0bTw7OEp
OmigSx+pypC2dnLX1/TUNYeIzE36nMvffEtTgooMEnxtkJlM6EVBFOeZhFmDBBZH
yS7AjwiBkEL7JoxTReBmE3bxngCHUbzbBM9LtKOSpNYhUq3JpYnaDu75fc0WcVzJ
eWck1fCOqEiyhxSaXKSYJOSCZph8fdWt2K13b48DXIGY5saLgwgF5B98jldHVCw9
kNL14DFluq/ZUsucszD+O4aeM/UypTCMkN+tO3MJOk2PlTSt+8x8dfgXyyzXeWcA
6XAKcL00RK04TPRHE7e7ZrgdeTwO0/CI9yLl/OdFqu3DF3mKuQ/9OtG/Rz5b87jW
EREY6rMQWO9CE0yjRZ6yi4VTYlODgXc50eVubGUXjDj4U8GoCd8LyDGGS0Im8dR9
ibaWJ0+IfqCmACz3PGM762JNggcs5ZN0WL8bgP001jsP7A+idj9W79aDjkWl5h+c
DIdm+jjVC4WESfhNHyH4E2MNGYmAArhRV3/1UQLNjUqkxhDsdg4Ax1xCSXiWZ8JU
mfdGNO6JLTwT4Eh6qgzKGN4uyObbQZxe4szFRjEqYmCYanBmSYiu//uAJPg+P09T
HvOVOgkpk4ftAkL/UkTO3++dn40qMr+XOb2jAaxK7hf6sNtv5t2gU1JLBqjLFsoJ
JoMDV7hAGTRzdPmamLopSaO9GYG0PrksvQpwQ3Q3qvnRK0ym/hFYmatpz75WdJKj
rQofF5GeFFD13ig75jDG3+UMMZAm7XXgPiQ9/vOLZIUciodxm3DZMue0eIkK9c87
MUiARKvBLhUmLFSdwkZv1398wTkdQ8oMifROzozi7gvtgkO6+/RWrfFhU9DwFkDx
CsiYTGEb7Bp+Jsq08KdIEghNPkWvCtwC3Q641QTHNNdSnO8XIF838HOatNwNql2d
bXW4OvniRQQd30wmjil3Ian62CKLm36N4GBCZe4zc8VyFi7f5vq+2NAHqZG2p8hn
pF3exMDtK/rJspiMNtJ2svwp8Lfb87NRLyRc4VJB+aySE3K2+/2SBYzVb2f9rqNc
6szMSLHpiSpAy83PpaLNZidsPqClj+tUk6HmaCyNxgCs1y4i0frWiNiFvaNWf1UR
aX513L1ZwPWTFC2UGPt+qwHFeOHSGjE4hMFRiaz4shMU2b0G/stAfC/xiwYSn3bv
6Yvqg4ShnheVfCq07AdLdmMbDVwV6DaCuEvSQbgWLmTBImHILs42YGzDMCCqjOh9
EbI3mI6r3n2lpkQhbQtoLw4a3WMdHyh1Ap8CULNgvYU3uimzdsaioX+4hmRbDqPu
q2GNl3ZGMfEXgwLrLENW5GWRo77abiqYToAvUn9gFs4tRTgGqk2wBkUpRcq+Zie2
Pl3vc2Bm/swJp7dMPOazTjc1JZTT4eG3jxWxzrF/5Riw3I8MStXTWNscAojeM6tS
7V0/26xcegsrwnEBADCQDTRp+pVnrOBYE01BA/W6n9R2RqE8fQOon1KEPKAQiiBe
T/UNZv0NZkzdyr7gejakPBdtVex9VFGTs9TomGRvLKomlmlrHnesdqzJXBPIT3Y/
pt4CN9b5PktoNgEss55WrWtGaH93UFWGsE9cSKaT+JbYPGxvcFpI93Vyt+91FsMD
PlFhwn1TGi+nWlVrd2MrHGgcLKRlOWjVZRk4TxlnYZCKCy4MYmAuwB6MOtkMkIkD
nWCSE1Yvj6ntBvIbJzxPJQw4wz/RR1Eh6Q5tmJoHRoi89oEejD+MbBnDW0vYwtdH
AMzrtDzqFpSf4JtZI74jW0bxh25ZcNoMkPv41NYjCthXIXbQLhC+IvyvmEjXMvlX
s1iEFg5gjIZrZJdOTJYjIgGPuHpqVSWLDGlsAGPUMAeZseDQWwabjCxRWfKEKozM
PJTbxKrKENve7Cvlh7PunaKpA10nv5JPOQsDaehmT51TrodBCAfORSv3tO4FrIfg
GVYb8AEhKhfM/4UVV0M9XfYtbOvePOrgGbmUkjBkxnTSINL9Q9EiRMeeb8fyUHxu
iz87l5Ar6D//ANnWpcBh8Xe4Rv/kE8M4xde+VD/0NQ1scMu5ewFWmMiaBnkvxH+T
fvcQn9gKNSR7KBpCM/d3HTm04S2dkncVN+VOtrbV7esreOu7Jg133IP++WwMmB8w
UlCD+Q+UZapjPz9quidzg7nBtCIMUyY8+vb+4htytRmDS/5lUEDrFBLqH9PdWSlh
skS6CSH1bxeDXReLPzrjmhb9lxT3FY4mkv0BvhngaA4Ve6j3lZDj/ZhM1yuWZNX4
QUBtJ76nnTbSlYoyt0S2KzerYp02gUxJ7IJclX7WDC7epc6vwqg7ibkbsNzbaDCb
NXsGBZ49NCPddzh9junelUZpw/zlmctSbe1k/yxoMmw50j2td0Qkrf7Yxyv7ee2u
Y7IjZZVS0Xl6UkIX53pBUxP/CYZhXCbKGTKMbn/YQvieKMabEXXDfGl8jZu44ryx
wfwlbGU1wU1CD5QycXRkkOnq7ZNdRT8Twtmgqj3BQ/5+8QLsVTRG2voX+pbNVCub
J2RrL4BcrXxwak9Xm/eruEztiiAfp85btveTBSx/5ADVXbSp0zMJkkpB9QPjI8c1
PM822q9KDSKk6KQh10kCOVLITx/ayFEJx3ll4iAamKYDEzGlUbDF7oxwfAkpj0wB
VJKPtThJaxPKzGdFv/dlkjxcdo5CoO26yN7U/OESXrFKiRk/qDh22xnsjF2KzODf
ihmUeOPLenUbha/OL4tsZ1t9gw6kCYHuQbAywrpK6AEOKhOeUpyuUj2eQT/AbFqJ
ZdYJPEw1z2GNPpmCtEajGr3OYL2drGtlDQxgBjqiOwpER3e1bLMGA4/68uNZDfPh
iJQYBvrHrLDyqR/pbJ2DMHLFolt4ZA+gNRqvyZGR1D2hURIETNDfQW+R3BeRD31J
lrfYYEQ2BmhTN7B+2rUCkuh1HTGM4d09hDH8bDZx0ywg4JDAapDtTmgnx7lU9z5v
FFH4JSw422WIzACfJGr7icBuCdtUVYw4LEQjUyGZsnKpuvahkHQo9D7GRsZerEC1
fke4fOxqgK5F4vFLuKOKD+zYaurNgGlcig3kIQYrq5CgQFirXedwIYJtZA/HlB4l
TVbaNv0EOjPSAqlZW/uM877gLOFti2L8CTO1iSRmYiGXhx/fx88HsFuQsvpvqBn2
A4+U1cBDF3KJR7duy4nO6ujeTNR5bfH9qIKN6iCoVZaijmpuwwDQEkk6KZqayHAx
LeW9jxQsUxPGfPcRshK9BwUYv3tAq7kscHt+sJNHGOC7VXY6PZ4j0wlomcNG0W6H
lh2C2CUvI+ze80pOkhqVOYswHrdQErq5c8VnZ5zrD2Y453nwhwiDgEXERZrOFBhz
QdcI1l8WaL4Z1Dme6Yz8GKWU0SKzAdz8w6O8aeum4oELWFlGlBhcWcIXyvf2MMGa
7o9vhN3xkIyXS1PAvs2haDYAgi25ZoMHqBmZ2f+a4Di4pMyoIZ4w968NOWwLQRMo
i2o6tHi4fet1zXTVuJB6tyOrK7itfNjsdIlqAXnJg+ZMm7nEl5TC9H9ouDCo1/ab
iedrgZ8K6f3fF8LrrIop//w03bNxxhH2Al7XebmNL+ZMWNGJcO6w07vQfqOG4fIO
UebRvsj+L5RKKLB5m0qrziH6WodDGBiHcV4DJY7APX0OubtJgF1eyDCmNNGZxDkx
GGbU0O7QtbmakNK8QWMOFUqDdfY0PMon+mOaSr19G88AczmqIcnyc3CZmIlZnTcY
ThGakqi1CR+bYt/sso93bZs+Jnm+0R+J5sr9ojfzE6mRX/sjISFiGzlHY1eRAlEZ
wvsQJ8JXvOEqdgisFV0CW7k4styAyzvQBDrF5T5Iagx+nzfXU18BYVeSBwAuAqiQ
G/Q5vwlww1vbdDrvFwj8tGQ1+4Vzem/MwP/EaSOCx6hmh5mKyKhIfj4EiDl8gCzV
hqfllEaem2HANjDLQOx+4kZFSniOLLO9YGbPr5qMsuhlCZDIMm7OknlrhyN99r5s
KrXArwJaCKDSpoKciCKQ3cQnNrjb72pOa+Q8qx5IX35Z8p56tXsSh739HblaYJXP
Z+1dgk7R3noVkKRRIxKdAUltWy4Y+PeasyJ+Or8B0tzauGBQa4eeizH+KbcmZ1DS
TPaOaVwO7l+rujghjn2IWmJYSZXjeLCmvGQXA2DYUrs6ensKL9CGcd6Ir1zblktU
0szoCZHQ4ws9WrVHW+8gqEk6hxo1xGVnc/0CJ5iUbb+r1i+e0fO+vyOi/wF9YS/h
gJzMtGnduT+AapgcYlvOdQOnc20sWCME+p0uWBHas0JwVGU4tPQb1lAj96EXQYVe
bCt+4qz7Re00INTdDjOBtjjVaQrD+CNwOrV9eI6va+LUgTujXbapJej/+IgPiFVR
B20ZPzCGKuamu6pXGfqlL/KBH7kYzBPShKPShzSgZtLDaMLemEtxRY9aEPOgitJq
fB4kWel0adlK3N+3mhtFgrMPCiwUCYf3WzFII0PCjXVERPsrwIvXA93C9zCkB5fJ
TMaqIfLvAiorBLlPJjGs4CiSlBvc5UiDhwOqlaUK7TWj9qMY/SlTD2CHMBipKons
njlDfZzGG6rfweb+W6qN4Ax+i7x9abpdjKlx+bVwmB76yIwMDhsICiIPX0Doi5cT
HvwNlx6DPqqH86fxjnyaEILUXBNNEBPXlIcF59aI8YyFWy4BbBOQyQYoQR4V9qfv
iOGkEOfE0gZnLnnz4mFfqGiA4DAxsSe5xWKazaK2slkSg/9Z7PhUDzjsuK/B4yOT
fjERhzfiWfphVSdDdzul7OteQQpLgkuMmruGeVdUKmYHNinWwLzaTekGc5NwxJlN
XXUA9xvBElCaJPUG4f2udDmXNsndeMvEaLza7ISMa+1pzyVM0bV1xT/CEKB6Buek
up3Qqq3sVrrQJFsYWYD3XIpXZIk59Z6VbAcm8S0WjQk9/A7ruu1MdZK8eghwEgKj
IyKo5OwwtNuixy/LraHacp0kDno8i4c3krH6RwZLAtsFEKwEmRfSctjDdaUMJLrP
/sA6CTBlvqD9Tn6BxHXvZ2L4cxNibuZSmU8W0JXHJk9H+cgh+iyDf5QscE0JsCRf
zxafu3hJrjUy4HSeY45VUM6ZOCqLT2G68qX6WClOfLweHQoIgi3n2nEqx/0iyKRk
hpVlhJlwUPnzMeHuoiE61nz/Bl8DIXU//p6luoRrWVtIVEYzgbWJfLFt93ruUjY7
epywXmu08yNlcMaa+T7hkl42s0h2FgSbR9iiIWYBjSk0DNx5DkG4boUOVXgIMeo3
LIRHyCGhyZ5GGogZx4jm1RhqOiUZhRFliMc1/ShBS1dCWc5beKpUNWih53UFnPna
FtO3g2IlgH/JaHoOeVac1g==
`protect END_PROTECTED
