`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iE7Dt/6jNzOr51bl3rsEhcJPylM7fXE/i2J3M5yLNw6iuknfFhMJL8CPPRyTngrV
Ivl7HGK0eucYLuIXCMH+RDKsVe3J9thlW/ZS2F6f5J/K9iOQjRndrnjnHmZbwcdN
2i0p/24n+Rrwrc6jySjxu2JQNWSvC0iC9tnQ0gd0w8OoD8FYUDohmSc4mexAJVnJ
po/Ng2WsX4BBr2VdgE4gs+ch8bL0x68GYJ+dYv2I5OiSv3OkXC+jiy68BH2wfrQV
S5SrNjQe2pORwptm1Ni8jjyeUy7VZ+Wcn5TWSCXGMxvAPYMydzDk5XhZrJvUQQPl
OxsU9Xo+Qo8gBhBrs4MIae3/mvjJe7d/JQ2nL8ZG4MwizvTCc0/twNNZlIkbiIPj
jQsvWJer06hubwHoeXJ/yAHEBwUGVIQRzz6BySxjbL9Y6RRgiPxec+wSn0eLjTM7
bM8sh608S6aUiRPIbtVzBZBXfZP9VqEoVZvUVUl1h2OMgH5oqL4OV7qm17XtUgJ9
VOc326ceR7rRwdMoZiDC1rwmCqWwByJ03bEjBWl98Q37GrD2oNJ5WD1fMq0B7lX7
urYY+Z0hd8t0Kz5xLF7knN9upnZjTMErEPIu1h1kmX0ylDlhhVC2SGKEIXTuHW2U
Ed/Nx9gBeUnrEtW+N+lAWESYy6Eb/NdqoBP1YuFscW1kQ/G3PSHIc6W869UIUIp0
SaRRof4ZiohyLJsgC8VxygLUkuJ7pfgyBxVcD3DiXZ3s6r8UkTFOSQVZNz3N6ipn
iKbui8f+adAowAc+51UH2bly8m/vAGU++xdfnV5LPlDRnSMlBTCL42h5DRnyXQJ+
NWhzZ17nAq+PJ18lRwNTSS/KeLvRd7NI4SFb7ITcqfw=
`protect END_PROTECTED
