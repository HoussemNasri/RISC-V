`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98+ouEY7zQ9GAmoGiYq0ZdMFbN2ADJZzYwaCZL8HIp7VJEHW9CvXPLeto6Lok5gy
k8B2aKDOnnwn3D6Eis0z14of2Chmz82QxRfNIIofn+RFhj/to3BV4WtLfYlcJ1Y5
w/dKGQ+1T8h62CLlYJMF4aezYTWn0iWwctQSS21eyOGbd1bR2+LJhZ27afoMOF60
oNd3GrJS41IoVV987jcXYZtccbEsVxlK2mz/RVi8AdWOpzDZb+wakdFoVjQC702q
BQB1wQQXJZb11YwDaJ9ojNACpW4zs/1hfcamGd5mNT+cvDyzSk6cQkStH8R3v/dG
xYLB2LRSlrp03LD3x7t9lS0J0OIW4c7E3T1ttwuEKHcQCDIx6I55+2bO4jke6Qqy
lfWeoanrdWMX7OUgssulmVtPL4WgkKB9D3vnPh/jL420L9PUKOws6bwNJN/zwiGZ
KrZoLPxR7KE5ZHpat3Xd1AppxLa0miPTmUu8QW1tLFKcqteIJPTqPcQPXmABOfOg
2ZmWFA1RtvB2bMc55PUEYY/NgepN3bA1h4FWK/5/LY0LH7NiGwcql6WCVgWlII1e
TxyVCyDJMroazs0MNhKSS2wJC5JL3R3RKYTgW9fP6/I1UoErfYUg3bOutmpwgnYz
X0h5F53Tp2xr22xt44oQW7e23qf7G4UT+Xlz2yvFo85bWpomUff1nsKKfAHvNuLY
WLad4Ku1kilcIRgnkEiiT48y+vsH26//J2UTKtXOvqeaUIs3T0kpyeoRxXDi0FlZ
LlDtVNorDlyVYG5comOvu4KyB3xMmSF/HpQDf1xe6Lcbex9AzTHJLkKInLHFfelD
vbw8f3a05vkXhvtZUEdyjBUG2aafDrlXXDC9hKbAOAZG1Kk2u4efUiB2Bh4bYZBl
k5Qc2BpW7Yexyr5rkNvvr5I9UExPBD+kNawgPlJqM+QNiQ4odjim3LbugFeGOhFN
qcbNlpDka9GSRGlRCZ2mwwNufx6PkVY/ZL7aGeX67sZ/Gi599nESoXO/NRqtKmYg
QZZYgIqBfwMGobiO2ybkEDx3i/V0EGRGmW72GJtdXDKCSPc7gZrXsdCJuOI5yGYJ
mIYV9aCT9r6xMWtZlC7VmyUmpkHtU6pKO8pkA2gRW5qHniBFezlAl7gmASOPhqiz
G5GZMJLpFEFMDhp1mN7nn8xGGZwzeU8zd5c9pxmJM2Io/o+aoy/3nvjyC3dAiZ2M
nv2MJo2+riqGJNANpBB7WB3kTi8E+iOe4KFTs9E4ygNsJIeayuF//dZx2xtEJgZq
wFRUf/wvMwzRhMnhzUvsR1z1qD4r6Un9no+/RF32qHiNYhcnoChgIm9QAAQFG4rq
je3c1+gz8BGefDWBFSACZ2Duz0e3FHMKBL/APhp/RIfnBsGC7U0B0J0YgjSUZce/
BP04L7SJDPf4JEj5xyxPoQa+iUa698HJRcQWNpXB/UWdM/UBChitJto0Zc2ecycg
qwnYIZhb1SizXo90pBqM4PcIxrZE9t6ylQ5EcE0xytKZIDbDfEhS8sxob/tp3ebL
drwiNO//4+pTp8nOH3qsPirmc12az0qN63+26NH4BZQe1/+aNplB1vN4e/FXONT8
za9dvv7YemEbgAqYuLtaJpU7eEBj0TLnfiCnpnwqnvK4uFq9U+yVkd1OUiOOxQAC
xT0hGQQarkrVuK8OjjxCW5WYMulRee7mP0w5FZVsO0gD69Eqhc99dBFrFW2rbIgW
NatQD8A2VLJ35QgQpvqGjtmQ554WqjXO4/asnbHd6e01zHjR9qX3JNlKeMJk5Fam
nrT1H2K1CXNIr6YavZdhfQygG9P3WstApdI8F7mMMPRnTDtvXLKNnFWAiFZawWwQ
+sBZo6Gev1QbGGHHIJ5Vn68DBtnWgE2DHdOROe67kXEJt4Gm3pLnKCHPO3TP5vKH
Hk5dodZVzORu6+714DVa1D6B293R0ZZYwCsbAW5LXGrFZEDoTICJgmKsBnDUMf9h
6lNjX5dcoOEyO4bom+Dp4ISntM5h8OfVZoiOLI5eyzd6JeYZ86Zlv7eD0H/x05Sv
pRk52tq2SCkavQ8Jle3BLUCENtE5WUyNAKl9FiUzA/yPizzP9LwlJK5smE9XB2/A
mCVn8NsSHcFA/y3g0etfgsSde5X/Jm1u+WCsWoBQmp9c96OrrDUDPeDkdaF6qP+U
v41FBxMSQKF6qxgq/vucn4wMyvERK3aSGs+QqKbZBVnrUKf+0hUoDy50O3dH1vJO
pS/iqquvy2S1dURVeUnyPpRSzHzajrbLSoBMo0DigRe7F88gDAzL/9zowgOTm41C
sPhBgIuxA1cRkzz0m2/TdqibxnrKf53WWyNO/lTPPzXNoC4fGHBPq3EWDFiClSAc
3E0TeTgMbiMu0jzd3BYIqUk+dwBPQKxg6bC6RaF2SwH879cYKtLqjoSbhUTbx3XF
nBmJJWCR5lIweEdt8pCtJn7h32Oc71wK/gkXZlUQkpThagEb+5ESsOXZEcBMw2hc
fWpCb7bBOxMGE6fxJJFB4NqlSbhnZ8U3ZBnUgwZQSh74EbI9y9mbR8u7paANEzbi
KWc4Nj8srvmsKy7bYgPaj9+BMjfkVVcPOlNRT/XxV3NldwUUj+MiN1/MgsCLR8m4
O943q/+ahdm/Vzz38FnriNeRElRgDVwwA7WOnn8r0WHuV08pgYHmrV1VPX5PG9WS
aJk996ueCm+c6SRdBe/LKhD5LDYPmgIK7Ez+9lq4ceclI66fw8Eso0srGu9UhYLL
sIbhiKUVJQ4s1VviK/WRI6drP/iGLS8dd7k9Et3FJIwVv0eUX75tgwCA7T3CSL6x
23uWSPBn0nQ7HRCb/fcDivcU+E770iTy5FBTqGfNVD88nH75qvXYt9m4U3ZA2XIO
J8Xw8iwaOIprAttkG5tCpdtfr/R3xnuWtrwsM4afIXSEZ+DkqhqwVdXdhxP+LiCA
skNV4yIGuWEh/ZsKfA6XN7O/UIuGwTOFEBupvVS/VLRN5+NUo4x/5DpICbSDF4qV
OrHeWNeRQgplFU1+uL3jw9JBT+G/0kXzRfNZXeeYJxWJLLZegtvoDTOV1+kPVUEP
YiWk3Jydzs7yKi051bn2sPqqDEbjpvAjpYscGG88gHnm8PqP3nJ4nMm2UFlIs8BS
MnnqUvgo7VTbwobc6P7r/NINGkH6esxrHOdWTHoNWJ/HhKrZG6Lo182YjorP5rMK
X+JKFo/PhaMVSdQ7BL2uGZa7DiDJvtkbFZbSqxk7ZKw5AusLUS6LS57NrATALsrN
DDNdIz2UO4JyznIcUDZohOLalCAIvK3CR/Tc7tDc4Ch3B+3qhmgSZ0GXv4dvLvSi
cxnHv/+oVj5X8xPMtft7r74dj/Et6X35sdkXESFIOtWCqhoYG913y+eXrVAPivvU
R7TV2aW21210Kw8pPdC5CkEHvYCW4EjqzSEOfVLwc7yAEex08LLwqstfiBe7Ugrj
OqYPQd6RogtyRpIH+EYa2YsTphvtO7OwfCMYyKVs0yfLHO0da15Sx96BmA5NZdtD
H5PyhX0Z/EWlJ4k0yTAx8wtqn/7/I6nB52na/59fSFoFjQqUIdgIQlXngLUSMoZg
u8O0oQgUUyJr2uifoLcOF9Mm/go/fCHPHXxfjmflKdX9t9R68hrvlaWJn79rwjmE
CWTEEzJoAY6e5M+K9QNG9w==
`protect END_PROTECTED
