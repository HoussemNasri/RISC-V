`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAdMq0bQDmBmBsLPcPZ7f90SsZX/7+dDlcQEe0JERIrK30XvFUaZOm6jTKn84a9S
48WJpUh+zZTybqhqXxgXrNcCo6yh01hMrQkxUiz6bRxPf9VDjsmGE5BpsHKalDmA
Fx9FqdC5bPDQL5W4eQef5afZt05eZzSy+bP6etTUsLU/iXI+Ml2PoCUgNJBXP0sI
kELuwMip7G3TyK/pSA0dPcm/WtxNpYcJdwZ21g5M7dHEN7H8gR/35Jm84XhhgY1L
ctcOYRnC31WUlqpHJEpyhO/G1cVJS/jW+iEp01foZpOvRQrFnd2OihjnpKjqq50v
bnhOz2rGGsAWW5raWkKLqR3OW8tPVxEpNwtgjk1V4t9fNu2+mE/jWaLgMe3pUcW1
MD58f+Wwz7iiNLtqoec0W9AyXpqO35KmVtx6mQ+YPB2s5d9OVUYk6UeitPPWPawb
DenMadrS0oQ3uizfeofOUBQP/mxxaWXGixBsk27Kh9CzVsWWWze8HKqtltnS5QjR
m8B5e6jXg4b8uZgP5QpPBfpRU+WORBYCbTt8TaOhHAhsbZzH8ehbM8CE+e3pJk2T
DxaWPsqBADyVz1/JeFoiz7uOtTkyqne38Hdge4Rg7xVvACQq2OcnBnfi+I47PZsr
3Hj+rMTIN1aVoejqGGbNuYcJYR5Y3Qf6i8ZInW52gU23wF03GbRc73uDsDI9X0cV
5VYuqxYNVCywzGdyHR596EeIL16EpzUH+d/LIi+joCb6+D5nqqCbpDUAzMsjbM4w
FDX6IXySQcboGapko1gqvqf2b8OtnuFjkxzyLt9CFX5lfjb7nRT5ldA6rU8TIeZ/
3aKB1x8/9suGTGatIgINy9L6CV8ydWXqZvt26FkLPtm37D57Fb+OCXNEkqpx8j0Y
Eq9nZZpA868H0aafHDCYi5QzYvsy2txf0/QnPM587PxKqc7yGUxpgKAyiFpCr4Mo
ui1mf1Evrk77UuPTBk4JXxSWFGAWohIe/AyaEzo2VuBsAWJZcVHtU+7AdY8R9N1T
HxcS6DrlOEY/p3jP7APQh86mksqYAlVBv/yG8SnZ6cABhyoUNRAu7XKF/BtWBKS0
BU7VxwhC3IX/Ki5QzIAZYDauHds5fOHJ2iuDaYVzP4IhXCQiaLF1IHrnxPf3sl8p
ZC60gnR7BW/0qvPC4vfX5tIqBNK/TNC7C2wLFDCdvob3NZDJcxDGi2hw81HJoDR9
ukv8uVs9yAASY5L3wNxdxh8nJYN6K1WFF33sQW9L3OhGpoxvkvTVJIaD030Jk8a7
N7YMF5EXgB+pXQVt8uWvcJZ5jzKP9KHHgbP0rtovVtRfdPQUAhS6SCCy699WOFRr
GWdyn8ZbLABTYn5m9GLsnGrnk/QhxfJM3xNbS1CBJnpLdhDpiVUHZgIfnmi3UYcH
enPwFcKpRBcofLpxP+uj23nNjaWHek/XCvf38VxYkjD5iKoK3OtDZKQvFXw7aAUf
AYDQmmrXj0sVa1TvACGvP59y7hKyQfunQz9AmIwGFmIR8Q7E+KP6h94gNLh4vk9F
zWc1/mbPXp08yCrB2dyuPGjaaZIVoelJ1RHuatwDUCzVLqtOd1fpt8F5c4qHYOlM
x8z+LaQIHY1oi+1zXXSJflL5WI8phMGqBSADlhotMllXlgpb4MsLsU/dgeUpm0e0
/85vXDA6u2jp8c8qTRI/lmPQkOgqFzsIjE9EcyUiQNHxyMr3K25DCnkDw9IUCFqN
ULnejB3/IKMkYg/GI+9vkhy9W8kgpPihZttX7D/GdfPP9hKPKaj3/Tigh+rI1ich
CU2ziEP3w1ma1zjlBdymdy9ZjbrKkg13P7XBS+V/cMVgBMQE83K/pecaVQS6jRij
ZOB8zLo98Zq/PS3xLjlK4Lf6eIcpf1qR23d2ZhZ6obmslkmS5ky7so+rxNtUd6LY
1UvtCbOJOf4QbWbtbARGr/StdQjoQaeTIZ4smeTCaJ6b286px+nUsfRjArHuwXhT
Srw1EnpgUVaAxwqaaMQCOZ1aCX5qpgrVWGANVa8OZQUXnfKKcGX+4pQqbww0Vl7R
TrvLK0AjqsirRUbPzh0FyLVE7HlJ+lvjUoN7FUdpDszeDr+4h4EyGT0IJkEY6pGe
DWZuNHu5ExuA7+Tk0e9yUO51aMUj7AAXDxc22XSEuRZZlk1HGZIyMl+eCDoHs4mA
w8LxV5KHidTzg5/7ybpdBPNDRRgDuXowSpf1Iviw9JMODC+BbUXNVzcXV9McdV/l
iqZmn+b5Z9vxno6Wynv+Zc6w9R5Vpg/2AH6zZ7GJjX2vyDc+CCGTVuLDFsdiFSiM
NUNBGAztlJTSuT70jlO5auqdymffnjgziQxgIdvGOyt7YdepWklAN1eZ8LCgTPaZ
Kd3gjgHFd77sylZ3E+AB7gisekofwJKAGKXIQE2JuimzWYaNZIIDcsCyzq0BtkvF
YO176tCGvWYoDexUNKhyU0cSXzCiV+aOCAWD/q8uDLSh4PTNq1xWIqzYeh8SYxkK
WlfH9yoeKeZF1iGbu6amqQwDLONaCympD9RDjDUMgbmW43+YasWFL5ekKr1xYjbc
gpQt+/K6YafvXL+AhGrSbUtW+evfDw7M8VroXakJZSWxg0SJ2oM/MMohSr544zTa
jd63WhzbC74zZEM2FFq0kyv4ITvUEWiwO5GwXs7UqXdCID+dJebF6bpV2WDWIssH
IJNOumJmVTLHWBNkNclNH9iM6kwSzwlKxZrr4PRD/6BxK/Cg1YWDWe9mbLL6g1XL
m9S0RLRJo4JkMy81fAcOvHkwE4/Gvv/qQJYx4BLXjqrhsjG+zlpW3mEvuwqiX3UM
M/s6ahQr6pULgZC+k+KePl0olCZ3f179hfh5+F72fEnQjhRQ3FbcqTEGzLDmv8xY
rjBqAaTSKMtNHjRAWtNop4z31y0nW0ygUdo0pPOw3tc2Lx2k7b51wX/C2tJjYGyJ
bCbEtbdlBnMfIJGCtzkGcCmdq82OWG32kyvu/pwOILGbX1aH6JIrCGxfQMRjmr06
ICT101g5OxV1kcklerja5XNEvDQb1v/Ou0OHoRgULqCLDD1KKAheK8iwwY+bPSxI
7AveyvUu80hv0ftmJfc0MGW8riDZGEHQ3K8h9tk1Vg/XhvjSfQ9AXIMmECp1JeqY
p1f5KLzKRItpB6P6XspaB8jJRW4dCKgrLAgcXUlrys1WWPLcGEIOwNxbdTLWroEK
BuvxTJmoN20IlJNpYFWYKu8QP0sARkgsN/UFginXr3WoNPvNvPeG0kuqADT526jk
6oAjW8AfatAZcF28XjacY8Zgb7ltk+TrVucgUQ1+ZOVvYSnEdWMlGBnXw405reJN
Xl0U2CnwHysmSqumO5pCOgoBnzQt9iRwhkPtFovnZLWmE9BPWiSRsmqDUH5BYm0G
uT4wkBdvN2fOuWOCQ7bK9K4kbeK4Ag2QlRCCJC1lAmViLjiX2BoZFYmA4slm1MSV
EQJKfEHG14vq8CPd9YEdxd1YF/KaIheYu3+TR9uTQ5RMP+cA19yTVE5CM4TrL1jR
KeNsNnU0OpFsxnbqed21olSBfEEbzZHbHnfp+Aa9cCcrIECoUb0iRLvRcJFmklDa
9yLmuvS/5CTUBoMkSs3C6dyAEFU2mxb3PXRYzr0Rkp867b4UUVdYhxlq5EoPGBmi
2+fcH1IvTl28QWoJ5Wr7Ac+s/+YaDhmnEBaIXHsNyzX/I+U01C40DpyDkDMpalXN
xpOBbBTZOiubimMYTGiL578peSWquDIeBFxHMPi7+2aXzsk/AKPX8KiJJ0cZL99r
SLh+xaUGGayjzSP0k+7rhN5fOXMp/5K+7xNNCszTGZ4ws3ph3AH5j+e1ZrcbsIs8
CLQk6vVjgOnjHdnOCMA6ylFTMRjjzH8H/6sg4Ozz9Zy6Nwrhph2fj1dIeQflqPjf
v/z/RIUALs49Wn42TjRTUpwdtjPdsQCise8T9NUn+K8TOYZw3TfqspfZ+kIKQPVF
Dsgbfx//zLBZE4PNlHsKawoOGUL5VOl9uwgRaUTDD/efc/14vXl/1s5HxF1tx3CY
Q3zkaXbmCy5HYmjwVrPySS3Dv3K/uQEhpL34Q52oQCAScKo1W/gLoCJIk4+GnvUC
WPmRA4OpkbdwKuPyAhNbvviAqB0hDEpsRBF7Nqxs+ecss5fSzhTLQap8TQXI83/g
1e7zEMUYrpuYRcsOYf1S4esvzoZy/B7ToHsrAJSY0bS9XPMSCzLQjFEZTuZ3WBim
zqAVbp5chBSth1eQ26njQSXDYnn66C304B3F2hxWZWaPv5ONnJVOr3GykZnB3exJ
dyUfLRcBeg7UtfMVPxlVKUPydIyB1Yy6y3Dbcql2Uoi6hbMjwLp6Y8POhLew2Bvn
sPi+rZXs2GN2XHTplLc9YblhAq7eTq7xPdHA+qndHOHUkWya6yODwKE004YAO/7M
sL/ABXYfgkVb0uZ23cuEM4f+8kfvAtrrzZUqSjHSNrIacUcUTVe9zPOnFGq3rlGb
C+gMFAcXXrxyFSOyERjBbzTVfrAEW7HvNctwGorF2zEsYkH68J4GTYZIHnTqZudp
sFsSrFr9uqVIASEjww3YT4Xr4kBBOOd+F6JiGu3oKUR6BrjsTBT+gjOoTVuI2f0l
F/Q5fP5QfR3HL3vFyIpNvej1sR00Soya0k7drzHw2Di0bjKtqovbY8EYSKYNL/22
OjoKWgBrwHkbH2nJDH2dxCJzbX6IPvBOf6olLMf83tRGbK3/nFfBx1+9+L7bmgfL
3neYIIxLaYsnRVdR3jLK2zrekMlRlQzzbBLObJGCSDzSyle+si6daKIVCVFrVAq2
elQa+N8HfxTgFeIwdQi1s8qvmyyjMzZZjcf74JwuiInl/k5uGashX72tN3pAsgWc
HHJmesiQ5JFsGyliEK9offfCX45fP6rUKsQQYxlnXPXyIqq0NDjDFqltcrhbabYY
os7Kmi8RShAi5HNUGBmBccGWZZrhoFhaAjjoscNg/aksQlXQSHexnciDlzzP9uog
ypG+WOddlUVg7YE4BNh1X42+XlkRPZbG6n0B7X5HolXV8ZFthCEX4eY3f8a67VhY
gF6VQobcFTvmsunIg9dMsjubwkbpmTe3WclU6PvR1Eni82wEuAgDpyKtiYsMBoJD
PJ05XJQGDsIrMvX2gSlzNz2q5ZSCK/GHKG+uSUXGnwqT/GpytQU/Be4R6GElsHUJ
BEcdhRMaLx3/7c0MCu8wHe6eEgeHoJogrLcNpaWrIjToOZtFx6rA/Hl8SRXSrDLT
CnPmrxuwv7ACvSyGgH403JfGEmQ1V0+OOzws2g8XgDgHChteXsMc6uvOioFaFQh3
v9kRHKhqeENoyZnjMHiIqct9dEltrfbXwTN8fs5asA1W5PQ+csmG37RMCVgsdtoJ
zNP8LVjmxGYpoSJO5FV0tgbPSV3W3EvkTHpUm9MhYo07JKKW190UyXDmv9lQ+rHt
xCBlXs1Vg/88a/TEpF7Llm7FUu0XgoaNwHitWiNbNVFZJ3A7eV4sCcqmh3sG9Dh/
KHCPjg+d6J6OnxPv1qqeMTVDgDKWkr3NzuYfqWyVG2M5DOq5WDFwHAdmgNrx03Rl
OedWiMlX1zs6hK4MILDoG783Or4F88IcpCWdxiU9wO3Sy4QjzCXi8aCdDVKYwu3y
dOT0bu5Pnz03iYbJfpHp4r+GYM9apg4MfZ7Of7GOfplf+sIgxXkxFaML1IoDCd/d
6nSFjmMDFsy/D8h0+HLC0ViulOlpWIF8bjScZQaEg0MHNQWkEj/buBihRNnqB7EB
xRszgI7guyOlSNiIKVg0bQY4UWdufsgRZxwmQCpQQculOTLH8iymb4qM4U0dpvu8
UdtcRmPdo6qWIZVO+0VSuyl6C2jooonUNfSBaEW4Os7/6w+oUm3V4CMV7etoODYV
ouBN+GBE9NVYSexp1OByB7NWju3DNAGiRSZndTr/tb1bGvQr3Zy8VNjDWoaonaJu
Zvnk40h+cdZaeiQAMLh+Zb8zXGZyX31pVXJYiiC3ut0GA0eftUtccL0ptlchjCmu
e1xVAD0SLpgOKQGc3hyoG2xNmR0/URez3LgZM3RNP5/xa6UeKQxVUwdXLd88MEy+
Mi4I99+LVX1cEREsp/W53XW+eqfhTHiNZHIEC2LfauT5GMOeIFXZKqWoos5965xw
8j3TMLsgdAvhB3ffMAAEWhDp6V/ZamcaR/tUItfk+7HTDwHnnBT+m8eYRm7SzIlC
WHgdrNZlsoY7SPWieZ1bAwUZbg/+DhO1JqQradBtNBX2aO/KdwtAnFPs6KTVxExR
xE4rDqSQ4aUbToysjnKmV9OC3gx7kaeAlm689aZxLFKMXD/8IqxBIz+FeFzrv7GV
sBu8EmtbnDwudxAo3SYxnGRzgVARD+8YTaOywy81CVsYvP2ys2L86CxDqLfDSWff
OB/sdvTj29onoPeEc/z7e+jE8y2jIj9qagJedHrRXxjHGS29C/+uP/t1PjzBVS4U
Zb2aC+qHIklIKZdufWQtgHz9j4qcGq9TazeeJhILqFMnZtGUWlazRPbQFNJ3eXpt
o31PjsPcR7hYH4Bb9JpHXO/aUs2u//yf+yjsCSejD+FkOvOoiAqQsTtOOsJnpJ7z
uYqYJPXbbsUq8bXcP5TxYOcMuLzNQBuibHP8E2UXofDBCz2rQSRM2rvIJnAiqj/A
6ZnnozjUxN5GubdiLPFdIXugB8HgVcxoPmtAILc4LCgYa+2fFx/NZmyUkUgz15IV
CH7clyH1MOet69e1yiDjukAujBZA7bHb/UA4754TKPr1qXU28ZacCZgxVkLCHHNn
JIAwJtkXDn5FXSOL2LXp06WDxouvuS1D25tW8r6+5TgF+1R1Rcq19kIOPU0UmHGg
qFIO2FJ8/1lhlaA2IXAf7UCOojHa55NxTBvwJY/KB7gaTER93mbPxxkFfgUu3b6m
jDNcb5MCUgGLVf3TfdGUdKstXD7ceAlkL8NU17teHMy+FYIXfSK9J/M6nJxDC+z+
O42EQZAgWinVULetBOQFABE73TfbMiMNkEGy1f++83kYKgm1CCIf85BBoBbo+iry
pV7p3R47ZnUS2B1GjNNhak+zcshYqSnAsv2fSmfYisR5t0+U5MjG+tiAanshrDbP
mrrFlsfy1jTOqBNEsfebFUmvyT1BdYZn7APjtmhSx05h9PRbNcVsZ6U7V7M4bSvV
P/74WQ4VgteL6AciFuRVu5yIh9NYgAvPyP189B4IPwlAkM/JftM7pFI7ZFRzRn66
T8jkzpu4vA9Nho2jTbh87RttQvS8UuLatLBfMLvnFIOAjHgxWQMngS+ybDkCVYj4
0TiY3Pjef0Y3DFcU2C2DxOVnP20iQCNJrZRxfAP7oCA6vX4Q+FE5qTHusmRap8Yf
bgxwrpn4vAFFiORAlW+bvUhApdROi6uU5d67PSU1waRYezmK0F5Tf6c3Yqf8nLU7
mU8OW0NHMSR7WBpe5w/C1zf4SmtfZrnbG3Bs5kvZ/tOsH30fVfZq6Di+KTSvjAAz
ChAXiv5SysMGab27vXOPbeJ4mwnle8oUoDeICpkaqkdn8JdXgEGzFwWDZ86xQ07m
Oi/5376bfJ2vB7oMUA8IdJdZjnr//HJZHkJ/ekg7vQZG9Dl5Kdlz1rAWFFKpx/iT
4jfpbyvJcrUuwZtwaJAnycaG+47LNiNjl4skkutCxlVTiCluSwCsd0/stNm/AItu
mpR7bEDbOfxCPQorVfemsQYAQSbLPksZoP7k3Twhmop1T0WomBONLsGWtesGOswC
YGOzWQsCET3c4Iwzf6dKWhxkeIbkLOFNXU+vT1qJj6wCKCO0R+W4m7uknEL5pm5j
5vvAcgkRISbSf+uioPv63d4FBZc9/0KUpSqI6AEtheCOS8WS2OBsoClpnGH5eliM
B5ryqKLZxRV1D2lY5/Lo3ZNjCJoCO8RxWHXPW0MGEDGitueeOpQr6vfMU+SVF7iW
daUyezG+iBVqcu2XCiqc05sJplqp86/qLMqMEFuUdtL9kKMqoH0kIUwAu4Ua9/n5
JyGZGPFla670JmRDagdZNEtSvxDOrTgsI0VjZJn3TLq3M9b/yX6NCuPHxVzZZ8ss
tjoASbNErtc/ZPBPn5qwLN5F/H5Nnw9viR7R0sTboAqT1Z10N+z6106MyLG/AffX
qBkuxSlQ06rZ2HM9ldmLpHhVubDN6W5uXQhJG9oPWALHgOuybzz3iHevv6yeno2M
j88G1dLevbUzYA6HpFxqjHzKkye1F36GqzNBJdhPqN/hHerxOp7RDHUlxoOelLKT
XYL2BI2gqsykC/X69uWRsRZeDbZasU8JifrM4R6qD7Lu+bhCZFrddBWBl/4mqX2f
zXMIlUs8GiROgbFELb6SkG0bHCme0CNXpgNnXV+w5AvOu8K3iCCAVApuhMp+Y/bL
ACKmwfK5xy+peXPVr6UOE/L3AO7UA0Wh36Abuqe9TXFvDeeKxdEqWl7ozj4Rwhz9
4H+QD/2+Y7j7AnU1gtsqjGeB0pL+XicXPL8wXVRYqXF4mTbS6EQ8iod7/fzq19ON
VbPyvDGmYBveSRmYTdvTs2gGBsrVMSL2ldZhoy96rsWqisNtf9ZkPuGTDXViK59j
rJxBYr4tJmDKGMENmeh3SnXP+8EjUTdhhupx2Wgig++N8S8NZaWTz4bh4vX9iHsl
P2QTc+FwGlvsVQJdbp03fIpT+2RtVtmjh5wvo10U1dMNIbpmeUBCJHKA7vA9Xl7r
EmdS/dq7sc1p88k7VZjzAUtJQAxg6GSZO47li2fNqNbDqr30zqLeqYs5ZAPrgQ5m
Yng+l4qaiaHeDDU2+u7y+vRtjAJ/BTfdDFpo56yOoPcJfYlAvlZCeUVrBc6br5KV
3ss++NluIxgPAB9+Wrwlv0YDW9htabt7lvLtCpGJIWga44XKdfckNKAsY4B5qxI3
YhMSzWMH/8CKKUkuTcMg0DnYkDkSJEXKUYKuDPiFC1fx8qkwDhMI3L9vWgW92+c6
nptuoRp+ziEHRkaO7CNdU5MAONCTYkC919U8J+/7PsfDvE7mLGM75+gf9blI9sNx
IoF0ePWuWQeabDN96CVAdbnRX0I6QJgAPboee+xhHS4dkU0QQzAmI78/szh8ZHmQ
LDBoNR5+R8z9w0pDXDiVnqhHtmFkPhGldffqwOrTKUlV2sp7fhZhaEOBSMoV7vmG
AxIEbE8Ytn3XiKjU0MZSvDlO25JMjHip9NBWN+nnpILi2v4+DngWaAUgPh2rdymE
TE97yA8LOF/Bvt0BDOg0I+y6CfHQHougpDCbaL5bl8k1Yfpgc8ALQc0w5oos94i/
8yTvVMQLV8MIdMC5y5UnWtneg+1N9fn9ktxWNIeGhhX+m2MOYig3bQQd7mgQ/h9L
9KW9UNqHl2clnUSvSN9005WMp+rtiX4kuYk1hzZ5W+15Z5YfMu7T6NiNb8Vw8udK
cUWPUYiUYSOhpFX15TtXtsZ+98xgJ4LL7zUU9+rFhmuPtH6oKe7lXk65Pign0HR/
HG1EbqU7wHBwGHcq4ha3mWBV/wn/1mCQWAS9wFajhXvOlGh/gIKmyXLo5s/KlDTP
SRrxBiZ9kYHAa5ZiG+Juctvr6/nUkyKriUqeg0XOjCnalWbK+6JShJg8T/9ZWhqx
EzPYB2l7FAAO5OkoDv2P/Hz2uWdcKYDRHAXx7wjNIUb0dtEhfOVyzumvb9cYkbJ4
0mPYuOxUigmdLHYTTTAMSPdd4sOiahqUAd9rRA7QNhML/SNW8pIcD09fiRU9ipi0
lhHnhJqrv6Ok659+Yo/NzYf2ivEK3mlCEDy0nhauCPV0YMb0HIzA1K58HOYF9Vcu
O3LbtmdxKQ51y/HZ2HJvdtRDLE551zIb25gaq4UKScxSS/CzpSity57NNPSnzxVG
T6V0GmrWFjzGGkQDjFCF60QGXoxv2AT51ZLkGHYvdFsffMkpo8vtBuRgsGIAlG07
LFEVQxyFrXnCixrPJZc4b5dM3aYHQS0WkZTw9wrZeoloNCL5mpN+rnPvmoKtU2Vw
TIVe8Oja1s1YrEbbzVYzemqBXFsaF2F/q72WcuXxDCXcM81XmW7wp+vpelvios0D
tEwJSTXjMzzjoq4pg1bTblbK70c+VlqWZYAUbTLRjIw4BMcrZ5jxevBmMMAvF/cj
oOt5r4PuDiYwneQd/T66XB3Ngm7FLzcB88Ug/TzAcuiAW+Dr3tnBMQEjhHCEEADx
uHALBE6NGTLb9IsCmPrqYQRrPLaKK89U/YDr0zbU9QyCUoEAadVi4UOTGBXdW6gP
Kt8UH/R0WRwnBq9l7ZRITLQh9r0tOF0bLl/EfIrwQOOaXDDiTwLGmmQg1QtQN0J2
w/ZG2dUomHBXe8QwRED2UrkiauaVxfEZF22QxkE32nxsPNOdjJ6M5px5iJdfyaSx
m2F3EjcmEs3k6ZPfIIqAZk24b2slrz+juL+xsJ7U3HTua6hmXzh9KuzvGtct6fW1
CnTbhkSY3qX39i0wc74Nia4lmVjFtONII5P8hEx/K+fz9lUvP5b73voE6V2lmPUM
u01tAOCbdTVLF+qsCyvPNvOaSgYWgxn4lp746zxe0OUeFnKhDWVwV/1es7yI6y5q
xiHAwngZG8++2MmF2zdApHIrA/dkkEIrWMUNOHAtU3rWQO42Fy6g3bseNXiKVv5s
cR0xks3Dinup3qNMGLtJeg7/8OYdKIi8wrrx2N2exVYuVCxsonIh3pSDvtJ/LYWN
O5bW/C4ggVm/MNS0zyxNzWk38S34YIajhbdkVU/iMmbbXrMof0oLN3t7nsO/vc+A
WwmDiGXc9N5e2ZvaL2dlR6Q4wTkZgEpFKxNYWqd9vQ/Q9QcF+O3nlYDUmblmnOas
Yd7jY2uIdVA1aSS1yTpm+wWL69gowYtrrwASFU/A0NmO8A+Mj3mpesuhRtZDf/XY
eG33H3pveej1g5atrmvuUNF+N6GQoDm89O/8OeTo10rq+mJ0XrVCQN8Jlv+X9pTZ
mpl7XlZgEyAD8KnHEy+5zBFq4oIHKAiJhXkV0j6YW9HlUphtpaEgOvBWuEKhIUP2
EQBjbgBIYwjBPCFcnoA+VZN6rI4K6kVXyeoTwfBU2ybfXy3M69+6Zdzht7cYJzB9
pIU1Zn3Y2CNQmUWYyw45HL5oeio3DPP/xZFJLBKEPXWIABkBPbYVzEXM8SKe9UsN
qyWicr5P83hsfufJXShpVx0tcKijGBkLHPid70zvCzoM3btef99qk971oTnBS74w
eYND4n6yN0hwkDwMu9wpgP2rOhERJ1AfcjieMrTqBne0JEefroEde994YVqhRNGg
EjQ2z6wHMa3w9zFvTtf5EmNjXi31MwUKNP2paRybtJ38qdo0xChZTuGspCZ5Pm8V
VVQ//ni98Rz/fCQjB4lFZ7BuI6UtDKrHkv/0D9brdnbOl6eI2NQgCKdyPFW+UENz
c18kvHtLIZ55aEqNR+qOU/Bj82D+dqBgorHJqu+npDKyLolWGg3V1im5jfyNuztZ
vCEWQzF2Q7YsAIKwUEnSkQuaXDmWr6nHenWeQovdwL/B9cyFoqVV7CsPcKrz4Ugi
yVM+YtUxRLaDWHy6NF9r4jf1deo9XiEBdfdtdmucgPGgI4kzYKHrXyifl+IXqSWa
48Ls+fscMQv0aNwl5ri986wacGqDNV0HbPIQ3T+/3EHEVmbBluVW7zyRzkpPwhOL
JQVO6hT7VrExxuNx0DBnKU7sIY3oVUidfv0yh+ULa52bwhzgFFm3h7QJ9MKrD7zU
sjVU7fGpMXDhr1oPQmo6XXsQaIAB+5nxbfTRJ13ZUMI56mJpkVctv7fanB7SFETD
a6sLCipXAG4sE2tQtJ84imkDEmYqky4vbDY1wlegO5RESsijFGUmZRfKP6f3/daq
uM4eqGqfyhJzGlyZIiCBLNDE/xQi6TQTiUVtgHNEKxsbqmIiUMlrt0kl6SSbQ57N
bJoBwadwwtW/bdUStuPsvS0t6UreLX6fZbe3rC/dsWV727TkkjQdoqcKXK34UQQZ
fFZtwZR6i+zShIet2Q27NZFkZmzG7sdcsPeXDUYRUZIflm1o5PeZz02eVanOJbmW
9cEnJvUXq+TYLMy+XguA2qVmb4HcbJTmESWeZpZIUu9aap0/+q2txOXr7ztRggi7
3KM5yedYxvJJL1vaKZg6Nx0uqfipTY7DsbBFbiEkVg43ph4Ntrl0Ci08snMwTQFS
AdlNFR3vS8W2ZnifpzsRcMJhBe2Tw3DQmsCxT2COhf1sqyUd8wWSnYVNJ/ANsqVn
Ucu+RKQfijTGO+AJriczP/zsEPBnRezolzx4oz7kpdO4kdVECzr46m4chvTjwuFa
X7rSK4pxayYnFhbMZdX9RrfXDOkN8Lpq0Bl5z/SeezXgHaajyyfQVhcpPKeKysbu
dmzz9JEjOGvkXXa2xoUivAW23vawn+2YhzJLpo6BZ6BJTMZ4bFrFYzU8gSXnMAV2
MGr8z1tjnB3qv44HFJePBCZ2zRMBnm5Abvnh536R99i7knBB8Jxk37N/Kq+MRGAN
/R+EMa9hYofwln8WLlG5vwBWaOLOdhFanmIBcEjcWqCm8O07YV/5Jsm8W50g1vnw
CKErvN5HYzbgKLse1mL3QoyNikcptJVzDqCKjl/K56OaiTCfCFPl8j5u8QgE1Z7T
7JEGk0W2VltzYrpiKD01Wu3HrWukvloXSulCrljoJNjXg7S4m77gv2+fMG9QFhUV
Cz8xgsCS6Fy9i1t2CH1yVNsYsk07k5/+IEfYOsJQS197WzRpqfhv4+RgRFWgeLYl
AiD2Wmk6x1rV2T8MX7N3n2zyW9Mot8AqrWean7eiB4I8MC323duTJmz5PYyMIiP2
r7bgRwU30W6lpbreBcR5MsJA0NQJYVmOqw+xAGZPENliDBf5XqEQ3Q771ZaZC0Kq
gMyZluflUlRzD80HCuPPBpawI215wHKbUcbGMIOUAwBHoavd9vb6tyFIrYBKBUZe
KFfZITIEPtJ2CBe717DZ0m3A/KJXaEj7dvOTexh6V2vr3mw0jczeF7X5hyYuLQE0
lZR7+MGt3E8kBM9d4eMgLwJTLJbYfH3//nK20ys3OoedrBwsU7o/YuygIRtdaOG7
jJwMulT8KPQ5wquyxksuUgf88YYYfHYAl+833JmTuIEy+dXvEbp73hAP/9M2GpZG
Cq9jQx6fqY+sb+xBFWas0Wu07CrQhZz2mdsF8sMkPr6/adyTiEahFqhVOFzp3pLk
+rAaZYXR0rS2OF6Sl5l5F8GObg+OJXfGJjI2aMGeyRWnlpDOxCgBk3bfP7ES7QIp
YUBgdnfStG5/9M3SaT6vJp4bo4UgHjW9RwAJAm6lj6toXuOnmibXtaMKNtt0zsU4
SpxfhAu0JfGnVXwrBDxMms4K0Kcyn3IE9t7rTgbzfDKeWAL7PCiPD9NOHJ4QsB8b
ikB84sMiC5w365UcMLrH9Ftdv1t2eKVfMFKP2zsKTJQ0MQQr8wCUrZya6N3Ye0s2
PVLkYt45hT75y5Vytmc4Aaq0JvpukDbxcfFspKyAH1UpAjyRGrYTtR5aAUx9Cn1X
iEUBOhSeP59lEpDPHZr5/7TD09lWVAq8rhg48DKaxnTCU1jIO2w+Iqxz+YKzAz8d
V+6EKjL7rOF2WnxDNVZK3bIXPGgp1dsPlHMRusDnRXNYtaq+PzcBirbM+sm8Xu2O
CWhVyGeLLyP6ZwbJFUdHnKYGYQscPp6Nx/I4TXUYN1k5LkUsB8IyYxUE7t/sjUhR
55M5myyio1G8hMOVKDWxfreGKKOK+ANGY4F6JlwsIBN8hRGy95Ny/toQSsFagsTG
EMgUSByvMRbPTJoH9TIXpC3gS2yGTKYlUYxWrgMSZUbHOF94tnTeZq5mEq6BYgUm
6quqws27rBHAjQiZY5Sy7OCPoh4P6quDazQXejlWqb4tczTUoCOjbTXuJ+tEeQgb
GMdnm7+ur50rSrMtoNmRuJ/YiM0eAqxo61rlvydEnsfRhTUeH23uwgk31znDLm9b
DjDQenyRR3FvRBuYWHKWR1foXQrvGAh3IrB7VCr35Z/nDEp5VzuCT/K6qQY32Op5
OXDq68nIQq427AS2w3Plrx2K+5Qf94RfkQoHUIDFl6UfvbA0vmmRpxqTUPqrS2TI
lg+gl70HnY+F9Y2sWAFP9RWw2lsRuz09GFVY3tSxUGd9cXB1e8jjSIA5DTmnZ7hf
/jWPROt1UKVQWvT6VujVn3CBwRl5vwe7uPTw01SvYuMrHcjU7/IC08oMFbayx7KQ
/G9qY3BDILvFCoBboFMI6zVK2FNukef1K4OrnZ+eGWKAz10ctNSAmoghsjvoASJ0
8iQVck0TG29ztUziWcct8I/vuw2TnzLFlRGGKOYdJpF9wP6ps2XaZXH8e9FfNWmu
sqPY5gb8KFN94QiAULnxoKzkOCix/JbvEUftdddtbZQH3sIYv1R7Y0rpPBWPpn/L
gu/uaKgGAykDc7Y87dAKcPDyprVZwzK44yIUd+ll0ZNmdL2aarcE2sEPfS520VT9
qm3uwwsPaLCFN9DrJaZ+l93AQacHa364fcjJtfUfwoCTL2PUF4+xD8b9LxM0OVMQ
NjbwJuTGrzf6DFdUp/0iUiIKyxffCwziznzg81mQwYKB1NZXh4XSnDRzY1q3Sz9I
27Tth0ni4IDAjqqo48Qel4r6PA1wya91cxi5LamRQCnF/29oD6H6Y0R/QetEiCoU
VQmeTMUvE9ep53cRXKyyt7OSW2WBsV8NrRpXUjghJqFd1VWtuTOkEsAY0eLDVDT7
4iWW3YtQAcEwsPSNEKTUTNPq4cFX6dsX6tUpspBgfeF/O6ueqgyX75rvliogq2cp
TgLnWECffuF+q7Zvj11UG4Ae2VIJj2cEPgOlLwNay5J6EwyjB+9UsOPwNq5y3sRN
HjvNlA2Kfxfz4NzYYQF51fUJD4MpzdHkkHKua/g1N8mJRDXQdUPT57S3JeTCIviY
taHK6HN4GQHab09vNcZOR8jWBLLZH83wgXwhPLO5k28aI9eNdy1vguL8g0SRa5sG
OBAY7sQhB1dLOrICbr/QHGRIfTWOg9F1tZGy2EYoGFo1hoQlOwUlX2edMwQ/yeSl
DCI+Il0/pLB9eNIEP2lQrsQ8FQRtAAr77hut21cUaYTX4lpO8SaMdc7XDrpRZZgU
fA8A5GWGD07tNm5Z2c4mmwPsNWkTsX2HSf0z5JGLKFrFQl3/xJSHCcUy1UJwXtqB
s+xRjc2c6++pkaAhTppejcDjEyvExZlNQfmvIe2e8my4u5aEXp4NpeCdSkhKwI/5
Wqtj4VgU4/5AwHhadohm/pOx5Y/LWEpqabowZ38oWAm5Q/S4hkrBK2tVhf8pFas6
RUvsmStXQfMcke9iLGsnL1tSPRY2+qM5mBZbp31Dn7wD5x/uxYOIziohyCSla09u
p/Ca9Y1yvVKXj6aDtozv3ThvakrKXq6S0EY1cFKT2mQE+iqsRvsan8J/Pf5Mi2Ua
MnNCX2cxQ+F67K+BvbEiDhXJnmUGo08BogIE8fDQnMN6pzzz53a9moXEotxDo1YK
rH5A6ZO7GwWQdcmo/Zh+m4t4QVTVSDEU72im4pk8S/tqACHOrzvx+Q04lJSyahDd
HQNIlW73e7WQRHkzabY0SlCGzRv96Q/KKU+1Ltzq7wr2CO0AUKW6fVWG7PBIq0x7
3Rd1dGzp++Pbnj7kMe4DjdTgpjCNcRu6ptmluL1FcRpLd78C8IyHmzS8Z5eJ15hc
bHhJx4I4W4Jb3BPeMRtPMmIqiZ4OyOxY3ml5oIg1BvJwOSVaYrUNSQZqkYCz4haI
6j30LBNtA+1slu2U6Sqi8wagKG/7TyG5/O3zPDlh10nxDhvi/TaJrAKMT/tSov7G
5RIPXBlzbjZsb+SHGOyRdTQTPAzw1jDK2enbRVBm/fPu8ERtSHP+a4rk3lycy1E7
1aGEJVNPmKa3GdmTATT3da1ktEwbqLtjYliuT4GHOigcNMcRzk9l05RlIgh92b7k
NdFJlrD2zBaf7J9aseoD1Tz3tp0Y8m/HlpNYbyE2OYEL45623H5FwL5lGlaDgQjw
yUSOvab+fOVuxlMkTrz+7OTOgfMBG06bUVK7sEZBreN1AFWVtVsaYKxpAl19NAv4
XC9HOca1DK/UclVZjdzsMTyb3dV2ocpCQHAZsdTe5X+VEP3oGN3eERfx+oduz7CJ
AwdUA0xEbtAEYNhi1aBI2XdwuN7uEsAcP+GMoZiSgjJNjufTbbD4RrOsSIS4jPro
SxuwHELXc5TJpbBuhOnArS908JA8m036rowDRKbJYZlbHcKVuin4h5JeSfCPN6Op
YFk/sHD9Opz643BgodFr8NFjtrZMUOnk/OsqkkAtwfII26pVBhOlbDTYOkMdhE5U
BtadQFr8rVfZlfcPJlfbtQxTkGArLu2pKE1gDcOubIba5BO4/JdUp7uC9/9QXuuR
xskqcmY3MPnX6D1q0qWceMJ0bQJkDC5aokZbLs0kKuJI7+6nfFbdk6Os6K0/kpeO
o26ZeDu4hnJWQtWpzfG9QIudQVO6Y7dWXKu1RtJRO39mFt9Y4i9Th/weYVELomc/
fF0lxJtoyrqDv9i2xLFOH8GkmXeWywuxB7wxe7tsK4ZRMWLdKbM1IJqnBnBM9xKf
h467Ysx+kQTGUIuJNOwE8f0L5c+j2ZtxqBwNs9R2lyMuD74AnRMixhnXvKMulhCW
Trr/EQz80KpeaZkbWHLpGg9qnSU80qBOXosCAr8sH64Oz6CaUhs3igbWGwVpMVsC
PoRDBuDC6Na7Kj4RRAIv3VZ/rohS4/cS+BqWdBroW6z3uTT3T30+YqTwR2ACUh2K
GiOrnmr7E1ab6ji0QRzR5CUvlKkItQl9Fx0SiLjwn7GVg9a4THFSomuxhofJGDR5
rgbbR1ZN+5OrRa8WA9Wg0jvJUtMrzHQ9u0lO+iFFbu6gtsW3qP2bl6c4ElFh+JBn
gmfo0xsOhIP4L85C/gTqUOPCI0KIaTfp8EkUBOT9uYzneKtc/0Ahz4JNyEqUz1YY
YD3NrD9YyBEPB6ZspyRLp9WmFtnqrN0tuEwdam0zxq0AEP7wICuwa9300jMtAdUM
W44HuuMsuJb5Zo5mDO/NTn9DLOriN2wyBhosDeTxO3+qv4aR9LYVJBj1IFY9GjFH
g9ebHAVnXvGxeUrlucaoW52KN74zIKZ6yTAmRMlye/ZH4pmfnuuKukxxw+8V4gED
9YCAsIWsPoRZkTByCf49j1EdzmJYgZUkNNP4jH8rP6/RRvdJ3LK0CBwMnS5CXzBl
PHvJ3AhOs9HHJkvMe5rM6aUdzDhJilxBxgOsFpr2/rQbmFYMOO43cu1dfE7tmWr5
4Ew2bGtu3zLUoZxevXqqDuerjQhAEkCQto8Oixp/wSsi19jKuwAu7+cEk8wYCe+q
92vxNOvalDrLmbKNfSnt9oNbdlCACTQzWzCH7s2ls10Vf+nukRJGtcBvhTaHsSu4
FsyO7uzs6ZtEA78H0ivepYTRw4zByiY8BruN9ki/RpL5DvRj9hxVRw+9gW0umM1y
Bv2wNhIVOXlAUVlZtzz5uDT9Z7o+nPmuTE9AcYmV3LQpfM0f8+8dhRBqO4BrK1Sy
wn/7Kmechh4hJQwGgSsnXzm1zx+eC3+lV3vs+rFJGTzKd1fyUKTBLuu0VOLKWowY
bllQTYJZRSO/eBRWgbjRU5R2Faj6YIWguvsIIkJgJTODSJPmz4iRxK3z6H4Ya7Vs
SWQ2OqsJwQxX2zi0QwR3eBr6cS72Du3xuAAPzv76D5xXsq+/GluCQVp99vmuu5Hl
EOzZ5hGQGrotNklUT+giXS2FAVHXpNQ8wobS5so6OYUqz8evivVN9jdusbV1x5GB
yMTICdVNexEWEzTkCFtQDTL8wgJFhENGWN3U0JM+CZ6IJdUxWpcdB0OgDoyFuRpJ
NR4Z//es+ppQxnymscmUj2NltnHPaZGCa3YetAJTvP+3O73ucJUytDXQn4v2CoWo
eQubLsv8trmEP5rf+e/YKxSrNMiILt76nUDBlctWymGF/i3TQu6BpDHj7Ti4X/rF
H6w3MWSQJQ+lrb66Yc4mKQoD7Gzz0Z//dHC95LNJLTVkfQt5OnvRqJhltjpC74eU
IAq9GLsBNvlx5MQfBgcdqjHFjTfcGLfNL1o8zCOYa6BoVk4d+cO4J5gwWJfMMN06
amdCQegAHImZJ9ahmfLw8dl1UGKvlk5mV4NO7lItDl8GCxeyB1rMqsHxiOUCffw/
epcp4TxajszjkoCrbpKN8L2aaBwIqzQPo9/XkSNuYaXcoHZrcYE/JOSPF9hi5yhJ
M9xPFesLHFjxL+/qeNy9fwPLA6kxAcr1s/cKfZkflqpCUZP14SJ1eLkimAE3YnN8
TJFuH3cpLhrljEYmlY2SmZZ8VJpkKSxOQJPwQblY67yS4VR6F0opWcUkfEJP3Z0T
MieK1WGwUMgInxx4yNz/XffcRIuJuI61x3PGhUB5trBtqapGrj6gWegmWopQWyEy
7pGC8IAnQi0Cqg0sL7sXq+mAC387H/gwq5fTGOna+UHr92MsLd5Vw+DZvWHR7U4P
sCKDtt0eQXTqc59PFY8EPNDqCY4VSDipkeeFy1RvnIwt7ph15BAbXnkYKByhEMob
ty6hbK5jtJAJkjFmwBCQ9dFc/aSu6UqICjGr40NE7Bwb9bMhUHw60P7xmdxFmo++
N4qIawOAR4h6Pjv2DhkfpTjDCXyPUrfXMsZj1Z2ScuCGPq6zXxWq63E3QrWgHnNf
5Zosg891idMVru7tpAwxFhfVYeuHXGzET1Dht8GcCR2MVJQnlaMXAmD6gP8IE8gm
q0ZMqkdaSo0DEag9zz+jt4S0kvSnumsDmRUYQfHotGvWLk4519Crcjc28qPU0TpV
0+CEoq7ZoO0KKRm4pBZysuxoYFBDc3IZdXKnnd+MhTh5HsYCQMqcd+WLl4lvw47e
zJe8PwzAi8ZzRFU6XqL4L3LRJ9JdTrYlD5NyKwgMPkPKUhmigEmvaOEq2zPTzSSD
QsmO5KGyLKI20KbTolEPQazAzmxvwgoDdoDw3gvS6f/rejvGMDrXbeoH7H2DuUcU
9YZPl1yz5KMMaazLAuPjFXfqoRS4qdvLqfYpk9x7gVo9dr/xJnyehxma7441irF+
Y7OFGOIle/wag9rk9TaGNyB62YFR8Af5hf+NF4w64r5oUpZtNI39KbLGJyNiycCX
0+eDy7oGuFUzjzqCgoAIoC5+xxkN1VwZ+RaQyIVGmn6rE8iM1tQzZYN3x+1DAj5X
5d4F8vbKYeZDmkyE/4HsxDzAbFuZhFJGcy41iVirPJ8kpur9/BabTwNPDlYGQ0NN
CCZWEDbgUjGPct/rp27BJpAjQzWHceEv2H3qqiN42x0s8nJAAkmsDoJwc0Ut2lTB
Y02PT5KHm1HGmgeJbl7nYvvt8EsZcxAYQ5fr0Ew/RlZJ+HA+mLUbwiuo6rX2NMfn
atSnhMGk264EOyT2sk7aRidAylg9vvMhu30awvetmw/iUiu3QR1v5zImDt88UkXN
Uu6pSNrv9eIawGlcbcpQdlUnOR6nvsS1Q93/HJ849p72pEPMbGmUG8jsTVooy8Gn
ZAq2g7PBu1vI3A+jFMccEG/s13SGCCnRAmITzLOCrh2VyG/vvI1XUUeFC3sUciBn
lVUyAtbC8/pvhX6WpoQZ3mp0a3A/cf9eBmoECosBIRaapfw4Z40wt62LMtSifGFv
X2Msx8iW9R1TiBiWuxycTG1zOXG/Jkasf6nRiqxU++si2YoxGRdzvUDgcgo6tE2Y
N4WqvQrdW9JbrZGKo6hGJWiIp6z1F1mNSPpsk56ba3S1wEkZdokHDAFYdPcCPu5c
xO+fudp61RowZJvo+bHRfIJ4G77EaRdzwDepBu//iHBtxZtPNRE7pZU9gGRBwxO4
jvykUiBDtNRa1uiXG5iN3i6r6zbS6d0cflRg8xUrwRa+khGgEa24+7cIW0bHUp/s
T2DnH+hmwEMT/Fosob7mA7MMiCw7hxxnzNNPeIh71oaMagz8SmNHg52ajEr3EJCP
GXQkzf+ac71UI9WZB3KTlpsWkn48sORxbyP4dU7kf2pQfZ7G0Jd4DJwuB11k2MzF
2F1qsishZbgLF7c0+vr+Dvw/xNu0sQocQQVPNJ+xHYX/HfV/3iNhDGUuLodhEVZS
XCB/Lm2LNxNgXdLbRnLlu8c0sDWMLOGbUcgjVLjP9LGroGERDYh768D4GLtbX/2R
WyQ8ncmI4Qh5s72cOpS75Jv8HlVe7y97MwDYSplwHXbJfKIGbApZc7qVGoAUTpmo
u/dV2oezkXrmmnOGEWq0/JrAKojZU8oKKEyXouzOQSb9GCuKw/eWxOvgoo8QkNMw
qCDjLGrvW1bplft6EoQYXQuh2gVy/hKfhDF9A8N3tV791zEMA/M3bnVGGfEFqP3g
2koWm8lnrQ0XcubQHiTW6XkztJg1ha4G4bDbyck4MM5boN7rFEGo7VYjXRFHsFo2
MAS17etOKGjq0rWG2Ju7bJbBFiNJbaugMSM96N3knX08ze6fNJfwltsUw2k+mYs4
mZFgkqVvd1z88SrW7DHLldBEWAMrGH+ypnW5ZecNPDOC2YJADTuh5e42xpfsDGQB
IdBJ6W78MIvQ19YIF0MSN1gBlJzQ4RWaqzQ9cgqDuG6N7BMv2cWBM/rfSNWHry0x
iZ0upCyZcYM62QlZO1660Rz6oltl3L3md0edExJp3YmoPgxQn4hN7ur42tfpQwIW
cSTd7Gl2GMsoFm4HHzO9vKJbAANlnOg44sqa0evMswfX84jUs5bsS1esY/5BMGmW
hSZm8nh5dlXyJk+uh2pzSq2ML0gFBISvq1TP42blzYr2z0EDvQVIjCyppbJa27HO
J+rQUa+Zb4c7TvhENKXwassakxRi12bM8k4vVjHvOCe8KyBNwQ9bh4QlD8m5NKqQ
lhefCVv91HqT5b2eOR/0EfU8oIF5F4jrqXyXM47561dlA30LTYfWmokPnaNyA3kY
XJ4zjy1gylhE36EfBGYwtV+byRQBuURa/93XxXiM4lianIkp2Nz7aqosiRw5NFrs
HE+B0npoakVA62X4wdu2REl7Q/R0g3SFbbYw8WuH2P8XvDnDQ1XI/FiM35TFOwJ3
VK80/NY2L7PEcZX2NQdcd90yNvlype72QY3g7P6Fh2/y5j4MoMbQmELbrMsF5IbF
ttFd86kdcCvlI8HvuZn+3imNK3Myh0A291fXgzJhhwLT7T3UXvVHbSIYHbWylnZn
gGPTSwnnwUGRlsG33Rp0nBhweqQFqDNJiRPreHUSEraC3sp6mcRvSsSqMU5pnjyD
omnHgu9wcyM+FgTHH6zzk4DEWe9WLMUUDiw2C9UvJa3f/I68AYfDNIhKLLfBVI2t
HsSNJJNL897tSCg0z6jwt0ByBd+gc0Hn098Kdfl6cNhxxdGRCnW/9OoRRuO/OzQY
rANJsWDr7JacHAR5kQLS7YM0OoqIa1o40NDYuseuGgy8UbfcCwkcUF4NrYOVs8U2
mLl7lb8jew0BrFoioJpIJt3CQu2+TlF7W4ZyeHC1IJrkCOGkr1q5QnwmCmNmnkgs
otMS/EevziD7cuWf9COTHGOzOuH1BTn2EGrkvHPYcNbpHEyNG5DmL7qzsMRZyuqz
F1mWDqG1/TcChgMP7PpFSrgPjMB35wjVdsChy1/KfmvhQ8mdpqdeStwB2p0M20+Q
52CpAZBKJIS6kt3CLi5Rlf+RvQi0by+odV+I6B1GyRXY+y/5yZBF2b4zdkIaMD8R
yafrXp4+0/uTVgKo8wIT6uoiAk2K7fupk8i4D14EMUidELExyh691gisZ15JW9ft
UpayLAGRqdvizvHP7Hi2AuYdYyLEo+sQu9/Rxsc1n32ftXM7nvqSVQjUV7ZZzylg
l18lovQyT/78oaAAm7y10TEEs9wZv6uhxvOKbgDLmob8pZMZqSbJf0grxoKpz/hf
J19Yexv27ynrtzHtc1CHP2IuWqFJrfSGSU8UkTQRFoFNWM22lzQcrGT+WmTJFHCj
waaDbG5p0Vc58sf80wthf2cMxK1CzD8cQ9ode9xgaG6KJiNzRbBIT7YPpgwohMz+
JyiJARuOucS+EeMIjfdjuEahOSWyzAc7Ggvb873coJlND7yTlpQdeGuyukI24DeD
AW0G9XwepNs80w1Kax97nPYSNf1HvYmEA6QWuFYvTnt91ZBwgG4kv6yw5ICimque
51hAwe2rR+E+CQEIXjK3RkafAb5ZwtBacRJuRJLt0o22GlPhToT6e/3qRTJwdltH
9a2WLdUn/ByNEe2xQlY5z9+Qn7W+Xs1GqIE0PSiU1UFTH1hD7wwxlr1oSlUCyEvP
PpanulJxcKytvTj0MSDhB1cE+DyoPFrOk2wba0Da57jJtrR4ieqOzXFGVHoF9xdm
gsDtsP/GfaCZMMm6xocsUgYca42mUhb6cNQAUl5RnuvhD/arU48VezuxmtfMZurl
BIgROw15gZriyo5AoFYcQnbSkATWh1f/pQeTJJuYRm2I9WJr7AvBOwMTKCeXqJwR
i/RFzju5VNNdRCXlP5b4hTigGQuibB4g8A91V3RWzt6VHO5Bi5w5D1k3KIbQHPHB
FWZKlNgicohoIRJl5w7NKqLxsXZ4uFcTTmSYUk8Z38XxjNv/Dt7+QiO/RBLcNCYe
yb/vrsVIbTAm/MzGHtVEtUtXghaRKOgF9TuzHWy/SgUWriZ13H4paXrO5HQw0Jrf
ajegfIgN4rViIBksU02K4ii6lRH34GT4bqphOZzZw8Ou/myMGaRXnY0lrMBme1IG
DuLn6FnZGQE3hsG428b7ecZ9uZkOtb8ZaPcmrhPOjCUD00WM0gBcyjOmYIJoGhES
SlEIFBn8mefWu5vf/baplN6nbG6m1aTv+h2U+qAIYdlNMw70c7LJoHEeI/9TA+4b
zeBAns6hbACxCsINxiTyGWIIjU1o87waosMf58w1hIWhBlgd62zUr6jlORY1yBN3
vjBaRhSPvGTXcjPvBUF1PaAU3z064KR0joGe14o6CRtx/JEkyTignez3CylNqNpu
IywI1apbHCWESPK6ctWnZT/Lj5lpNQRJGf1svEZ+dhN2nLAMFiNvUMe37avihQ5Z
tOEKbp1x2j3Kn0U52Ny/hRRgWguVc58ue3rd2A/FyyzweA0dfsRK4wW34Dklm9iD
ttCdmWm6feVYU1I1ANoJs0ohzdCNgV9vKfU8Bn3af5uPIM+KKSMuiL1YWAM65z9t
fLqf4UypJivhKz8sWe2sGLbyl6G4/xu7E/o8uyaPr0cx8Fp0Jg4uoB7mUF3gtvPU
Py6RlLVd8mPbOeZquN9yqwFPqjJArgEKWh3nYUdfzVPeOSCTwlFrw9Jbpd9o/1aZ
DYSrP4gp29cVUl8+OFTrVk3rSBgyx9IlncRRKngddy7CqxfUeq6dG1X9xIveYJP+
ozwSxuL6LrKA8Z7LfWhMPIowKSoTG5VppAUUPGxmEpARoIpWfmDSXHpkBPRxz3Xz
ndMjF2oJJOMxogEy48KffxiWjOx4wIxvsIiVk0f/1KybCBCly77+Ms3Kv5iXhBWD
81zXCBjbCa7G4IOEX1wDh3pTwsU5JjCNx5pl9FeavYTqHxcoEsuPx+Hg4Wk8WRmc
ijsDvgniv6O9BARHSmCUv4ku3+1huI/8r+htRuj6sASX+cjDkIh3PBcu4WzjbVr9
ScNCZsTdu5a17DC9FXjYe2NMI+3aleiCtmlbZZxQqlFIppu/p4/a6kN0xCv93smC
uiqGd05lkKzlLcOLJTO3Wm06WgXaICJNj7Dqc48oMslkb3Cn9gHWpwnpIOX3r5en
pKzJsHg8s25bl/o+VT6W2w5LGxM9CMhveV8dVvzCqf58EC2uV3tRksO1Y+5SbqoH
Ugj4GoNhutxhyKwerWPkS1UHYqfVAFQefOpD1vQYT8uj+MiRUygbSZRIGVJ9QHPp
lQv5y0ODS0oPR574A36JBqp/x6TKFimfUGAnER8bpLymyuoJe4MTpc3YYEueBgsQ
oTgc4kWdU9o6WOj3b1YsOpk++n9rIcwpKGbyUu1fXyUBVdGU26UtmZFahZoH38m6
IBBMA+luOfRU0mvWJoZVstZG8B07iiAQ5EQvmZXq6/wIJh/Z7A1s79294mLIBlOi
1n/9CsfNRVjg9tfFzv2bPulU1VgsdkRGsIZRD8/ksxUF608Lx2U+OC11GlqPngNY
Og6gf8gOAdUpoTsP2BzcXm71hw48rZG+uGtfSC6bNl0QrHccfRJ4unBjTGVvxYcP
r+FSnbVMpiIu3EMsLGTTbkWEYjMwFc2jUkqBDgpyAAnWarIJIBa3w0vamYXp9e4I
y/4V2PAHAfqhBSWMpYHaM0RmlzyCQhUG9QC9v16Rlu/S83FI0+Em3pUBFrGAMK12
MxVBrdzl6ajWj0a81pLox0NAXzjQ/4CCFBLNEMf6yP9p27DStbEvFsI0nmdF+0hG
B79NbiRhCpVuasUFByq4XCfA0d/YEXzBPCzrivWo1mcEWzQQYfww2eR0RQNjlXMF
23xxWUxyyQRvg8nMk/lzuZQB8DsNE/BQAILfnJjqD9S9h2ufAG5yK9Pr5uupzYEa
WSdcJ9HoQl1FMwx9Fbp39yIEhkQ38yvVzAmmyS1WN1M/vf8kWLIUKNawA3eUwCqb
rbuy8bLNPsnm9pipw83NbXod3HofofqESSKFvntm6XoyDHXznT/k+i7nD9e+qqbQ
75wm2u252qVM0riiRjyv/Ae0C5Ca65nxHwjixVAkmvdnarCrgsqChG3kjEUPNNee
N1XFhKX2F4P+dLjuD/Sb0HGtuBrt+hOrKOmi/DVMqPAoqsNjscs1N9dcSIlqZT8y
RiQmV68ObDXyo6IxchkKsSEfzBPiygc8Rbl1DDHUjCapomEsZbDdDu1ov6wV2kF9
Xz0IPeo1Z+V2M37Nq7XXbHwprcMPG9/YvL7w7sKSQpJ5lO3N9zTok1eQrE+5Ep48
EDV1T5KE5noMUdVZw0FZBr3cUQV5uvf8H8yK+PPjBMuFRv3NWfPfkFrDzJXqytwt
Ln6TsPBdb0aexaryGxe//24zVep3WslBGdwaaPo4783yxwno5/THb1pBOAa7LOAl
6MwBU/u7lXsJ8vg1wSBGff9xiDUUv1nMAmUjCNSYmN2xQV7N6qKeqBSmONWZOVk3
IjdTCymaHlTfnujqQc0m+XXAelf7z57p0RHKwhircFsAgY81G1L2dQYLLNRMtz85
T+rsn1eiJ2sbMDkZY7T7B3UrxgkRk3soGNPnI0bmHip1hczMvpEjZ4NPP6MAAmC3
8YHNLawClC7MBq0bxQm4iQ7PaQ7tItbQ0FGMCwGCg14kQFqgNeboXyC8t5IWQDrq
h4shwJ6LctOHCMB91AIq3/SjYY3PJGsgEQQFvVmps+IEFR6q6l5iliUYzgGd3VQA
/u3IjWkwB8m4C/H570jKtB9cp1gR7SfR/xxR+uCveyWRcenX92oD2Jo+i1Z8rraD
QCAWVEwJ1AU536KveE/VXv3go7D5UcUzuMvZUSYCw4Ff6veJ4r/7YtVRdh8Oj84C
4LayOqfn+nyCyc6jGKGuDNCD3cuYTMlvPO4lmo/0nRVG0P9bWqMMrJnYULFFBVAc
kE8svQiwtfaXIq4rTYSxHxyJ1Xta7drgCPkYHNI0Kdzz9UJ3b9KtqSvFwJj1/Xeo
TPs9uxb2kV79ePMbCLPLqjDOWPC1EU/WS/O11UPpiZix68rWdx/Sfsc2cK1rdiDY
H4FG7NzXfgpkR71rZLHFr0DSR95d6jcSQjZPKnFMbbKsBATQWcZNuWEpP0LzFyrX
/NVVEWiKrCeFsjJotdjC3asFpfKwCC75BjraTW6VtUJCg6GqL+ORwL83R48/S8ph
hreD2BylRHQgjCVl7AhO0qzJmf89c+NyI8X87hUALD47MxEJwUur30KWxTD7De6B
suR8vn9ozJKov0qklOyD8TCYCKfqpdhU5Hi8+VFJAyTzR5QxAfj69k01e6W9EBpg
SBMRKsxZJ5XeZ75dwhAcMutImBddLX86Gmrr6i7H0FJQqGKxw2gSSS5Ks53YnKIX
I/ofb2DFN+qbWsONIOZL96stdePU3ELBtd7lB4quCfXZmDPsHl0ric/iuCB9Gac4
uMENXOBpccdOp0oXdjxaqftUCaHv4tMoylfual+EpKVDlg0ihrsqbQRK4zEVJPCy
Dmctp0nL421rmbkcY2G4oRSsTUq64zIN27jpmT1MDkIYhMkbiGreQZPP9hr9E8nn
XL6VruCr7Vx9FXmYDdWNtOnTdqcjCVIH5jXe8Ec1R56XIZuM1E4TYC2U4Q8Uf3z0
Qur1SrcM56pyxask108/vTZh9FnQxHknYsopKn5Qdi9l2xR5h9OJrik1w2uxFpM1
9had3CdnmH04hwj70Nyoydv4nyR8N8gvgRwtg+IqBNPKnN0bY2Uy5tdyS4q/RGvj
ta54ZVFMaJtf6T6gy49o1OhM4Sm9hvkDj6V+hRH1R4WFdtGI8XEmtzEgUyUe0XuL
ydig7+CfYUKA6gpcAtLhcW51iNzzEHY8AEe/7an0Ol9JPKiSraAP0JYTa0hA7eI5
WOWNrb71HFjhkS/XQpRtqq/4+33r4Xbru0CLmewVvD3uFkZiQW9rGP6Uyoz1zTcl
qj2/bB+yjL2CYokG0xElLqau0J+0vJ+uPtauZQrxxSnPQlclehx4I3psIhcOLs48
AKqyitUKBJfqceRJXfn8cE9Obkvd3z7mo+tiG+tv9fs1YUo7cqaV0iVDJ+pMJJNY
mdwBSBqrfJgamT1dCAAl6sRmYLUB6F3wvrxp7qFYfYGVoWuoOawkcQQhhEqLPHjs
Gb3B6yKc0yH4ioVnWO/dzZkTOiXRDb4nxdH5cvEybEd1yXdvwajaiLhiLRNkvsr0
e+Asne30+73rHmLKNzZBSEv5HJm59QMeER+/BLbQWOsJkqd6Sh6WSuOR/cAZluQ0
SjYGOLD1bkdIb1BpOPFLJY6oLkmhLoBDa8xQcE0rSSYRx+vsM6wkNuCqG+EoBkgf
reEx47zHMaw1Gj1uHdBbARaZsDcWVEkz5PYdiuVkpv2sVMG/a+dg+NBGXYlKsRKX
86EitReTrzg2ofzNKbiBJtsWZSo2GYbl2hD7pxrUOFwi7NoYO7w51xlk1TKRkb+f
7rTStCVlXYUlQMX0aE5gQWg7AmIhbsKiBk+4WIzLweMyP8yzO3qBdhQcjY8Y8Rmr
F/uSF0vH11frdex0aJrak6k4JEs1FjZd3EQL9Ipk2TfuVT9n0Xxewmb2gNQM5VrZ
WQ7Erxu55S27ZovOCRn/Xc0YSlT8nfOjksXb29LNxbn5bEFE5+282GXXKtv+kI0a
PRDictw5/RjZcelW7YGnGMtDhJCW4XSAnFERsWlbRu0LZ9/erWAfYH2jhhA3VUlG
v5t3yHJW69O5T/TsQwBzOt13XF69q/kaeWI0CfK/RHGYgtdHeMBhU2QaI7r6IrxY
v7qjb8yvIvNODnQRZy74SGmpZT2eu/yhXiWgsaAHcUMkcBklLh6wKgseY67+WBpV
PKkzVJ5QF24o7VhOwTmkvC0PC778ieaz/m0ATJHa5K7JvwJFBEmWEG/J6W3aqmyU
ydDjpjnbZzn6HxI7alY2z9BUzyvSpbmb+ZotLQCIA1h5sCPLVbDxO5LsRtHI4Wq8
UbAuHnWDPU5ikwwveJc2H6uqNHpx7jvzoSsLMF/l2KeAxTFPpo3dajhDjsbud8dA
JVXimqs1eH086NM/htZQAKuzh01I0Ou+ya5TwdS4y20TMc5VqUF4V3Kf5UwBMcPB
IsMz2E6JiG0/0JjVI7COgc/7c1qs8XBHU/Lr2olSZYeKYVEVSVEGBenhAIQEywLd
trBL59clJyR2ZiOJ1XQAtNm94BZBXOYEf3U4JQNs9lMvJY20xiwyyLx70f38eeJr
fgRLeyCYSMlrQHuFtGiCzBzvmmN3ZFkdfS3IU4pv9KiOWDxbjAd7oHngFX4wDqmE
sZ07k5RWROBnjrMMeIJ/SWZBRXZT3JPtBXNy7I4W55orzr7FE3oRjx+rHrFqPUwg
Nqi4Euc4qRfKc7CLT1SfJiFQGq66QcoY9NiUBGUjiwu5hSJYqkrgxNAgSay/dp1r
tSMsP22AQSlDhIjgaaaehNB2enaglvnyzvK7NMrmPUCWtK6d3vwccdpOa0r6X3p/
YKMTIMblXAbAHXK1q6Ec3skEc35OT+8LnKBsOP2rfsGZT89J7XFMkTCvF+bXWBmW
4cHHFGClk/ZgRtZQ5lwYG1jvNRlMkCvjNf3zchczrcgAbwJWqk0cYTNKBKwLZ2Kh
64QX824MGEOSn1GbVmJyXvTmfilBIqC/GGxVddpjtlzE9J1GowNCDsmfdQWO1SJh
+t9w31hQ0lsMNd5t31st2DVZIckq8hXvssmr3RZ/usYXNhJUkDZ3arduGXLVWehW
1oLp0VjOdGO9bnc3s0rJFeaNAtvLJR8M5hQ2fIusECxilV6f1XC6902vjrI1GokA
kzc3SWWJt/75vhSGf6Ls0ZlwIVHByORr3Q7RKLTqO3bIU0SrFaZDLIK5wRTK4e0h
u0Ax9JVRtpKtmzvP+ONBMLgylJt8uOGuPWQ4PdDE0+z7iTo0LanAuRCo/QTbiYUo
CrIMgJ9n1BqzrYGsCkui+VURSdtBm3sOv5QVWRjwzDb5xSRnPlhVfmiZnXSbX4az
4g8BE9S57DpRTwFOU50HWL85WW9SMBjwNah+LzpAAT9gOfMxZkCN3QbkN/McANfT
h0LTydlW+0Dd/4IdB4QPfUKs5PkbvJibtpnGdY1FbtDpJQPURzw96QAmG7Szbry2
fg9ddNxgZIgEN54EK1bYoFgN7PiulC4itTjMtgv1cTtEwVuHwXUrYGdXr0mi1/f2
yyGHBIrFMOdRcRT/DOeBcKLI/YArIMuX/d2AgYz2KgUHTTcXt3Dmsea3tS442Q7V
i6Wcm7hnvUir1hFIxjVGXqc5DK8KLM4WGJRRtIwa99doB10kfNGdsN5Jj1Zm3fDi
qGeFIG7iAFH4W0g/VI47fqMpVQhvQZt3DDz/9CWuE34/41KcABT5xyqlf/+CnZZt
5A2CS4HXpuof9qdaUa/A4dOCE8VGIT2pRBDaIMujjla9OZZq2UIERbYHvjiuGbNj
lppFp8H1NgPukzdm8MQ1/sGaTSvzEMWaEwHxPL1lF3nOoikoKdni/YvrYJoTkgDG
OQCGJE+7Eqv6olOE07OD7zVe8k9RL1C3BeTrVydfm77BL3HoeMoIP/GVrzRXwKem
L0Z887q/Wu6TOr6AYWwiI5XpGCNO9d1eW6CMREBfelWtH3oyq1Mo37y8+st6Lo7A
dxpEF/ynsKwPk4/z2SHQhyYpokT+Owul6XAlapTClbESVYZaHeMOmQs1FAmArV1A
CZcf7oqK1UIGQo+sUZOryIiynMFCItz6Tf9DNnyiiyb64ouzqA+tLfudqCl3URyR
Cul5NFQZlrgYRsx6vdhHcjQ/tHiGg9n5Em+k4Ps6vnLQFvd/E72ywIsq6NM3/Kz+
uzaJyhALwsSr/dSyk3hNAe5JXbi/ZtMyp9ECld0hE4p+vCVdbQhlReqxpoqIBJmJ
T4lngk3ms4JGFBKWGfIbY2qUqr63h69IvUaQrG13KAR8c3C2MoneVfKfn44hXC+f
DGOgKmpk5k6T39+nHYVx6Tddm4WXxPG9DHIlzlqBErsfMQ9x5ZG/Dj0X7WknsTZN
oh2vI24KZsXP6ucKhVCFt5SePBTNaFnZWNCdFSwjv6I+v7Ki/wrvudSBOu7+igNY
MpihSz7WpR6eGgovZj60PTTDr4tIW3olVw8ZsufaA07yHpWTflA03Y/Pp1uhH3Kp
+lkfQE2dBrlNoMq0sI+cwINY+w8rDrOIkZD3+XtUv1ZczxqUb7FDOVF5WCUcKq5q
0eSAeXPGt/CICPXOrdN1vXqwCHz2lHwk5FQ1EdOEU1zBqYu0gXj/CIhNDw4CLSCU
F89aKq66xIhCAHiHWWc1zIRkHI97Xkvm0vSpng2mEX+4Jcxwv6xA0apH6ETvii0a
JDqfqA/T2sbcbkeoIKE4x4MSRZXtadtGHrDEcEj4REUjuXU87kpSeh+NFOZ2xtUX
QOr9zKCL16WYtDERwUy74wHIEcS6PQS6Necxi1MIdvVqSNDOorNIhrR8ZWQ61HBK
a4GGEvbb9kvpDK1/x2UNMWpxph4XDhK6sdZba9vMtj+JuOwdNEFfjHvkvdIi6QGG
r4MGzBUy7bL60SQacbM+HsfmlflR8IX2W3VDeEIL4AT4AuFcrYk/c9saJWcVdgVX
sQiu7/pGVtaBXsJHJF0zw52hkAnwFP0gMqmAUq3p0+E3hVru/fLIXnK3mP4CvwQP
TS2u9dVSPyZuuX0WYbx1rnCYtS+jV1Aurl58nKwR/+Fe6vb3Dmwq79EWibqbae9G
Qm67V5IOvd+D4zF56ldVRXPsLWALqb8mOTBImDR0vcfTlovDRzBa74BT7/DCTR50
YZ3oQMyWnetEICk3w4TECf8FhnjlbP1viJ55gvCI5jBB3caOEoo90iHSnLO8fvJl
lBWbYaXhM/VwxkDftBcXI10h0V94UadvPi9EKvgb7wYcgdCzLHOPYApvC+Xz9+ad
yMtpnkChR+ZKZjb9R3orEwECkqqb7vJI4RzUVX0MRUakJk507ASe8U6X1ZnEumGk
+n0KC7y1D9imurebgaL68ufmWSvgzfzkb7jT2R3u6DIbi6jlKN7A/BHpKW5+pCa5
mqlcZ0Ibc+cj1H3HskS4pXr2s1tjVF/dNP+1h2/bahefFZrdVaRTRQc+fPV+i9D4
M/FETahyYLf7sRPaDvdUqUB8E/RUDYHtOuVsGqEuo50cuap3bdbDckW0SUR7w4fm
PzTBahyA2xLnLq8wpXvaL49YS3LsDa4Y4AWmEshEmrILlnD1upMCqa0Nd8k3/U+D
8zwHu6I8p2TnQFotwBsYx3ZS6HqPitNZC/Z7w6FQPEEabtKLHFTYPnx9EqhcvcR+
JE8iot6LEqPiexv9jlhGW3NxvoMwgAaZPRTNrNVpC+CSaAKIItQTD8A7Hp/+h7td
gvlb/f7DhO3jgZFG20XRGFMSFRoQBUtrl1E7eQ6I0P/Zm77oI1+E/+S6KGZd5ZZv
nUjMMI/qQzuJf+5vEtlYS45jkMRfxecpfbCmks6WfawLI4MDrySIRQGkhzntuQu1
atceq0t6VczwEZ8KljWvq4LQrKC4WDUPZ+Ax4gL2U8xnpHS0MGhdOlGDNfHGDZy2
2ZNCCEYgs37iXB+e4w2j+9z4AfjoqqjPYW1EX8750xStTeVKiSwAwDLkpb4arKpA
9G5l+tYaAn8WPIRBdx73jpdOVat/fmgFiY9e2v+GLqdDtRP7zuHYwlll1bClPVba
GxrQjVEhpQypR7QEIYa5MbLR1c73W6EUjGh7sW2XRqYX5hWWrsPv3QNbBylIupOz
n6he6+x9b4pZV4kjVnFJUaxSv0jMeMYm3rIqzzMQ+UXFFyfBjfNNMdYqFlC3DZPg
Js3orxgc4N07khqfYo4tL3moE9vDfoGfIZbVuZLx6Xubkh/iqLU9+F9the8rO/z2
Y6tjrEqvidPP6FbjtsEHwZuyulnf/SNCZL9j0aUUn8O0IEY403ur9KWdJdKuO9nW
MbqFAaf6+LuyHYzGFXeG59R6PYdDBjrpo8lsqmBbtVWUyBb7fORN7+ZA9Aj5+7Su
GbU1eWTpxX6sWHtYNlNWsZIRZL9lEX3m7jYUZ8Ugn+fp8gcsc3DZG7CzTrmC+an4
fbh3hWbBAIlSYgZKZCMe/DzFkySCNk6/Rnj63J8eZ4JarMFPaK47mOjHNCKphMfG
rjVv0DpCZTTao/pWfqV37pzIFBKf4o7xa7Lx+4g6AYO5A2WhuhiBWCbHLMCBI6Kk
16C8sQK23XpADOg9T2NrS78xDJbGhtzmPTwHcty83H6txwj7S2lhzD32h5nrqgs8
K4T17xUJdFgzDAAa8FbSuG6vHdU24C6+ymchEmpDKIPI74HdcBCy1fh3EnmYn7au
s96yL1rT0mG97Fx5zI2m9sUbdE6VlGbM6E4ww+z91ZBEuFpjOdTXqvGgqwsXBcEs
hcp1e9Xo5qrtDXTHZHxzDPjQV//mQqxn0vtZEPacL/5gQS+wSP7qoSbFyWexM7bu
J64DGnBxcMWN8j+vjFoy2M1RZrRTCEhYwFItKSG8yZ7Gx2BN7E5auURKGoyR7lVU
QiGm8/QYaoh5YRq7NZPVOTDYcjQsfCHNdGon/P7ksvMHoL3/ohk0LPeSs0AHRCNd
YWfPbVE21K0mOwoyOdk/V7IU6fZaBjiML9VoU8y/5jzHAlA0MowEQzEfU6t0gE1n
C8XvCNYyMgEsgXR33ZszSRYtvQqtLqUipV7AT2AGaXjE58pOiIFzc//SuwKtpz8j
pNPPQVyztJ/T4eBOrXUSdYW9R2SZsPGvqmko+PP1bWfgGDajL6v+MtEvxY/U2Bmv
oEEF7UTgYq+SzQX/unN5Nu0AtDK2ivFIXIYVvUJQ6OYGa0yYYgFq9+rLwbksWIlh
KvMoYfvEMblwcL/lm3VdS6Bj+TOqfcP0k9IoOHuLR0WzR0agO2zTMLVr2R9vgV9c
6yHOZ7L/JPbDUcntKsuP3lA7dEtGLDpgVU47AbSmvfP0kjjwS0y1SUyA6kHBc9v/
h9BopB47qTTnzDf/F/cVy2FD94ZCCZrZl71haiecSobXJK/3BWRQ9xTD3IXH84qY
X5+z5EMrs++a1Heu2EXqvTVFkCAJ1DaFKjj6ryw1Tgqd+FwTiDUJ5BJJBKC8oRas
Ghr41BEVbWUYFXJVwV8n/HIkrHcmdGZ1umP9MfPmU3kLzlvX/rEngp7pU0X6nUjU
WeM5WWJqTm6SWJukQwn7NgPzReMd87KvyHwnkU5JhLzvOimZbOdNbe69BhrfTD6q
2lPxUe12OIQis6mMrT+gv+hEUC1L3Mra6wU6r5D4UjpLGJHxdsrMUwqqC1OCSoC1
Vt0WdYdLICqHIo0MnaczL+xqwrkYKCOZztEVejdks0+KHjIbDxsPbz/mh2F73VbP
WUKWWLczfMS+OdrEWjy7MWRUf0JHTzHxrpHH1/FaJY1ZoI4Sv19NmzHQPHmwV7Xj
pUVwYd/VNYAThVvkvdSJobE+yHlGTFozwmCdtB0EmnNIMm+EkSrc8TRTMOVcwc3V
Lcz0+6svr6uGpU2u7hL2w7dz2er+wfg6ru+YayPAmXhIoxl8tbzmnR2kE/kof+Vf
O2YT4g4VCD4DkcZCa7tq35oIZQaW6je/MPbbgcKdCb/srlVfWeXNrlOakmI+OUbD
kTszaTB4adjdk024tHt7PixIgBrt4QYjx7rqmVFgmW1LRXyEnzPYbVd31GC1uESr
fM7A6uirRkJH4TsmWqj7AfwSrpueDFbbKoIfSLQRqfp4/BioXmxAGuy7BwX+t2aa
4JFbpl+Pp/xRpzIQi+VeK5n1XgCzMzrQsXVuOniwdLt6z1Iq9WeTEchR0/H+WH35
54l01ff5II38HF3+31KQEa2HpyZA67MPCLyQERZ96FkaAtvcFLMyURBuog3HJeAm
665ouwEHsXC0kmtvxabLlJvNc3e/GlkoXxRzjO2tz0DFX5ELajh54ycFEUlyBhDH
u6dSTpz8aszuWb5hg8KuHiY3hjAB1iPBrd1Uq6kTDFqsJKcKdSHPIAg3WF5qLx9f
HOyp+Uv4+6gVVFAfVyKUfMaakggwiIZmST+4NI1o4hCTG8IxondRR4mh3FZejjgs
dJYSy5bYivdUB9K+oET+NoJI/tSVTa8iI41LeorUPqZtBpgOYvaF/vSoTq0eE9ny
Ziyx+NZtCJVB1N3kEpsXxNojmqFLhJLm09EX2AWbmRF/uqSM/Mgm5T7+YFByHcOv
7tWFuW1ZgCl6o2+gQOd+34AGsiIH8CAkH5BJxobG8TiCOjGo9CYQxaY8tnWK/loe
VzcFrr4qN4UsZlRNVAK0ABR0VykQQB+QmEU45UwcXFcRD8f1JX4DtWDfs0H2Evk3
wSY8SfjzwgTRCya9xN/DIYsls8YYF/RAHD5CRJgK+/krwcggpmU7rlSEfYkpem3t
0WeRzQI9Lv7yKgwwR9nxZQk6A9lMKrzSPreCSW7ScIJ6v8sr8vWMQQWAyKcby2ot
Kgi98jMC9zT458kV42+z6Mn6jT/I8sMt3bB8P6REaRkcPYedJBSS2I6P2ZmoV8JN
3hfsf2ya5qUSoxUig61pxaYl5PS/P4eqHD9RqGXL2AXsMYGDIQCRH2YipxnQhZkX
GRWSIak+HNdOT4Gl5GeSqKYfXnDiVumZl1ujLKUjml4oz+zdSamlMzr2XGw4/a36
O33Qd0SfOwKKneovsqpIQGtpgbGPmvYTqLBOqTo1vOgXc/gB+44v8c60uTEyEFdz
/f0ioVx5xVjOif8mhMvMNqjlegWqJ0s5sdTwlpeNx/eo/NqeOLNo/3mt8xQzdV5b
Tl/2CGyAQiJS0drEe90f9W9A15uvwglU25xfpsghROMl3yiTylfYXsjFlOrZHnTb
Kp3jIMNh9poffRSMIVrLiG8xL+Ejix8GRvZ3DMNqRuzFws8OMKMcFtSlVToccrx1
RsJDU9vN0kqMXp1fWnwH8PuCKuXdEB+k6BuieIlGZX/iRS50yN3YieVpRlfg2Igp
JBYI5h0JQfmh0j/41R477c8ek5Wiz8XMCM031GatMtrrc16S6I3O9okf5v4+RXXl
/b+SVMwMxBuT/ZHAGq/MOGv1A68Gu9fUptMigwiopQw6F+aGa26a3nFyNsrCnWlO
DAiT4GwgKqozbRW2juolv5Ueb+1mlDY+YDfm7mggNoBZJHjDmF9WF1kaCOqeGJEn
5ceSrpdVUvoqcyAqgfwcZY6MrQUBJuhNb0tHbnsww+JJIvPbz+E0uyDEnGYVtnvk
ZiWE7WkOEqhs8B2ovz8W6kHBQEA1hT9spyCKG+eiv7GEeVtndE4CYyNhFvzIIwUY
jt8oGjivS6KwoYdZKIAeK3xTwdwNtaCT2DPwo1XJM/Jk92XD+ADbV475mcqc/gqI
SxTcMAT8Tezg7c2nCxuL5IwJVpEhyKldXRD6zVV91r63SF0+AWPnE0yXaZpdR2bY
4Z+nw6VipUhDyye6UOK2FASgw9JE48LglSZmjrp+5dF0esM959wV3y4Z6qtQRkbj
NI8rxLOR9FNMGWUw7J3AaIFULSSQlwqWhluvdj/ZLMLUhf0wDM7kNWfLPiXKC8PW
Wv1GIzE19NGADYDf+xFMbT2ACZQLOG+dws1DXtFRutTjQgTNZwX3kRAPFx1OzTmy
jMCfUYeb6Ow54PpLnxcOj1FcCO6zJoLmPmzPly7Ov0hTpVK2USX8C2HfetaQfdJb
hq4euG72885uiu3xmH0Joj0vNp5Fj2J+lx4XQ71ssrc8dbYqZTXzuhuF7lUIy5HP
wXb4EhmjuQJlWFDmfklLVPkkHcFlqtYs5rwPPlJEfB89kyiwCO8g5svAV7+1hlWh
3WBaEA9zwos15AHr1petAz+DEcM5qEB4R+DVQduRVbAxawFiqyy0my64u5W1qDDe
l3QOqEktTpasillYsqV6U2Xd09sfUjm6MKgRkhJNjGqkO3/nohl3OZ46ytceNUJc
bwXLCTVEsqfiJy6HMPjsifEE7m8c773j7we+8Rf26H8nKFUVTnLkO7IgRY+4QhKA
lh2cK4O4grl78wYxpQos8W7PMBcrB5AZPNQGrgmGfR7k+WTy52ybqIDWmoqAbrxK
sNuQ79UvOLC9DTXtY7nlmEO2zkq/XfR/Bi9CqI7HwgM2EeW1vuk7CybCMrsTLVUb
v91rGr21kAug9AP/52NCgRX5R0437w3m9mCqs2UPmX3RaLwALWlUJXV23aA9OePy
Q/qlBTkzubjbG9yCezq6QRQVjPbWVaChKudVAeM/z3dRz1Fw5h5RdA/i3YCgPcbM
MD87cqqSguruv4I0Q8KvtriuzmWSbUXbu9HV/J294zxhrOc3CLyuRcYMHIxTwOQ6
PufUpPTbfrA8l5O7Dmbaq5f1EfVtT5qbh6fPzP3nHchqwTIS7lj1v0wT/Re4IR8v
H2ZbQLAaGV0nIZi33BR3WeRzsMmmdCPg0ubxB4QNovfF9SW6x2oeFGoayQRwUgWq
a6Qmlme/QNdP4SEzOTlz77OMgv0oPyfp3h5IDGE0zM3uO4KOwMfFWNFy/Rx9traN
9ttzPWlkStRNX6nQtRDra/8BKvIB+3GpaVbcM7qbBMQMDZI5DZO7wVWwfuH0XrxT
Tr7j9egyzDJL0REVIWcpOWVZUehfXGCOhkTFLkx20PV9nMLeJKsXj3TN+7JQ4JUQ
LVHEVe0FeKoKhf1HFnh70CagxCJYJAPWLEBf60FH0GsEX4OywXU7LP14ugMb+Y3r
Pl2pjUf9nTdxn8uizO/1XSF1oGfpxQL2Q/DP+hCTHhgs2VPM+ozd8OUD1NiHuaEx
KxbJHGk0RjTo9CTSaXqKf1saZw1JYiL+9KNRTLnkMEO2YL6MNPLegICOg4Kg4fCR
sPG+N93wbqYdcPHafBm+o7qjPzod9KXVWIfSvImg3LtujM2QpDXOzZ3D3hL3+iLB
O01wgR+IKGcICOKBK9Gx9XLNVZHxsdETe3GyL4n395ymih/pH0W1Ry8qkdRoFP5i
LZd51deWjH6H/xmRN++O5vjj3vHuP6lV8IqtACVDfgYo0t+ikqvLm3Md+dzzj27Y
A3jEAaPjYVLflHE29Y7DB0+XpuwQpJIYPsoWyx/7zQme1TjE/UiGRl2ptP3Aobp8
5EjCw6as0yewoFj87HqiDZoZSkL89a7s3LlowUrKdHeYv9TVwddXQsgnGBDzSRuk
09rOkcb8A1e8za1Boc5K2VlKZLutNyZmcoz53RG1I/4z5nhbOJxgoutyNQ9G8Gwc
G52KWshCDZYCQav7EQgiomMcj4wWXUadgq8iDlZxT+n1tpjmu8tVn+vWlEzQukIA
xP30V2NpqX2WVBiwO/mhW1B1sFckb7neI2BnRV46hmoM4FnWfE7fiwpsD5lyw7WP
+jwrUTwwu7VA/+asCBLU8uKFWR35WwO1dVN3Y/C09KdhyfpzZRF+CY1eCD6q/d2l
jtFjhYGvqob0Fayysllv9h/JHyHsf8nhcbla7gyZ8XdrMbA97+3FTiR83sAqemWV
PTIBDGWwwvXNA/yX9JXnE5Vc/oCiOIdBkmeil37gC+Tnd5B9tsLvt+diMeZdHgEy
ivQKhZLog0zsjvxKsk2CPI4IKkfpx1c6tlR+5jK2zkjqVHKuARSwE+ldxJpgFxwr
cK6z16eR0rkhRLIjxT2H/2SQH1tEff0/gdVNx4JmyuuTVrhJrVZtgwbyOpeSgnDn
4iFEa2KmnJ7ugp1seIoDYV/iVTIUuMwEf3B0yTP3nqpTuNW9twOLvYjrtMgVxj4N
mEdUKa5CNAOF/AlgXIMwD1JPTDSnEdlp1kHPUJX6Q6trQTqJpRpvvLIem0EfTTt8
AQdfHMfv2ol3tXcxLNsoYkYZRlidxye+Oce3hlsMKxhZOXxI1hzys+0P+X4STWWI
EqvCQfs71nSgkagm8HeMg3ahcF39Eym1i6GxNx6X1zR2oi5LRZ8ZlTMagp7UCg3R
eZHJY2BMBAHQYky7w9QMwihs0eGuf4/jnpjyr6RhLCemWbbdEWgIGFt6JrZxO7Au
TWrO29pdpxhcfN2FFcf1DvRkld9gPGxpzVYy1CZjg+PqOZtb4ehUmck0qnIYvql0
9haehTp6mg8fnPmI2JNQuUi47sea11Vx4EhduVbps86cVBzty8pVH91JlEQvrRT2
a1rn6o5Ertr+o/D5itzmXNfYcg/A8zLtXO1xuYKrnqhfxeBLCAodGOvuXY74RQSZ
ZqvWfBT1zDhU1oeVJ8oVo9oaCUGY8gHj53uSflL1lpO9miSl1QF0JRxdPz5e5jqn
n2MNN1oSENj0qCBzLtT8WYmr4KolDicdHWm9EwvqzOk20rPWAgneUVa7MtgZXqkl
hzyfc8NgQSpQDDFLnqMSSobnnb1vOAXAWh5Jx+yZJNybtsrgc7umswRP88XpIKfn
LrIWypPdZqEQv8UOOFVLeP1Yv3xr82aKGh7LfOdly4gRJSmSv1h9cPQapX/fRXj+
jY8SCIlKBu5ZE+wYXR7cPa+BMEAkuHYZeM5D+FIZjCsleBP+5Oo7vhRqCEb3u+7b
8RZvZJ+nzc6Ea2cJU1ZCx+DZS1p4yXn6iNRr7GDhtsIK51zm0ZJyAmeGZbQLZBuS
hbIcGdL69mFee9gn70vIPfIzmfFzwHoNquYEsXD4+f5XbRjfuMzDJGPKE7sE1mIv
yl5XX9IVChqaiHomdYEflmF++4oDdHBO3N8cPJMNSC7/iA0tLKyRs7C9CBH310Hn
EqR0HUB5s809ReLbGVL92KEnGEGz1moBDFCPwmHKVeVNwSKxVcmRCMc90kM1uwQs
ZCTLDUzCdpihtdzlWwBqZlZ/hPQU5DsjLbJYbGH7pAbfaMI9I+LJ9xVF4PtE6j0D
fAKECu7ycWZ92fmg/iJ/eYl5bs8iNQGsAhU+kAxCekJvn3VDP7Rb+J7DMs3kLuCK
jw+uIjIWz1icBRvSNunYwG+wu2jynW2VX48A4MOdYZJ9UCRpBbSEmlJt2luqzTBp
woE/E1U8/eeAhk/YEgCL5yu0CsawiEMiZwpXdLstCYg/3e11E8E/YYPVKj+/+wIY
EkROBClMudpTxGWF2OGD4rGHKBlFqWHSMmt/xzNMcVjhDqOny2ebOB1NWSIGBR/S
ZtGyWqhS8st71JMsH650G0AuXFPCmShxqdtUzchp2Vk2B0i2vnppvS3T/CM7MPXA
smFdF995HnB0NZ1nEK0osP7O2WKgNHzKcXKHfW1PbZR6DSwQSJQ2P1VHCiHi3d/R
OKW/vkYib4GkYDZOhWXu8fnIUDBMSOobg74/Vjo24TIaRsxt33MpgW5cKID2ayOJ
ijOGogUdpATJxhL/bEFhHy3M2KoQ68oBZR59qJbR8Zk+Q8ten4WTBfJYhI8X6X3F
IPFhCElRIc9JcJJPwmUzvxJMEnq0g5mkAIiDQAKrMxBsLLJ4YMaPBeQGtdqTwafB
0Lxj6TiZyOMAEGCqLdvHEsF14GQaSfUkB7+yrV3ow1FdwXZ4PVJ+T9BZTZMCLYtv
jqcaHEy8iqQpayDEKaTRO+iiB6KGZ42fKkaR/NTGLsNp48sITljXP06sJHS84PFU
d8TZWeMvGJsCFBvQdOKt07lhV0Ng7Zzldi/hNYPyo9bi2JyPmRIYaH7/gdbkYis6
i21SwqR73dZR+bISiL2cOI6I+5iq2PRzt2sc/GNyZ2IzvPV35jvSk2KYHLrAEkVP
kgtO875wjqADXcWIvG9Mvfx16jg1bvkc1R9bYx8ikRpcGgqMzBYjCeMmLDh/hzM2
xhmF5feJbmULmP1WkfkaNBRwX7SKBxd1RLMNChKNnW9Q7TeHq1BEPaeMdGI0brKC
BO3Gib6PyNYdbC25+2KkDiTRNJQJvnlDCRLq2ExH8ih8w855jlWt8Z3cEN87Ds2B
CAu15d6DLchzyDOHsz8twnXEZfWmPQc9gGJQtsNLjKhzQjj5ZYVkwRAjxs84yyvo
BeQ35UiitKdDfofcnJ5DWBmJ65uIFcJf2zQIQPqpUqblVofePY+RxoiI6EYvAKXJ
u97nUEkoFBZcsq/DRxhFzpR81E22wwg3PYU5yNb290WG7l/TurH1rvbAM0riEXjQ
S3eKoWVWYrMEX7zKmT1LxxDg1AKv8mQXqACudJ7unsTBEXXzMw//mrPhoVrqZGq/
qA7WVOdWnHtacSTrn10cUxJWF0dOBp7lxqK5l3eWbWtDDwuIbMnkNtI3h+TqmIRW
yR0IkhFfMiJz80n9XW/Uei00SJylfNxXT/2IJVe54BcF6V/vUb3tTuctUUh5HHqS
/02saQC7I/kXVu1RKJ3cyHuwgQR0B140a6hW/ZPEwaBJlh3tPmIst/qS4v3h56WE
i0bjvLUlFv4YrK6IqTg0YsDGMo0zeEdiD4/tLeJbyU3JoDE3Qgq4IxAHSd48ct2l
iM36G2Cu89X4eGYBN/9Vy9er2Uc6T2iVZTupcVnA2K20GYj/pZymKbSe+A+Qp4WR
e5VO7QbwQR8zOAgRO3jgp3zm4WVM8PZ4G+2a8JGZtM67GPHwhmwXUOi/PoYGTOp0
dBDej8BqxpNMCZ1laN71BUf2EwyVarA8xJHbAyEHfFy6ZCN9omLxIZmtNltxyJYK
/pyyJZS1N/p0LMthylW9XxSSAmkmeyVN2jN5288jtmJxr23n7u07MNcio/+qrflO
3BNSdL4Kl3sy1EOqQ1UFV+hdEE3peOKAuYpYMR2Q0JQeconYSBcQe8eizxeHMof5
j9bohGNRDxgeeBSe6OdLxPH9ugAOcIazPI+cvn7F8WZvdrIShKf/5+8I8P/eImwa
hwG77i/mjzRUF7+9OEOe+n5FYkauCxQvsFOZojoPBGlylglIMgm6JmNu0y7G+pSE
w4/VjIhxClX3uW6XgLxpXFDGhJ8JmxIdJKQzJ50FzYWVr3/001tyKZtOaSTMkNYp
t+uRFBn2dlN9di6MAPX/F0TzchG5u7dUwNVJo6v32Jt+SsgNL8GZyyXQVuGzPEog
JMBQQkSoHmY9GyaUS+lZMG8xlZOzkabG1RWLop76nIJdo/MyOs2osRITlu7A6po1
w+SYvKZJVr/sZmpkPPuK+y9P1eCyMQOIdL/ihj0GSlpsZtMCIJSZpd0Cga+ngGYv
SWCyhbA2HsfJSrHSuAz/zANbYOBRAIP012hYzYUhPjcKJGJg/W1ACRUddxdjF+cF
vEYXL2NW8Z1XKvpyZk0gDL44342t6aCGRIZPr2vkfgPzCfxGymc/na2nEibIdXbo
zjSoi2yqwzXmRvmUvorT+rwxBOKao1np9Rg2HCqaDelsWT7CQe2LruK2hqypyIuT
A5cr7QLo+9+IY50s0e7nWFX7uL26YBCjQwZwgyWOX7nnuQa6JCnDZ7mGQd/KjWeM
vZ5nqDYl0kvAYIOwZ15A09tP9bk3XoTk4AVrrWU145/sAWkzFb7BQrdHaBNqw7vC
rpejXrb5pkXAAatFFiKYUMoCl9jjLR6bM1Jp2F+kY5swSzVtHXq0N+DBWATPLf/C
hrQTUBwZKgFvek+jjVEy0TXR6SU+Yjr92CsnLrUxqdMTrFlXiwn/SgFtTfjCxPuI
47IVXTvqK7CwYY5EQuwVOax72Bmvg5xdvERVICbZYuGXKBB+KK4GlAyaG+wzGgYT
XHJ39dhCf69sGXZ+z6iKnifItkMV/Mtdj1KKDhkwIsd81ouvJVXfzCTt3ZzVitJf
hS5NqHgCOczrf5eUtd9mbqZCQ7dgwrMHDvq/+yx0qaVOHjilE7p/g9Hyix0Lk+Z1
30V9317cNjQq9I2ldLrtKFPWdWbbWjU9lmJPlTnOo2jVixxnjcGBjRs9wblV1NUv
5nWZwD1/M7H/UdpK9tfZmnIYK2CVg5WvreKyrzs+RycNMTCRZ245pRX9DuogGlQG
JZEW3bKWQtQCi2QRDUSyhd2byNF5MGbVMByl4nFBxaWa3/BrSSRBzvyFxxe7HQUm
wNaId6dndUd1XlDpNS/JXaKcQBRZX5NaU7iz97jpiuNANmCssVNBOo1L2V9UvzjQ
NocQmhESh1WFMClohrMJiFO5TigOneiGLC2U0g42fvQrHdCb8cIVl/wrY4YOhKvb
HiPGh5Sjp0GwdeNmpjF5a1N/f+EeiFfyy5X3v3W950ltwyiUoSXLJIm9bpXDCSpU
d4uNvn1jjgD0XXAUDsmdHOkHE2Jh6jQwDAmETFT3fqmKJvv2BOOsshoHQU+kKJis
5S2ntWYxB9z5sYJlIKzpqp6ZLVT9R5LlBeuCBMcz90qa8cTiUIAeW6IRRcYvdViQ
kLgutm561FL4TfU4VQfjoqQIcNhTfjmy6yVbs3QDe3OmJ7RDk3yD2HgyVJmUYm7S
9gMiiNfuP4OUcPV1UqA5X9C9mqeac/4cViVRLmMGsfi3CiGIRPnhFNjtpODP25XJ
j5FMGWENAHw0w1btFB/5YziFWdQBfmo21+D/MbFToZxNbzuq7j0Z8kwssqqnTxAv
/yzE2BYJlbBAqEpoUHDEVHQaIGQbarekZorrebqGUoigOH7BIXUxzjdl91iJvDUD
trKzaBQ6efFmwaXh20x/+xzDraIBSsY5Byk1XXiSXtQNg6diLktqvld/chqYgabs
5Yr+HegybMhWZlyObzxqHt0Vgw0Po4Dy8ozV3tGFbrk5VJvHPL7Z9QPVTUcFqpIR
1MJcEfxakNG8+HEWxQmuziYOVEr7Xrmquq/Cpsn/LwwKbP7CeymL9+SQBRuUKS7M
q7LB7K1GE0jm2fiNN+a28C8C38YRqcrwFguEhZMjxaZ5BtBCS3eaHsgxYbfPaLPe
2sqiOi8RDjuIDQ+hvWpg5wOinjUsbvfD4fqOURd/86w3YWU81ojUcJUDOHrCSQbM
RRvBs/+N6B0sUY5snKY5FEcHAJrZNskkRPe0yFwjr1S/ZGUx+OnwG2iXUhwz/+B7
l3sUOqLrGIRqyWQzTrD51lu9dJejCjk5ov77Lpo7rLpGvEU1Qenbt9ci/xqyhzS3
vUkGjqWkYCWl3h0AWR7r+S5VvnT4wHaU075jE05o/NhYGNnzFKGW4on4DF8hCl1b
aL6Tp4nvT5cNl7NfTPlSzuvEgagyo/32YxgCxyi7rzLUEShflJL7xF32o4YFd0L8
L6pScsUyvcYXQeQ6xPaww2c7/SFN/TzIkrxuAJRfbPEjK9BgEGdlzkrW5V3FXtz0
LRG7Gqy5f0B1tVcwWWehrYc20dInLhGZShukVff8SdVrQYn5w77/WSKQG5+7aFKw
DPNuhaOrCXZ6Nz8pL0WAcvmAVyss9pE7KBLRFha61Lnmq6GgxtVYW+k4MRKkOb/j
aCNew/VVZ4DLLJy7pslsqMf2+HdqJ2q4CXZp10oD4/piLB9etxMdozAysJBgQBH7
9TCU/84LlOoyUv4OHvCirNi+tj4Y8sjnFLqifDmdTNVbZi+qsn6q61IM6tnN4PQl
zLlxO0VsGR7oGh1seoth3MvaHcSSlX8U/XKTQtT/1CRQdEnJsyH7wBxU030cRagY
vjaK0/yqvDaX5qh7mh7+tiL5OLGNHOjiOdCfAHP5BIEwekheIBf/CJKe25JgHo0L
e8j2FmLCKRjJLy0C68MimHggtqExhz3WK2okr603pPMaD8h6v69W1nX4nKIsEvNg
KIfj4497noZU2CSDoIuvgcv7ZkNhq865fUCft/QTGQYXJkpKq3nhEMkzzar9SXhM
EXCRN07jliextgBvXEjt5ibtP4NKoZ6iyez8ZDhRnj2sYg+Gh5MqNCefwBcy9c1q
kjCr6RvF0n05asPwCnmOdC2dEfhVsY3lqAzB+4YyhcynboiHegb1IeSrGvVbe6Og
NDqb9KuLg/rhGkZfvoCVkKRGJSjHuFIYyXcj24YK/KwgITuxpOhCTrxpDEKfjXLc
ubqbBUNfmXvpe8hsfR14g9/IcBmpEbxiD6GC68HJ+7IQoC431YmXLUX/Dxlo/dX9
s+m457QAc4nTRET1HsvV6E2qSJoCnHK5EGba8aWREwLdxDNNLlu9+hm9J+1EPPlg
9cSMKDDurJuIWxOXA31UFLlC//NiLwPnbK+sfqecgEvxcNkeV/TKQbGV13UupEh1
VG1kyBDgxv+MVQTAe446XSvcFFo03WlEaJmhjZNVbfuYu0ssVRfBgK271a9nSo9s
0GAaKiI4PPsQN4VegIxEDmr+1LlZsCEtXf8WXzzJnjr+E3RVvnBQwz/6eAxotkA9
niAaqhzfYSTwNPsIB5fx1LT9p6pVewI1+I3+C2FoqGOAFVTV2+zmi1HC7FR3CKol
breZQcAwlbIZgVti32QA3B2ItfhS5VRGqqeJ1B+js8PTYv/KEJYOSLLwVh0YtCRE
li9g4Rqxk7mPhtscYb7y4o3g9LpLfs7epypSPCphcfQu/QPB0hxbUGqRjSZDFlKP
3+1CTcy9W67IixychrZdLNjWIdI3uSQ/A50rtqHuozNls5DxqzRg+KL52icHCa9S
MBgsDyhlcNkhfjaNyxd4BRJA1rLy14jFXJfYB4rS0BmoWAjuClZzoxA+4P5TaJ42
FF5vEPcrqWCk2FV0KVtzuLnbL1gqgvI7ggUIDCg7hMjJ9E1ZbK4pROjb6i9cqSRa
DR+42EyIE3NPmuZb0MAhwIR7m1/tu3B3eyclN0xbyP18urX0d9tyLqBxZ2Lp2oU1
cyRgJZxzlChfb80VzvzviCiGInkNUEyJYjy+eu3ttpsaYPbJ6sb8xVTzeXE71w4d
6l7Bjq8PRitR/ofcPJksV1DZyK8UL1tEhR5RB/jGVW5A8RhYYdDjNbG810nmmCZI
hID7A8S8q9TI/O44tUTAvnSndbkN8bItmPEseudbNUL70kdU21OV6PySa4OIzoJ3
B4Kw2ygP7EVn7Rn/QR+ci9AwICyDnXha14PEmD5/fGRxqX3DfU5cJjMkOC3mf0jL
auvb1CKKntlrlRR/Csf8cjmK4Xd4UwNfvtsA3VCeVWJdivRdbiOM8RoxjhqMCf+P
/lHxLWva/DzL1OzBFwDllgeiY1UKwIqqIIdg2KCtp2XUxIqwM04M1rmBJD21LWis
z8o81bfgmneKTpNj5ElG8GEiY+FzRlJoXjZppX7XWTaLrQ6CM8+Fmh0mqlU9Dx1b
4nO4AbJNhd+H268VgbUnLhR+6KOW6GudPeAFpQMeZcFT7bHeoUm5bZKeXOPVpqsZ
F9WJC64uHANRpEgqUmq/gRb1qMu/XunGbXSbHzgwadRX7oPXs7IujaaWQeehMKDj
vOOYDCrSH+zTdvJ+TGHcczm9xt4/ZfzN5tQhXZQMAi9AG+AhCSfi9O5UCblfQIpD
I3uxTPGEKYpoqVp7U+ufcZiYzMGXwgoUa2bZQ8Z5zHN7cX21Oe5F1qDNtv61q762
g+bo+nCLIuzIz13w1D9bfHU3M+hJjhg61XRSbVdopKKHyjOAcQt9QSzn0NRiUTp/
CcKsqGKNmD+j8MGf7BZI58P4EZ8s69D3xDcZ0bgk9QjheAwpjuYLJlWNJDVPgQY7
CikO4fMTTFRp9EZCzNB8aHY/3+/h9UFKJankMFSOV1altigXoopEJbVKDCUJEJEs
/g/fBcoJYQ+GPvTSyvRqzExqUrZ2skjbG6uMAovsjYhnUJuKmHmLSp09C1TgWUo2
PTrnTKO+ciaYSh2XmmbUIvr/Ok79T1N7QelkWa9NhZJd1i96koDAAX6+SXmByTxN
UzjXshsAC6kxPLKzLm32pIt+dbsN4pHSdTNoZWFSInl6Q38CVHJw6X9AhYqJpMY1
zDXtupMRkvU73G9KUwx5TVn9d7DbgHe3H26yVwqADjgXzaYi+Rtgi7W9k7a2B1js
cI+IOrb+1pNQ9g0ciT7LHLRnI3xxK387e8PiHhWynUp5m5a6Ts3hl55YBH6OpmDV
wlqq1qp0dg1kzehK99aKId7lkxIakBKK5Rg3eN199TfxXMSkrZQ6i1+qiCcRbRie
Rt7XwcrsuuGi/w/+2z+jgCSjrpzq5PyqKPpn01dFBoFz9GIwN0twndfkXd+pVSX3
2Wwh/ZkxkkF1BlDOrYl+HWjgZUZn+/NIidV93Ytc7QKT10gIP7ug6BBsWdgsNHAx
xkVjUD9A7bfMnqv+Btk5cjp1FZa8DXMLFkNutjEANy/7LVRSZZ1GnyupaPf8Mngo
qPq4Zt/zvJ2FWpl78/117oJwPDs5VSxhjLMAyvVVfaCz+A3d3faykwrfVV4qxNmC
UTbVqfxjIsxlZ0LAG4pYxQ9GLbMvZf1+//v5BNHXhS9zvz0GXh7u50JM12PPZTv/
e3wyR7YR4zDR+zUy+7WaNrtmdAb0UONCNTBx9Y9WQ3LmXZEXMkBF4SPWrBoz1LZu
wI6PmmzVC7haDhvXldgGudDGMhOO29D/ZKaodeK9gmiDcUpHRLkTafl0qYcfvnUd
Iec/SjqfOX6vM4qCq9RQR7e/VT5a2gZGR9rlba4f8VgbrprXKvWK+d2rJ2q2KHBd
jv7B1xxwd/X1C5QA6dofccQ1VqAMcO0vhZEy+escWuP11EIiQYiNOGa5nmZqxe8h
VA9UQ3ci+HA/7Ffr3U83oe3S4QI4aL9LfmVlpeJLndFAXVswrKJb6QHdvsDHg9Qy
3vKoUsT6lG3NT2ZKOSIt9OLQOgMWLBrWUInsP+Ljm/To4sZcHlanavDXcRkBKxYK
pG5u5NIEsUnY4qes5W9HnnQc+oljKDwDYMYQN8xbYIuJci8PpnmQ33sLVMEc0YBY
9xTRtTVIPPH1tXWsRi9fGv1x1MFam91a8oLw/XTb7FMITHSHtmnieSe/C2Q614bR
dVdT4B9dHJfKUL6qhZySaIv2CyBOcJfJ3Gh0J4CFZPozNT4FKTQeYsgn9c716V5n
dUGZ+zGeDDsvohiVzEYq67JOgSjKAdZzs4A6ooZwjG6CuFGKSGW3/l7PuSpfycY8
HdWptHrgM2PD3KI7M5emYbVJ6Tnlpy5gEeSFwpYU69BVspqR+35xX77wlbuwZune
lLHJvTu+fA14ZyG1iUf/r4ReHaZR05mwXVXKpKieQkWcPm3x+UiGMjvO95X9l3hu
X2lB/vVcxW8v3pkLoRJE4/a9/I3tmJR8mIQ4iHig9U0ZuJra/1yZBFFFx5qcP6Tu
1g/nrjnAKJEF1URUSuf2MpMGAfam64SJanvCqO8RXnEkgp4h0m1+KF9qAIz/QU28
myKBEUWSvBv3a/PDlblfr9M60apiHdMvdIZkyfOL/U7CrGUypvklEaR+KcBnfcNU
nh/M09/GJuBRifaPleMqJNf8DFfTTPcneR4qcwUS6v4IFT+KSBLiaGP7W1lrMAQ4
xnSax8mWXiBAITMM2ndvnz4B7q8jgHwur8l+ekWaokErbCYiTnMxvcp7Djr0M03b
SPKyY9zfu36zH5+a++FfCOVKiW6921Uiuaohz8FXT+Y3gQHDEcyxfuvE5tJXQ1fY
kdTg9LLrn7PZV/1Maiuti1b1Sh9fjJT4jjArfmI7nShUoMNE0JuhRXzp98Figc/s
PFmmhvZEjO3fVmCcZcXe/sbgIHoR8e5H+q5V+fiWv0fTJx9icQEeXYvsIr6ivL+6
0dRbqDy65bFdc4Mzf93oTMnVzxQLeI4Q+JIx8Y7Z5fkm7PQ61PeND7mkGHfFWdDg
aCQVLAkv65I8KWlkkE9z+VtfIN6xCHjBL/OpksWAoZm/dGbC7QrIwrqNxL9BP23T
naGDNJI+IOGc3ILgm1sYb9xZm67qZqtU1qGsQp8GN/ZPpVTzZRsinxw+QizrK/4n
t3MqgTo1U2Xi+HqlA1aY8WLOmYYGivMkGKpcqmwpep3cTWxhRU2FbgZWHxseSvbu
BqTLQ21SHPlViZxP1xxCI5VSqr18mgRQXNEmCgxQNfsGNC0fPuzgh5qqQciWTGx1
Ul9iSdrQDABfRCdiWUBaWlpDe8pNUso+RM9hnIrBp/h3lMn+yy79ioYjDO3qONpo
PqCcgZR5mBC7mhLsNN/3c2FKl7S6frFii1wchKop7PhMU6tdvQqSkxKnZq0eBzuz
JeFpLrNVoHRGsTM2UKzEYZ56vHcVNzQOX143tFHpuqTUdRGwHCO/YuhmOHEWM3xk
pvi0AUB7ltGPbeSUxh3Np+Mz2jpb+tehy9C2CwmC0hhUyeINDe+DxS75qFb80gce
QztHYfFqOKsf5UdQp+NPTCJ9yE2moBiC9byKk3LoUz3lR7X1EpFfEWdulIIGYUu7
pu0/LyD9EeWNEaqnmFsaf0IoYcGoV3RfhBSXj95qhzyEvadrcTGB0zyi61fGiW0j
XVeOHa7YpBiJLFcfVRnTi85Qwrg0/HqNEc3lbYFOEIHyniEto25tQsO/uikD0oyS
ZIh0431MrOTmzC6+NNbB08+L5h2VNJIAA/CfHHPtIl9S2WqjPcN81Ah1ywBHNGGG
oxyhb/GyKp8aPddPyQyRq9Z3KULKLCGuqjj63S1S9QNS1EiO/DLAhuBMKkq0FwDE
vBT2wylgknrBS2469yQxty+KNflA+cGKpYgTyimba6DXva/Zx5Pdx3XUhjizVxZD
BYFBNnfrQ6W5QmJH3E7IpcAB3ssgMMhKxrn0pR6oyQV7Ugiv/3F+DlROUPELV5L1
MdP+qn9HAS4Ryb5hMLrFWKkNMTOxHy8vLPyBpyitEMiu0slo9DYjcRtBy7AWReEk
655zwCvcAFjsdYa0hJwWzSlzFobD+1iddP8PpQVJmCNbRa/5JUF42M4UA4CFT61P
IZ1QKMIs3ZphrYwbM3dTdwD9VVo2KEgCFSZm3PRh92WMiiyPejZyug/zFIhtP+JS
159OwmlTokGPL7K8mU8uCwB+CZmmM2k/UTkjUQ5KYpsxQuk4CmPM/vLRH/rdDNhF
E01nZKQYcJA2wN4RleJpBILNMd8S7t+Rml4pcBquMTRi1eOeC7n5gDewfrRMyzf7
5v49kc9RKjCzGdperevLvNj2MRLtsFKbsH+wktkQz7F/5mwym4dtwwL5qLGfuOtJ
mSTVxBtDxCeRR23DK8Z4LAsZ1BiPTpIQVMsH+aRV6Qwk3b01bnbyPt2osmtC5+Y0
5URhlwhqtpYE/6LRC4m3iHveW+qe7vKstUdHJa3s/4Rou7RUjXsYpRhCZvDwAjUO
hvzurVbD+9TBtY0YhOWs9OEUhDntVCU9CI7wRY4i5qknjZ0lN2vrYCqIyaiOo38r
GsSsvDJEZ51akO69UtUZDrLm054t5Er0nxfN7HYD6tDLari6jsO6eYApgZ7rN+0v
p2suyi7TvksCnQK7uto0CJbpkJi3H/RmtvUl0P+HDj18KLbajH4m9vUh8nmA+1Hb
aGEXeyBMjGjyvdlp3rspIkhk5enbhoddWGAyngjfq6yOwPiU9dFxCERyPQkcsigH
gImFQIGzTI3p/prUmeGPq3SAr5mAG4DmJsbTuMS7TgbEIH5qbUe/IrRlhQ6l22DU
qWLNV/uvd/EUAG+CTDY4+7/UljkIDTNihyVjeg3GzixsEg7/XJrZisZ2PkPn06aj
Dl5Ls5qI2yWHs0QO+WGo53n/GY3/+Q14rD2kqzq3dj6yn9Ue6CGx6Su55AhOKiVc
VTkPkmqPyyuRET5tZL/sey8x4Z2n5BBHrxQGujTJDFuQvOmhkWVxrTurbMVhjrc0
00DKzk18fwcUb9vmrxMPb5P4O2HQTB4+BU/UB/XJLWWNiZjnDNy4YKGParVTG3cZ
aVjKWRV3KA6+zVVPsOQCrEg9LTdM5iRXhvoDB4Yge+2z8xZS48axoDBygEr67Xj5
F5A8aHeE+amcqGRJbQWD5Bs3Q1e+t75//5cNfXPJguiLNTJUoGnngETW9cfIQEh5
bacc++YifUBogzQHcYjoXsXWcaoHuqaYEZ4lDs/bL+Ijj5pWWBr2pvkq6Xm/ggy5
niRyfFmpfoAIKiBaysavEgrOCnROlEwl3wSEzYi0RfIrMupU/ZHsuqt4cSg9ojQ1
ivHUbsrUINYnH1QRI2NJCpT2VXkEF0eDY/J7yDJa9ig1APTgNRiQbaAU4fVmtPVV
aC0npweaUKawGSSoSOxxm4/ofTfNddQdIf5/myIwCx+A0GL5MCLN4nsOPKWTLSCU
XON3+YUA3ta+M+B2nyf7EhJWdQtRwdtJb1txS6LsmB1fX7U3HHAYOwEul2kz7kvs
bWtBVX93vq/bmThAJCLXsN6axTAllp7Nvkik24EwpYLBT/ot8OFKMUVZoh/YTxBn
8Wd0syRE6kZHgmdvASzLS7Yvy7Tuxi0Ff/sK427bhzbmw7yoF+Gy4zAmvZywrudj
bcoxH+01d4W4IFembJlUgzzl1Y6FErONHMVUq3+nFT5NMILwJoUNP0F0SEtZvGbI
AmP8inQbcxXBauLEKFQhuXWLLsI+9DG1AYjkssvv5e/Sk8IgjlIoyXYwVH9IkgBT
aqOlDhHX+9kk0eb4m6PCNVRDiFnFCamOQJSVcnS4Q+Msn7f/QtyR7DwFQg5yfbti
xlQvYsja60BgFvG9Vaium0eeEIaBH2YzohKzCdhDE5FLVIBJImaoYxMouxhJfsTl
gQdY2Iua+44ZuYQvzhovuVhHUWln8lOp5WRNorQEWUOG18VXCFfqwtkLNUkn8noi
0UGLjVrzbQO+m9B6mtfYqEhRjBr5iOi6+KjPEINrZoFb8ZnJ6YEhxXuh/eT/3DmR
OD5lIPYW7OuXg7LELTVurMRaU8ob61wlLpdDjyc0WnPGp8crybBR/e4NKAUTrNJT
nZ+wUk1ati+DaMRcv2aNgVI1yUD7zTdHf+o0bzcgkYks69Kp76sgyoF/6WqmJ4oN
hYzzn5ykbzVLjQwcFZR2z1bTugKU4kS9tuq3ClS+2A9LxnYupPrrWnTTP0AxGtNC
kwXkrrRjJqY4oZy6nBtA4EfWerKbk6E/R+YYPXlF6IZkmcGgSxWbjxwhvBaRuxMR
Uflr6dPWLg7Wk+Fk56aXddLUxCgwkHIJn1BYFSXGqphrixEOIkwG3WrAu+6GIZxU
QFM3aBcuJ1vrEQTohiG/2pqHK27jeVEkdBxC6O77bLsfh8NCO8AgxSoGRE8BHOzW
qXxjEfnuG53zD6/V9lVCO7xQLmPHHpmJ+XVkmiwCCGEIaUDb8WTBTeRxg2+fdPlg
KP2b7zgVSa74sgDwzsZGD0usaXKzq2b2VNaokkhA21/FJ7g2oRee73TQy7WVPVjS
GIdlcsWo0t4gvdZMNQDGsPdibPu5fGq4rL9kVLCPyRiM+0nn98kxo0Q85a1d3M1F
DXppQ8+RN+CtvgIaz5QC3hPoEBJwVpPbq2XBjD653GvVtOP6ikizSl16n35m8yiz
PElcE10IUTVWAF0S3ROpIRHKWjY7E0o3CVFB2Xm+i9PmOOvYdfLkn7U9wIm9er+J
+d9oTAkhrdqJYNrydSjgqCiwA45Nh3uN2QaHyqD8ki93JnLdXBRJPkwyyKRq2igR
Y2dKxjsv2rH3Mvb3wIpIGw1IgMejfK5cgb2Cg6y9QjjcouwZAX/3IV43yCYnnZvH
U9I2mAdZk5uGAehCtwwU9cDE/nNyfWzA8MuA82Ze72NjZ5UwxMnHzH38rHXyUUlS
/ITwMm9Ej0JySI8hezZexyBoDB0vvJOXAFsB4iUBPLzT0xKtpcH7RW8CUwEhmqpV
YUCyxtghI3L6ww7AofUrXOU7S4Arid+o6V3R5+MkBGNOIWKA+l0VeK3qZGCJxoy2
Pxx7TwfKdmatbrRJdb4rGowRUfTyti9yXvC+kp+rEfO+4Fwkmwwj8NpOnT/OHRdP
ch0YoJL4CgGXyi22HD4cWLv5FwD7BzbGN8N26uEyutESE0RgXy/VtADjOsE87w+K
I9NW7qOP/w865VgM7TA87GzHvvnZCNxSTwaOSsSijGvjBuUCntO3Rdzzex5ftQ58
MIy98NUdHIvjvXu9O1ES7CT5xnOFlLHMRYBkE3Tk8qeOlyYbuRf4hOnQwW6XX4D0
5T+DYf92/ZLFp/wzN+d0dLONv+SPh5eTsE1BoGwPnMHFXKU6ysuhoISJ83nIdcq/
V4SynKtCPIymCqmcWfZDXDfXhrE4eiv8eSwaagejYcax6SgJd7gKmVO0+vhBSs6V
wN33TTtYOhl/6/pD+Tp6K8KpPpYqXJkQjvnLnJvbBTFAaloxlOXHAzO87SN2+/0S
9Ul9DyJVCXE1LN3G73dL+2B3P72ZQVPo78wihv3aplhzgT9FVa/ocByQJt86jQti
xh0brlBGDzonO3++bmaSOWFE7lgi9wVQv5CJeTupBSacPdACfivawGHr096/lxw3
vlCovooTRkssRaoPhfaok2MR32MKxmaf9OTJgmixOyC6Rzsz+4MpWZW3PuxF02MN
iy7Wf5cVPpF1GdWzG7IBWPGfB6q7VKoBV5SqaCVfzAYuqoWcEPYvk0c0IvOEtlqV
rbJbLJw05U7ytuHg08GCwdEZ6jCOIisZU/C3pSx3klsG2n7/30lCiutdIPjvqhCs
1a2jb8LfgS1ig9RD8NUagGcGd6xh7RS76ITFBmxKQ8srHHbb+ZmMdzMmSLMwXcvg
rWmnnPyZm6kuRhh47NVUZi8GC3wNGwqII18tzK/ic2kOkmZ46gmnwaNagfyCrVwu
fntrvEUAOq+9cN8Zt3vQQsuQnhAwCLbrzBhFu4VqE3b1dja+MWdy27p9oCC9Udg7
atbWtWIJDwD+AMkLBbL7IeKkkAKPw81RJuFc2rU+TV5/WPiEYjDNRzwYfYyBuDDF
pNdZpek/KIxb10uAskcigpM03NC/vmXLS5PohcemgDRqsTXNB0n4Q9vuCpIQP7rg
xa9helgX5ihbNsFAtMKk6xskItldhhhyv7Uf6XEX9wGLCu4T9sk8fmygkC3gWH5m
t+79KGit4gF9I6UNKZ8oIhKdkAy5hg21snfxaeW3OUn+kXnpCvHCCF+wyhK0sfFT
49UZFbfr+inTktkBTQX5mtiqt4IajgJoBjVoL1DRQ3at22DIWnRuZqsscJRewY8y
mToZOTY5wMazB1qUw6NUZZlfF5Wo1LYnjlJPWE5yXuCdd06Q2TsZWkb1L0a5ATz9
kMA1DK9v1dIv5HAKZbulrZCd00i29W881OhsvNXqCJOjrrsECwlFIG+JjIgMMePV
wD5j1Bmd4z6jLnRYhGdn2wzBhGFqeGY+fFXCULMbJYnOmeqzqAWP4Z7FjQytatob
fdsJ7HwCnciuPiR2OIx2cQmRAJksTbbK21g5BDXd1Y71kQTF1wio5F2qD68qQClj
8pa7s/AYZq5oZuLPGEtaJUH/kGp7lkhX3o7lpgAhRiAa4iBF3pbWB6MVCiCWortF
uDwHj93elZUgDDt9nQFVJLHSZDb7guaQmEloN0J/a14CtR+TtoR0NLlTS49SY8i4
2jgZSn5P5fLFkjKN1ewQT1kA0uaWiXZjhdXPriZzTjiKutyi708DMtH6SDVog6Bg
7xGfuwAazZd6qQZv6eI6TDf64KiyzYJ2mdalqQIfnjq1WeVlMRGb8FWBuEcyoEMO
y7inwFrweLMGHf/V1zAds5/gc++qCoBc+7wJlyYdUCxC2uU/72mr3jhCZeXE4DCb
3VLx7dv0zeHNHOw0ICn7mdd8+CighP76gWE1ycvUyyBTKjCvAPoQSaUDM1ls25on
OWuUqJLKluV6/k9YZT4edulh1a6aAujA3kuAlDLKRuHVBA7PzpL5ic+GYr6u4u2P
CYEDGsJ1TBnVN+1qrIhctSxdunZfwAzlvJ5Th6twDs6WJ9mrx/tV76sX1zEfojPL
HrOGz4aGZOoCZys70J2OhKfmFW6z/ZGtSdg/XOuOONdOdW+e1C5iAzZCxLdFtZ2T
Rm+oT17Vkc9T3anI37EwusR6bcwDa8NCkD3Q+mZ/s36qMOW6smA53gtehGZa/WxD
9DJ1/CSvcEdJNvf63EhOhxV5lMYqlW83KasiUHCgafYvcllp7TFwTtdHZPGvoP93
eDPgvimebsM/h+sBIhUgqBDrZn9KmZmuobEddl1FKV5LZMAEmwtMnHGNRKBJfdXe
Ahlw8/i3ILvBIB7lCci6G1czmEGW4+HliBx3XVSIoCCXgbuoWAQkQVRbs3T7naH8
4K+gUVS9vOTn4Bhk11fq2TnlcwAv2YUFvu0bpu4O9phaqCcCh3sZZyBV5GgW7SBh
vF6nFTOK83aJBnml355Ayj922R9m4sXJemLVR7/lXhuW0/V6CB3HIyvBHnpGFjPh
axBCn/Rh4pEVfehhaCvA1MnOQ5c6cmx4Sk/dKTo3Lnd/1uW5rTy2Z2nV/cH5BS0N
Q1vK8fcJyR9urzaK10jtgokmRYkOT8bfKAEqXTRdq8JSt+s0FVFgos+Ioga5oC3e
qAamYmf84qENpEyKIhrDbVFbRGTBubYwMyXkJFk0EwkOS0YlU2fNtu/Kv+QQaA2a
U3ccuetX1mCAIWDQ2ckB6Nw+9+yk4wVqpaJd5IRqgZf8vyAN12Aa+ffSwxgDgfEF
ua9qtE2cXFD66rvxgfcdD9u+8cwUX7+o1q06Gjwxf7srv4v0QgEnN8zsanq98D6I
2mHFQhedTdZRIlWqCve3XM6cxANy1nPm20ZieydbBLpjnSQRCfVDu7ePcwMq1rem
37rIQrSGDYBNEWJWG9b/kkYcR29zpOnLxQjtKNahhtButi6D6IxnMvJ1Y2y65HYF
HpbXAn2bnBuA2uh4bFY/UnWSn5Zt2R+p8JKfF8fxYkc3ppM9zTwHn1mlpp2awgfr
4QcuHtVtkXLUQeds/VZzIlSEj9T5B9Qbk6xByVOj6Nkt5zYo0zqsaAAyRhK4hIqY
hbKCaUWSvT+e2p3VSdevJyqIf9PZQwwbI9Mv0BYEiTbaurCaUV0Uk9BnB+eg4dJ9
BZQ1t75rVwdmq54kOnUbttV4HZsVv8ud70NE/lEu+O7A1Xbstne/BKJTJv9bhOIo
I/uTbyBrD2c619qm1pINLbFQW1IGGxut2Rdi8gsgKdlSSdvDtfFYyo+9qBC/9SRx
VuQGmM5xmnSEnPQLzIc1jG8qRB48RCJG4zzVUGsFutubKYfwqhdd9pJs6G/0/kaT
pGXx8lUSfs3WoAUWbgFg4hWdBPv5OAPR0lwSxiOPqZlSycDDwdK63NgMWQl3FgwG
yWVuLd5qPZMq1MIbVXagrHtVJHk9BC1FzjplefNoFZW/ZtVbDb/OhRC9B3tYLcEG
5fhn73qNZcC7S6nTNXaEGZTEPn+fg8atEr+/BUAl1E8teYPTbDVKo4Rz5EPh0NIn
IJJpOZs2Q6WcIMOdkIpfbO3HacNwCuMXRfsoM2Jwx5h6TeX5WNjP3rn1m2xt3dvf
Y1XIrOT5uHiiqPg3TuTeQI34zhZA+kmcNwRSf23Xp+3eDxsu9GRYe/ix4zyii06R
uL5Zv1WPcpQH7hmVnFZRp1Z1G8ao02AeOBQXqBp4wL6+WoaFeDRerjcS2JOFwic/
GcONI1HMi7droUHoNyVnOOD1TFjgadrb9iVBxaxwgmWyHfntdzCNuxT3GyY/PpHc
f8fyXUoDv7qtl7e57ouvMzwzrC4AjRLEKr1YjGh9vIyE6o4TJ+RynKWwoViXsVWQ
83ToUMTW8TTE2v/v5dMlx25y1ucXxVbCAnhxVkSrWZ76q1EMfF2QyltEJ7FZsPry
EPCpKJosXj3YQ8rJ2MryA7Bav2e9iUNMHyhjVgi5tlbzyAmULsaKjfrEVdWe3jQ3
LnEQruDOMZ9kk/PLzWz+onzgkVThVrDxITmhSmYRmLM6u16tu9/10A86iEjwgNc+
BMh3JErO3o/UCFWlxfXM2ePGuvgYWDTyu5sGuRGgtiZTJVhvda6nX2rZ5LVTnzWx
+MTFTEA+UUZVjnzxt83esAzpIXGpg+V3k6UKjjpMiiKdnrxy4KCnQXdXIS+n/i2q
HUrhfrYU2Gd5eisRezwYURWrzmYo5o5JhDm7V2IKn9zCil/XzLi4MJ1LijhKWusI
ZxYNOF6i9+hYJnGNo8cIQwHzF9E6S3F/us+eTgfa1Bq2DpaLZIErN0Ta0xJOJtDp
B7OGZf83GNFtLojR1JP/6Meuglwf1CpiDNborkWXw9e3vxtLMQj18aTp73wBjr98
jHx+bbJMtWWTDIgV6De9Grb2vH9ni3fTDKiDdIzhTbS5P710Liqz0CAzxtv7b6b0
Lpi7ZFX39qYMQ/kK/ghHhiDPyQUT03GDOpR4JFkmhED+vKOcsLICYtiQAlt8yRjH
NgbVen1g5HomzHcFHmJAreo+Az5H3YAAHMnH3B1/tvASsgRCSSWm62xauffbY/pZ
Z3mnA2AJns89yiv53UI2Pejy0IBoludbGtZ4oPWQy20rho4DGaFt386X7GOB49Fx
oFQles/nziWL2x+Pt0YA57WU8JsAZ1Yjw7o99JJzshACgBGOXPhKTahZxDpzBAqf
BKghlG9QIjidzkihLQkKXaOo5G/SucbYx/M79QuzMu+fW0IyDUu8QPRJkGH1VqL1
tq33IjAHtxnhq2FhJXZhiKV9ji/LYZm3cAQgQQoPPS0NkuknFGCa5cOVyCkJjYJ/
RgIjHKB7ZSwr2gyMh/m+wRgwwG/0EVCMYbc7/zuI1b725b0EMVXlGQIa7z6ksjgj
MYNJi+u6mB+C+uoCsJelTLv03yyObFXkGLtSEbnSwtyI2ZwwrZUcnZ+lnVIOoGzo
I8oz4n/secvJSrtBZiesk++ymFUUp1tThz84HNUrqeQVWF8UxaH9xviIwPnUhCtq
fwklRCcxsaKmv0yBL5KF85dvb6g18dIX6ij/la4DJ5NGPZ5PTC2B0OaxYmJie8UO
/8Dj13gZ63d/XIuyaq97NoXFq/Atq9ak3L2JarcpITqkjFEAgeAPeKir5mx6N8Kw
0nFrl9IkrxAIRcch8+P+8pRDzyD+uIzFwRoB7JJTe/uouXhkf0sdpXiYfDRKkXVC
Ypu1J3f6OhhNNG1ZBZfzh/iZ13WjpIpUOH/11OsyQi5rM1e+aEky0oPsKdGd1BTU
lCX/8mMQQ8QKdEp5jG7CKTCxW/3A3b9tWaYmNKMilRv4IIvLXRQpc+AQZaUjlsvM
nTtat0RDHKj04z5/KiX7qKeM+gWohbNb1fHCpntVD/mHtMni7YK0QG//nR/JA4+F
EAKt8VqVgQgyCo0iBZurWolYRwub48phRfeBdW95mU97o3pmmfk0Pt3G/S86ybRi
iLANyxvdL7k8OmJK0aauVs4cvE8rW+b2NnSwQkV5zcQ4KIhw0TyBIwU3cJ4sD5Ng
IH37rlNr5WbFlc4bgnYJErxNWoxhlsli4L8Rgia4Q5Klh5AdpCRevQAfkCJNEjw1
vjqEsZto09GTY+m9AuF52oNUYsnk71uyx7x8V859+0WE6cZVEhqZt3YJImnld6m7
HDk4a72qLzrj4zBINWUSZx6lNvgPMEd2ZF+BMjE/R27LKW++7mx6NXHuassYl6GZ
ndPxqGVnAvJaeB0E+gLHEv2iNOVKbFzQUtYjK10Dv8wXa5tkMr0tpm+U1tN1Jf3P
q/u3oUaaYAHkXSrIB0Un2ED5Gr0K7XYt5lTOL5oJdfedmYrRy3JV6dVQ/fcYJWCg
NdBxGb3uRizX0Gw7UM9ifTrKmF5Dgq5epNoy1T5B+29V8hfKCAcfTT8O/GUjTAU6
hnrkD5XWdfWv84Tw+IK+cDzW7Bajwb2htwIQ+acvSF4OGyu9U1+krSeNLdtTEFE4
dhD1FGToJT9L1Ep2hqOQnoXJu7RH6FZn5Pomk5pJ1nC8FuHdAghkI4deDA8WrO9c
8rR4Yvqmc51aT9l84hvctSsHSZRuvnUFPYfFG/K+36xwzBqHGjoUGICUloK3x8c5
t3wDe4WbUOu1+3biADhvoTdHAtufnTaM6e2x6hGPRza03LfvUutF2TGNTjeIVh2Q
PqYfZsRuRN94YUkPpT8HkRnSfuLy4hovKyZKQjU8cLM5w/VTJKcGHv+921MR8HX3
SNMe5n5cNcD0J9wC674uUjalj+amMI3z0ssvkeif76zn8G2s6ljl28nh1uk0j84t
yGf216iKzkJKScj1hHJW6l3xt1KLTEqWUdqFwwF2obIaTfUABU0JXLn7ghuYzs/O
X08YN35NN9sXPUZK83pRAP2pUhn/uoBoHqKQRr5FEGtPO9eq0AEhKfdXgcTKa3Z5
P0Rgx1DJTnu7cq9Q7lSpblhYgBDyOwuz/vFekDLrHWosbZCnQEZ1/MKjx2b9qO3S
Nqj5oTHO+oCXIuK7iIYlrXCJU4Uh6FVhZrJMOni11jSSfVGQ8TQNCpgADQlJQBP9
N1Lbewaz3EfC7yMIyFmG3+UOIofk5Yp5N/KcqAGNq48qd+Y6WBcb3AOoQhlX5ubc
ESieM+EC7QMRWFmYt6SrbBWAEVo96A3DF2dhLOrPpSSMRA067clprgsktiuiLINU
slnsCU5hDAvFKDvwUfDc2U3Y7xXK7QKXWCxKELjalyIKo+4UK7jyP1PPvPsPouiq
npOrpbQqR6iNWcLh4qwOjzgR3eNe2rN8/6QlcIYnXEGwjZUJg6kUBHB/OHZEzDrA
yeV5CWK1x6ZLtwuS3cnyq/Nh3cmnVLEyqhUUsc13JWW+oLJtjhoCxZvxhiB3/G1q
p+Zgymi1eaowaVtFUT4M6OFoM1qO92a7/3XFGOz7NNZmDkcbo4biFPRvPZaGnSPO
Y119jW0cjHUmu7zVdJqLN8dbE0YDnNPk4r9rbs4nM5Vkhz9ncreXsyCmOK4yBvjx
ces794iAwCVE4I1y7f+9E/50BO33Ve+SLGPqlptOKQa1Q04MCenwV7ev9kFw+i+9
i7t+llI8X3QkNAcFg9oMmq3Z8Ft0WM8przJLFCsIGnB8Q82eAxM2wEpcHMQvOAJW
GbEgUGJyCVlhlygRHiXPdxdorV1KBbDackLUz6ggdRsu/vsD0baPNEVk3WQYtfE8
zVDR5rr4eVs0OGcfqjHvkcJsxe2PyCSl7euzBg6GENek2OOLzp8cGjnB+DIuZ5+2
V4AOsQCUmvJux9LTLUwRS49qnCjftYFUJDUV1xaCs5nwadxZN4y6/XnEYMHTM4G0
MZkOrH/XFt5UtunfM2k2O+x9BRfTszijKWUtvLT/2r3iq5WkWkAhUCMG0jFTpWN3
U7MTudIvMQ+IWLCKdr0tPuZ2SvEgvj1ltl2zeeY5xpr9a3ko08mcoUaHHMITLwJI
gCAtyI7nPBfCELUsCOO+/K3g3aZcn1N/NgJpEYzjrUr+1LcfHDDu4Cw9NowZFgES
/8zEOdCIbzZWYBolCTsCSYSOQRswS2qN9ypL4hHkPXBKZfoBEeP7n6EThM69Bsij
O0U4iR4MyB52WqIuAjRtuxRsYOzMnIuKzhD4jlmn6mVOF34wdve34Q3MnswwdmKP
dMGPniL7oyZqA1Ur2Ts8gjiNfo14DFBNTgUTRWrp8vdGjFibfoiV3KRXv6AwT0JE
Sh87B3EzP4NlqE5WMG4nQ1D6nrNrHiA2YLIjQQPblm8NufrCC5ndwyAnAdOSpNoS
WSEEWjZM0BUKTveWGf4RFVwAdraco0Sy3kDIbXJJOO2MYlHq+DJwNyt0HXfrb7w4
ZNfGJatURpSB+pYL4PoDRT3rd7yXaeZuV2ZhaSk5Pe8mvPi1xls1NA0Qd4AVr7+l
otWr3T6+j2fFc228uc/sIEfSRs0NWXF1uxZW+U6kEANB4QR2JWtfQN6Qg+8l4EUj
SNnHUC8gv5AIIcfc+mOJgEwy3r+vLpmsRbRGGxpoPlRQzSZNxpVbVOp5X1Sqjb8T
xXqbAYjtEmIXNEND3k1zllw+PzykW48p/A89Coz+ndFV2pDYEArXcpsw6JDd9Bml
Ys1BmLCKBK6lEQ547cZ8VS37hWWZABU3Qs82QWr9LdBdwvtzTkWfHHD1iG7Ta319
HauPDp7zt1J8CVq4QnOFL4tJFpmdZRBDXvdvOiA+vEOxaaqLGWyh4m17Wb96ZhVk
Z5P5LgdI54pLaaMBZ9QMzbD52Yx/W0NQtLazWP61X/k1A7OU5GqzC2VrQGVJ3GPs
DyzRRcsZKjR45V9lKK4zZpp48xvxY8Kjpp6uvexyYWqCiI//2GmKNf2nZ3k7APMO
qEojKWOrt2sCpPAj601/tCtRzh7hxiig5tuMw8BT2FuQ9zBCgnBIdknXEjTTjhVj
CCQn1bug+NDOyHaXBlXILgFCh8VpjyW6KSKeNv1EbuMHZh6fzSLHaT9TrIOgfgPp
969wZtYVhCiRtxrN6Dj6kswi9Q6iqYxQxuP9gx00HciQRgWFxiXI1nNtIT5S9LfJ
vYqgrK8WWZJj6nDVDlfkfbFK8RkA4b9Wgw5zeg5E+DvrVhgJMi36P5yQSUq7mlIH
O+0HDx6vJtbndeggL1zRJqdnWzRooAhyI2KPK4kCcqknNGEl99Mdtv5izdjXW+xm
mXKP++90Yr2KwAIUDoRVbMmddGsZuS0m8rsBfy9FNh/4DEQWg8PJgs2FPjL267/d
huTiEnQhqn1SaQzbppomKGeDNkLcfQ95PruOnCMPdZn282RZP3u5j594mxHJu3Ii
9zOT40asWBnlA7X4dzjBTRpv0VBWGGTKRFIIECQU7E/95fG/+2mdf+Ut1Shr6Inw
Zlw6y81czPav5UNmq3DnNTN0+yUMrGoWRJZ9cuUpBuAykf3tfNxfTUyn6cz8jQKj
pxBxYaCWvz6h4PbJeK5dez9MqK0fViUSyjn2JEM96IaEhAn1OU2j9hKqfrZv9Nxq
GogMAsEYpMFLfFbMkRMphJ12G7UD5dni1fvzFl3wPzxze4MVUROjcTJlucTwHlRQ
qmSfCiGxz0Xr4JpbjUvuJfRi23nzI92VqYnMrH4miZC7URSa7Pny83Y1T9VyW0su
ztY7wc+8OfHCnMEHu4Ike3jfqOZrYCf1BlouKmw9v+nDsLYWNiidFWhjt3gO1wZ1
1Jv9v0kXwM9tK/NQbU+dEkJPdOIQxG7LWkeXKoyVibhyC0zZ7lvlSL9sHG4AgXhe
4SKNgn0Lyb2/QUFNQWOH+6/WzQuiLMN5OvaFqZcyIFFo/L6hQ0KdG0wVH37Kf31E
Q02xwcInxbZ885X88SWj+9PERgKzr6LURheJIauyFfRBkNG8xVsX1LStM5PzAsLN
mVRcMDXkuyirWHhAAklq7vrmW7TvbphlTJGAYkLJ+RTFow6hxG8RxiTboRl9axGT
MxwMSZ1DP/mTfA6SuTVwkXlrcgnaI7Mu7C/ZTZZXcbxVbL/vm7lV6Oup/5uBLE/x
4czrH6Xi/ERirc4lTKZl+HkCDL9XcBiqNywmvPH9X8a2MQCuB2hHx19imM/1UBYW
MjWX+/F1PvjdJmBzLxKvwOqpV2ER8Xj3R03nB1yihllqMrWrYfXnLPOd+w+HQCcW
rX9OpabILjj32U7LIvK1O+8L43dch6vqxpJ/MxnniRc/FGGdLxITZGMVLnXzGr5L
QJc4nMTKGhthtcDYBjsyl5x4a47xwZcKvB6ZNeYY/ypP31FQN2y1UkPkPecQeeCk
rW1R2qWIlkRZyNvvwBUiDaUU0oaQe81cw/johdBWGDPkGkbaSEwFeV2NdY57B1lh
tsCeLrRcDlNsQJtl6/wKKwew7uXs8K37S+C7bOunoif1glsigr1HLJXp6Pw4L6ce
F1wQZaWs4adCeP6EvSdxRe2vYbFowdlNK68ZBc7FKUo/9DWq5Vsr9whr1DE9vtut
EOn68r4+wYNAA+B9CtpCfAuoOQ5FYXgdDUZQiLYHOsMyzYbc3AN7e6TturCOjBiA
znIOUqBJ0S39EPLc8HHEdUA0EhQs7UtTo+410jB5NPgcRp6m8TdhpWK1hx4dBvtw
sexnwpY4tpvIX3NPfG01HJgg6OslMPfXmBYLs72E9FQgIskkEPa7MfDa41HwVgE/
vCvB2WHpLDXFNrZpTKBjCybxOJhA5LO6DrTvPuJ8F8atwjd5xtIZegw45GteovTg
gscdeCE87em6JGFuiXzBNRUm6nod6qh6iMa7qYUny9nPJ1LFwsXeIYf/iUKtgAMG
f5Q88+LrtH5/N95UOyYU3dxhiVZOO4OEHG96/zOiQ5tcQBZUBLYsVGZBVp43wRkc
BzOjwNd7wUvH8VZVR7OhO8C1u8afwJb0IXZzer2Zmlp0duO4HX6UME1CLpmQhdNn
KkqA0ILJm+lIBHzkjvsEWB3N7nEEVJjkQvnUVkgO3eKEqG7i/6ImQ9/gMe8t7efb
EEiQ2mdVBVoFOg3ByiaRaywzsWSrwY/525r38ZMiNq/mWn8CKw+Y1MNHJL+6xtht
QuOs/7Kq+57LlArVMVmetqfQpY5JNnNCn3ir9y9e98APTMqztfKeZ1pX7Iskpm43
X9H0OBxBLe3jkBtgp+yMPmZJhBiS5vLvx6772GOXZc7nzLGOmpL41jDYYfFoSLML
mIMId4tH5Pbc93r64/h6dfR5Elt5HM453/DulHr4hCGix+XxO5OFTMkRM4+9KSLS
l56ArhdjnXmQFKLXqG9tRTq3Nohfg5/udbZb8cLtQ2cLyEmtJqKBzC/o66gQw6XJ
21+zeqtgEaclOuiJXEVmf0k1jwAqbJ8KwVfgvltykeYWR4nhRtWJ1t+lWzfAoNyG
mdStuUG279rsR7CizKdLEsNBT3CwhF/QQ/ODwav9lJKHYMoAxqufT5e7CNs3z2xb
tMJ0MgO8MzqvskKfaMIgyDCo6dCVFgeNVRz3Pc0F8w1te4opIBKV7mEsIktTC3qV
or414eTd1FG/mrQ9ATm+LvHOItRBdY0XpuG4nOb2OhuRAhW59VPQvsWF7F2wuX4w
J0SgLNqjtHqMTIyAIY15b6q3/G0P7FYvEJ4HDHAlX58LHz87PTw/0emmAIQO0x4T
3OLBO0trfvWe9kL9Wb7IZkE7aIKWzJ71nOu4eZIAkFRGeGbBRlPn9MkSra8alXQV
VeYEJaCowYdOz/yP0yb+VuBTcGOrRTVJDZLT8uYwrqnzHoMswqX0LSddk7geOpbj
kDZjYYb7jA3aMjcEs8Qu1C+Zil7xD2adw1iXLE3wCwRTTLctpzlRy06SBFGkdkcV
erwagIj8E6vIyT62Zytm6NByj5vWa4FwAN9rp+3g2YmPYKk5obEdW+HclO/ou6Ks
c76sNxg9tsqtqfInIcf4E1ESKOcFstLu7xk7ykS8VeQTvU+X9mr3xaLk+3wBTMfq
8bKU+IEmgdpbWzNrM4V6gJ5Jdeho9XoD3vs1LjvfXomGxhNPpYdc4XPOTRQtl+/l
b4Y1mcBUeBi5nsIVivYENRScg6eo9lOu/g5cUMRd78jvEF9C+tEkVH2CAx3FrBzo
tNVVqKQ5MaKi+p2ob3di/Jsnre00WqS6wGw6lV+Zsui4tElQCUFKc+FZIoYxKi6c
3GBLzPUQFcXRQlyHAfqyNasH8Qv985DRs18NxqdRMohxG6aaGc5+yK2ppKS0y9qN
iqJN0+Sjriu/RfbvnNCqDth4jNiW60mDjNUWxU8YQGbtcO5tGSo8sQKbXYwdzR4r
8ONniMfDgsHxxCZ727yizdkRuAhuE96jHLDSPwxjgIWWzREeU1QKN1b95wKAslk+
5mSE9Inqjx5JI4Z6AOaF4/1bg7MosfRMGccJFEk66hit3wwCCdvU8WA24y0L9wAj
01FW5GCI21zFXrekhhmwVJ4CqsCWNFZkaJ3LXKcmr5A3MrwerDpko9s49O9aFpCq
ie4uX+XbILctx5lZwKJba6LSgE4FH7GyEvpFpYn+22IZYSNfqxmDbnzBAtgDGDhr
TEEj1gg2knWJZDInWkUBh/ieo+LyAJXuKvG7l7FbhDj4wEqM7UabUrEm4uOLrBTs
W19lQWDGBNnpQsvprKcVkKciyAgzPm3gL0+46LBPoq8q/7DY0FBeCkDhsh/x4J1N
hAm0YW/fj1jtGkudkjclhCsTqfbyYL58ZoEyRho4Ex7oEp5ukhYcZGUijKX3n8F3
UAjapnvoqjj1g9uxnbMc+ZNhvwgyya5VaPOY1ap8C2pUHjv+lzBUaWD3l0OQyv4v
ASltKwdwnIJkXqjHysFRGLtLBgzUowjIMyjbWta+tatHvLtlH4R5+32a1dYo7s3b
TlVi8b11LuNNblLg/IqnAGNID5UdNHaRM7nsXPw+qldyD8E+KyEjlNw2rSdMiTFe
EKwvVLA+MtBhXu9SIGTNwOJXqNu1qq7BTORxposIFUUMYYstZohlxnbSWYUJhUej
buBQthOhoKtnPJXLG2wrFV5fQwZKZYdQKUKtBmwLS1VT/V3xmP8/KsQcFnmaVOJv
nlrcTRO7U0y+8YsTAkweKGrwhSrRzNEwK9iIP+Z7SbdtpjYTNneVQRgXZRBG3s0A
VbNigk6ewOTYdltWvE5muAXQa8X1FGFAq7Pl05XMaDSQSfSR76oMRTt11XvsfsQ0
oafVU0to1N76b/43C8iNcmyPgye9oNUVwkJoojynFjBTBS13yEQp22KsGw9JBRup
JwJaOsooHcW0+T5MicvwEfBJO1KSN0+gR43/1GmFwkVGu5SFBPwqT3PPrxKoPeKx
AR6aSUp1PEzkidUX3eFxbFgm6E/rYttP0HXpPIOrOvjIp/bwj3JcJjT1pryY0eLI
p3WFFLlD2ZSZl9VyAiwipIhpUS8lTyoufJRgxWVcdxAzqajIOMZKIV+L6PUIGqzF
i+pfE+uBiZ5DTSDDR1o1s4Dewz/rfdmvv79qor0MiC/5K9Ido1kqzbCMXa5NvTci
J3cov9i+48Q4cO0IOpvIEt6F9PyTVQs8z8w6GoLH3g8ckqaUvwsweo4hRAUURp6d
JNTreqetllNUFh3w6aHK2WWMe+e/fT60R4Pi4iDmlimEauIxDIjwxba/JUNNf828
f3k3pUMev0w0w/1ZQlT7VTbrlNPscm0hL4uvaDyp6EmiQ9jS0oAZD5vqW6vTKZco
BS2hRnFx6kHxdkq78ogkbkKxDqQJcQqBzZyo8vSxu0J2JqvziiNtCxVaHbEs9MzH
4FQi6q57yX9HbQ20ESb0AUkOznAZWaPjRe9BQHVzecgTf6EOgvsGJYTSUiM0ky2o
dICZnZ7EH7QWSOitXtPSJzWeY0bRrUJeF8iv+5JAY1laKLkvoST1/UkfuJVA9NVb
yrtMIeN4g5hD1nnLbxjZBWIsMlKZUOvEAXslOArMMJM3JneLeBRlp0/ulFflc3yr
4FuIALBVltH9PcMeCISTLyC9t8uqaRELqjdFV7NLnilPo5rOmJYRth7Y6pasmTd3
rZZLckSZq4p3CDf0eDIi8+sD568FeHNYJqPZFFWli0M4kY2n8e+qk2GeQivOmWKX
K2RMLev5x3MewtpmsAkruAPkFM9sI+a9pt3dHGhkJQY4bqsWM4mtZjsUCcL9D+3O
67ucFReZs23U69kWHGx6pXpTWclHojEClMQ3vdPGG2cvLRiK+LP7yPcCIIZkdHbx
uRmlpwcHSLlIpmTf1O6VFZwQdc0tUdlnQku57398zoF9B8cafECsF1AWPydy7Wpz
m6Nr5T+77KE1cLmzYWLRX0TqSoKVYSlAR3TIJgW7m+qoOITze+QHCSTgpOlRUCcy
9DY6uqFJSO+bD5FMM+XWxFzZYM+jnqLUwLijGp1mQT62f4vzE0u7fnGHSwzlEh1Y
N+7rQD+ExsK/3gN6SjCsZ0NkSIFeU/2wahl8fHAl/M9kOil8aXDs0cProuYBbVFw
n0hL2u8CcDFzxle69FCj3dGo2O+MzwNN85xEYBDCNCk9dHVZIPzkRpZ0vr/SA4k6
mTs+7QBap3YuIP/m5dcuxALWUG8bLwGHzpcDL4tIF2Ev7hakgiFRqu0W+noSXrPR
hu3Qp9c2HXyZBqdDXmdgopyJyciw4EHOD31DsGJhEWCIhHUmjTk/WJ39LcaTksxD
mD5Rv8eOuvvtKs/tehnHV8joO31hQFuwJ9VUp4rW/gHzMhGBZcdEerYLmaAuCE8q
XB3dBXNU/HwhMsKdhFLjMQD4YF3RJTn2JweFew+8VUyQCCZFnqSCO3s0t1jZ3uNc
7PKzZYJgZ4zKO8TWuSNmQRH7Q27QSnLzH69QfsUACvo1ETgvh6lNHmS5DducjGmg
5Gig6ZozvTpWowsnPzfIENrOa8ACX1811EXEp7byEYsaZR/Uo+MmI4MrbBPgjzj3
jvkKS9KUjB9tWPNShCzmNkpWDUQaVKKdL+nKPzdYjhyillg24DbwvDUtHtiAfQyO
CFhKLPesGA66twbM/JY95F8bQQJ4EG6Oa5x6lJ04U8Z16eGTmynDCq/TvhUladIH
wZDBU5+K5cbsf6btrppuOB1Vhe0Duw0AGR0A0Umu6b3ESl1Sq43xBB16e4yReN8n
BX6NBbYp5Z8OM6VW4vxDdH1VDQdQY0+QMRRSnvse7UxYdwv+rjmSBRm3CKqmS2D3
L1LO+qIXaL32OIi9cv3GhRYBWcSXnv13gz1VQVqkL1TlSY4ZhIuUGWUMv3lebgKO
+EJ0QEuC4COEudnhU4zjBNXXBDDaqj2Mg+2GBlVD8mlrhhRC1l2dlKOjCNGRdV9H
SIzM2SA0McF2agQBtrbcJ3TodWQcByu/Qz/V17cDvw/SKCtQwT4RuHdRiMgSylI2
jwM662xBgAyIUDTJWC+ESDpndPzwSBeYx/Ilk3PAGByffZ1+SSjac3pTK+DT6vYy
vGK1zUh68F5YE0rKPr53V6J34bNygbZ43hh2laje7KMkRTxW4Nma3qcXDl17Bgvp
vYl/z03DmTNYBFxY4jl0iiQM0YmuAtzfT8moext1dHmyeV9IuEgDqTHj7PAIr3ql
9/quGKs8q7XYaVDWW0lXPvIaCdWmxEVJ7SUa6/a1r7m8ViTcAkuCQZXXUaBzHU+y
AfMiWBxyUFUMnmZbOuknCd7gg+Cx5fvCyL94BJ7v7hiFel6IwNtXxMRlGJuqpRVH
C5c+/fJyWDn5zLBBfwj1YEO6HOCLb+XVles+RUBesjLcgWJPm0pW0BASmNf3V0Hv
Yf7EV2OX2dtoXeVHOcU4I4tk8KWaMYh4Y/Mqu/7vXmJX6Z/8S3APmXxIo41UTbX4
MWtgcZQvit1w3jWLSJjF5KT7h5HEeuectdYBx0L7eP1dnI7GsPODPQsaCgEZ2JXH
w5I2iDI+7yCu1KHrM79KEMvGRTvjlj3f0rgDnZzYrHjg7vZiJi5mBxc3Fd2OA2PS
dRpf+AD+lg+LNI4GR7xGesqHtCRgbi2liLeQw+slTYAW7j/aLl8CmQHhl/AeRQXe
9cXin0Cy7AjNVJ+h+aB6pElCi9R32Sw09s5JOsajYDaX8cvrhI1ENqXLUqsz9iNS
pmXki5eEJWjhq3F5OQDGn/BVzdzVAB9nWqkKoGN6cWLv5yq/dHP2LS7yR5xSdE9M
5bO/XsEs80ZMY7ENgv6KBOf3NQNNu8/kIC2dm9rvtxkymRtTNB0NDT+pGr+TQUAy
9Ghtib4p+VaV6Jk2tD1N0azGfh0Wbg/Z04/0qr0x488s2A4Qu1W4q7YBSQb+njw+
loqDltHKKVQ+glVQh61L6K7ETFMnSsLghUaZomucVFkjn+ySj2mlA/knLGpMTCdg
2dt/WGJct3+eQNNQy+3iBRubMaQw3PNsLWtHfyRO8a0sHDbggD4DKdfTso+HKDlF
Y1/YyNSUaW5wxSdOtkvODYHu1jz1avebmzhkvuxTvB3JTZ0pO60BgXgcl3p3/4CF
ep3P5Xi84+i8Q9EASbvhUP4/alSuPY8ipFZinnmXIPiV/niNBUa/GEJzRwygO5tb
XElDHrq/9rg8sPjg4ij16lmKuJgO3CI0V7ucjkgXVC/gUoniM7e9r+OWMASSI/yY
sbzaqvbmIw73wbCCPi+ngs3NZcvIL0nulD1h0ZyxCGt4A4f7sH3fQHpFPfIrWKL+
SU9JfF4nlQnHtncbeeQqRSfndhVskfeBpwTHZb9LoZwA6hqEhdtqfHa611itYDnC
NBZluHn9lV8nE/GZHPRN8PX08LOYwPuOKL70TgmkUeIWq0VPyeuOw5G9OPAtfEgq
sYUXBEs6TkfVpMTDFyMu70Zi/aW4mnpfLN9DZxngPZE1fVPbprjinbYeM4izHcoB
64UXaZwHRSNnenLRfQYeVgy9mN1dV9YBCeXkWjCa2nTtf4N8C3dib7sEv8Ayy+Gx
+E/D+3v7W/42LDFiTbCy0n/kd8URdYKg3lPeaRz4lkhJRBq2+NEfO5FZ8w0QFtSr
6HHldLNKlgCkKxOdcNoFgPYZLvOM9heHWfHzqetUtRTN/wZaDKBLLDjVSQo2U+Wp
vIWLc+uOrtuy3c3RHmzs2s6UeyUBsfnMzOkWGW2g7nQbrRcRmnY13j33B0czoxg4
XgPxnQGlIIW/eKTf01ShD04SDcSAXXt/0/irYqr8vJn5nMKiHAxN06FbE34OaObZ
txm40tTPk/XiwiBLTPZAsIlcVCgeDG1PmoSHPbbWZ/SOa2nK+7/4c5WSFQy4T8Xe
3UMTFSCmO6/MUhZM4ZaYpNan41XwRtgLjl6Rfdw/3AqF4hRJOELXUnCcR5WXiIQc
gHn/GChyW85LLzM02MSgtLOZOfoI+pwcA3mv8STJRK0ARgf1hIWQPj/2iBWPh7Mj
P/WScYnLcEE/daXupZ1lryVmmM0lAbTy5HNgCPlJO2CwxP8XE7ZV8nX/dbxMVYFO
8Y+VEaFAgAHVqBZiedP3XxdUxMnrb0BY88YjUCs2qh7oTvNnLA6DHq+i+0GRP47w
HkFYUvygjoqNRe5cKWvUfUn+C0Nw3Qj1tShRKDd+E9P+mrA8VRmPx52723dIJAoT
fynfyk0bDRtUgFduAzAZhxYUMvv0uDUNKH4LJ0EuF+N+xqINLmQF1r2FdX47QjQe
MloAN5X+lkwP2ubcwnQL5BJ5eEnNItdz2zkmwIoTXhrznMvvQC0Au9FHadmMa3x8
jGiWm7Z/ChSCqMYReymEOpuJta0689C5cZSQOJTCAMlkSJEoB8ce4/+Gq2GRFNYS
EjiqSMjjvodaGcQicpuyK65iQ1KbpJAQyH7pvyK5NFBjB/I9O2jJbQcHlBkyluep
nKSvRDWmqZqKqtfjPYAbU3nZtptOmfviLfzAsOSqtOd773Eq0kmFZ6vv5DozIaYt
XdvrKsYIxyzc2fQN1UQ/SlL8Usrb9Q9ejRPiZ/anQAbU3gBeGAP8kv2hGLmeGavm
h68mrmz88cU/thhSQY4WkBhd783bq/aO5MrvRr2mI3eZDBs8RAuVw4hCyGusSJt0
ur4R/9yIWFcn7M9beyw4bYIrslejOmsjn90lrb4Rb3BmVwuKSjMeSdjfciVWPJxP
ErBEz944b/0U7bCbhZZnvSi1jZOCdPV4N0PIfrEEuAzm6/l9xWObzx2gaa2ciuwt
thuqajIR8bvJTv8C35qDU2CWy1XUlG678uW7wmfTldQt/a2zCRnCaFmLsIWuEfij
9j5amRYiFbEJ2p+yLOyD7C1ZsDYJfQeRBTPbKEQbCqRcHgudmD46+h9u8yBGgsJV
q7OVKh1JLXPWjbxgAk1BMAwAfUyuKpe427cNsdOeHF1qp2sREkf6/msr8uDNzVxu
9uPOeJgVNb3isOqzCk2F6/GZpKOhfxPLnlozTUV/QMHclZcHh8rIF4auKGzdi9qn
L9bw0DL8RJLLu3TkKwaiBSv6vE6nahWTWmkiPmyyZ00oT1GfisxGhHH86GY5yzVt
57ioWloWhQb5X4kXl36cRb9hS+lfe1NO+NqVLFaHh7Yd7db1uaY0QAd+igl/mrFB
+1bQT+6HieFsmDlSceugCfaD84xR0n2an8D5ORVk+x/uhRoRjzU3gUGGreXbNI0S
zDNuj09KBBgimMdQ1GAoaBZ+ZgFWw5FKpywngZ+P0qqXC7Kp1rH1YkX+DNhvPwQy
hsxc1asHgJsHHDNsTFNrWhjpZj3iXiI3IHD2v2FS4CjEceqHjxz+1Kl81zYLyJtI
cgISQxniNUmNHklWedlfVEkkEZ7t8lntId9iLK0TFd7fQzuZjRylSz6cbG+Yqm1z
rWoo3eixWB8OqCZCj1dAH9z2Hf0z9iHZZm2PU+nh9MEae9nI0pjFF7NXBTxoZe6x
8pXXN6MqeGouO1YH1y1YtkpdcWpqlBoVoY2Muf2WL+l//XD9BlV9ALlSukRTDsVc
RgmoYZXjYWOBq9fib5JCFaTLFRAlw5Xclxp0DftM1DdqLQhmVI8diCFhVvvRQUME
ghIb8uAByy1LzVQfcB+t3hosNMhTFzmwIXgjXCQM448sTS2fEYd/fZOjV82N7XLP
A+N45em6DyQ9UmWiFU4xUB0lKgO4+rMIEXhupzfd/eF4CVZy/el3fS7dDfF2tnWs
xcIRCPH8IK5DdT73mzVD3Q/V1daqCrPxXVeZeU/es+vXHI2uoxK+7ug8pML8Sxpt
ntAdV8NYjJG1H+V5tw+VHkdqdLkSy20OUcfdR07qnXEHs+spsGgFmddJDsXm3piD
IAPcVvQKWFsw/nvu1Zb51zJp+K99T7dRsG91sOuMY5dbfyigFAgcMs/IofhcvTFr
KV4KsTr9sNswDEVNgvTxw/ky8PdtCZxRI+rBv41CXyLH3+4eSqPyc1HP8OrC/KC4
cm7IktTHAWI/clRh3atJcBDUGLnUy2ITuvFPpo/9ZuIS1vIoyB9Mav7/QqD3YwTx
tVZXEBO7Q6MWAX8nnCeQy9rLUhu13xv4k1lsmEIWBONNPPvdDg+pTU47Ktwl4Wk0
J9+7vpNLsL4S8AH0TuZDFQq2rBz5Wo5N5mz+b8pF3Mmc14LIoafM5KaWg8A4RF47
vg3MUIf9fKh+59siZZpsWem14ds1XlNMmyKln5GOw8gFmgAzett0WjurP9d9ReDJ
e6yHMSdZQxJJU0EVr4Ybgg7ui7wMmmon/HKqiQgqCWDY+MdUJMDoom4JB/xCtj6V
xf2kgrgVnwtKuSHJhsz04req+jt+URZpRyDScA4XGk5yNx3U7uo7iOkijWCGCkcq
z88748EFjsgVgUyk5Sy1NHNfZKtAdqqwgUgEPBt9zSl6Z0Aohx6JKaDfVhhMfXm9
f4My5AdNI7i+TtSWf3BdEkYEEsRMQPF3LCTQDDf6ahmtMKMMHoOJ+cSN8IZGjj0Q
wnC8LnTAh/lUQqiMUienYbJEicXQ7Ghxhsi+0G6g8UTkwagcKugDEb+X9MxD094F
cNfZ6AOeMY1e9Y/3uAPfqxyHWoGU8UGXZ/KCQ+Ozeh9KTuh+KcdHepC7b8r70yw7
urtKPB2SVHqxMKmVIJLM2dID5KOi17qSjTSHe5F+jKJgRjyW1yReiRvXlDev8ArY
mVKJAhCeIiIQ6Ioo6uPnkqdkvx2aPOZirQls3CTANrctqWtsdfH0UoywSnIxe1Md
tYq9OEsFIp+g3t5ov1inTcyZ+n4IYN9dlinCRMIWDRY6MMzPNl6+F9vcfbKMZJ5p
QO2SRrrBMXntsINnDQNRNB3rN7eDbRV/9qiBIt2Lhpzqdo8rgVETQp1c26jqqju7
Drwy5267PALJJq3A5h5etCXM/wOLywkekZldbk0Y3I+e/BUgDPS1seD+PiR2Z7tm
fg/y0sk4rjUGHFhsXIISX9ltXuxtHFXlmV3RMhrLFqdVXRofpAC10UxZanfv8Od3
uNKLKgY+bzVH+o5UWEP/UrbJO6Kf38FSSkfdboeTuc6jWvLxdYYwPBQ100ugoFV3
DUPLA7bI2j44kpMs16jFrtviG2OIbytDDGSfxtXWZeQkyIV6vWsH8bgrK3bTY+jJ
DpPrsZVSUVALyqMFuUFCcQcerYOu+SgXbCTVOgkhDNQSxdUVRmw0NbdnScD2EcPs
7uwkWputZQNqBkPLwbn0AJZFEG71M0Q++i6qdFXA89sBE6+sJQs0+XUWnaATwYWm
oY79HLxAgCIMERG7RMMvVe5HbHfKyfjgP6B+7vprhCI3rBhcndVtWR0fE7acd3qP
SK0eC6bfRQB/kDD6/zch+NQVBN/OZ5OJ7DxJZ/6U7W6wHkvPBYNS+yHlYXQSt47o
OX0wJdUV7XJ3OPYCsREXFCE1AB4UCACAuGAzIj0DskKwcw3aBbwU/fsqtaKrXrlS
sKB3hmiSkh5RON36dLpmn8ck9WlBVCX8NBJpJueDNAJE/DHDwJrUsvoDVivV+dMV
/TPIxBltRFyn6SpilxJc+7LW8Vwm24louWhYQArqDD6dRjhexOByzqxGu5vR18pN
V2iL/c+k2wIhKlqSQOgYSkm3yc7+hPLUynjNZtrHkgX3lN4ip8F9X+oH9L0qRgLW
F5u5EobWPAGA0EOlNiXhuxpVJ40QXTG2e4976C0IbNKP0bVdrR9hN7cZGGRuEvOc
V5gN4SpwnQRuHgAabZZPzaMd9IaHd2rMWpl3WkCDI+B30wC1nuaRtrCedHZdqY8H
TfTMSJ/zrCoJL7p03lZqE2PpcCd3PUmrz3CvDG7ZDpCZIozGikUsQRWp9SD7EHD5
jsktwUXp5ozFj3O/pjyGt9qG7jUgZmyyWAAmrzDj35v7V60M3famxBC7TbU621DA
6WJUPv9jPRy4lsl7bHmTslWq125eEdUJigzQ5CYqoSSRGVCUfiIc/ylNOReJlVDC
JDjNKop2rBZqYBf/tfQuE+wNXSiCH5v7Q0H1NlkR7JGUu4pr9VjXXIZ5o5ZgbuoL
tyUX1pA+NM+Bq3180ALIuR7+t2xdGdJCGw8jj94U5DRpzdYCdFGcbs8PyXs+Ah+g
GyzWiOHwyqEThZeIq3acNZiw1U/YbfBAAG4KbuS5JYvK9IebnswmQ8cG4IlJFwUB
6V2l5cyBDv03Xnzn178zfWUw+KotWlDJLxgB+yX5fEIkR/gmm5F/g2ACFwOBgCvi
lxb3pCYoovWQzHd73lcRcaS5uunbKjMQFBYOaKgJPVm7+54Jyqw+WnrKPaWnjWKO
A7xUjvFvoCvdEC9WS1B4h3uwiV4Is/rfkqUGRmCuobgbqt4521OqEwkOF/7TGQdU
serUhdtFOTRyzBZdLKhu1C7iGIduJB0/+UyMVpl8TblElWFvoQY7L+aBDkgf3u7C
VUsJKWDMDrl0QsYfNBWnitv5CZEDjfrLUQS/GFWuC9caat7N0gwKUZrXb8A5ADAr
ERRUPwwGzcUG3mHThswzINayS/B0ckpVX24rw/RHyQzDJYS1Z+KsP41ROtHLBPGg
dAAKBUhClSJISI9ijoMbCw7C5ngLbq7CJJGw2JzIVSfeY2kwKaFxOwyjEqb2xBRV
+L54Kf8S1GErw4Hqt8W/M5MzF+TIw8jEZkdNCU4G5d2RnSg2m3oFgdqug4bpqWuR
WtDJW94L/BTt0/XTqUZdWkwRwI8V2WURde4WxffudZktkvJxdGE7X83aVy2HQOnk
MDQsuNEPCtTg/uRTGSBzbMKDDBKSNbQqzOyHjbBYV5lVG+ZpjE6WyhqTeqZU4yaC
tTXQyvlYXYCQOuRg3s2P6yOXVlwNpoNWwdafAkhrEBdbnV2xb4Z2TqIf74sgzrCP
Q26jnetSRUvfxY+/pPt2DlYFGmGp6T2NIceuSOQT6tRRsGH4Dn5xDvwQdTETDMam
jdsm/bpghvY9vMkc/F0f08XLT27dWipMrQUXZePMe4s2f4wY7IGBKea5SOql5R+H
2+vw/TivpzPwjUKpY27W9ZRkrcCWvAVSzZAODbVDvM9S/fk0TuXaw8R1cbvThRYp
9ieOw4hGSi8WbDKGJS4a3/+jPnD6kzk7x1Git8uIn24f1JxFUnQLT1KgXoH4eMH5
GGB8xRUNLtgGpex/NILGSURD7vnTI1JpKYetwffQe1tRJzkysaDv+2ATaVQ1uZzC
SBU0ir172r1uRX5ci7GdDpo96VYs9za2hG1QDcLmf5oSrUvtv2Whf7HWxcrr5qNJ
dFci8xQbNcVL71rc70CmyxmYD/TXbtDgE7HjYXxu1EAe1iiKf9Dge5KdUws95e32
UQZoNpvv9dbx2qly2twLiP+/tnULbtX7l7b7wguAo0KKUi/vOCR1Bz2nu2fzIFX4
gWDNUjl4gENj17OjDzC6hlK0A8P5bbHyafotCHsmTV00TpnV7vT/ufTlSYSb+pPI
9TCQfOn73ZoVampPfbCnliiPj1gbjedjlJjsyp8BE8Sngs0MIKP4JLFmcukxnnPq
SVZEx88O6fvJY0B8oFNVvC6rsibX66y9ve2kt2mpR0L0fkIdN6LxScumbny6bNOw
wqMeVIBSSkMies29IrChg6UxpUJy5s1ykOXtDyF7+I4=
`protect END_PROTECTED
