`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ys/8zWJTPVb9NuYS5Y14A1y049/w/xpraWLFnQ6nla1g3g7LK5AaCzos1wOEz8do
kXAVIy6cFf8py8VkUnsuEGRa12ugWjKeoDdkd16dXb8o2Rhb2zfA5Ai84NSCuyhe
6dz2FB6bxFLn9OX2fdMu5d1APAnHYqIuxmNrqsTHhRPFwnRvjOrsLVlSPqiJ5oQN
c9vrs57+LO9jvupmejjoPOkdFSMB3X8sccdT03NshOpltM9gpDftwPgLD6IeYSZz
lrOc9sBfZFRaOMbbvkdNSuVY+NRMDDGjd2mfeqciht8fTjW6XMd6R6cs9oQdLg5a
U3h5NP1GEafU6m7Yr5xV5WSmxIcmMSCRf03PmKUvWwfbw6JTISTvmlEbSWvJC9a+
4Elr2COJxVLMYo5VENtlCFzQ23zmBrvFVldFXKs1ZACI/u8qP/8++ai8kYGl2Z7b
qOo39S0jvr0E3uVT/NjA6RNOrjNVInHhGSWioNWAxkKCiLgIs+sqpK61cTWdUYdl
iVhb22OlOn+tv7XmnnlNuESbqpgo+wPb/eTtdiVdSaF+2lJwX9W1t8Ew2oYDTThr
JIctXraRv/AL7Y5ZsONx/3jTYouwJObg23x4WPBmAfOfngZ8h4Sgq84xbG7axZdo
Klll68Z5EwIXTpIFJnvfvjDED7pCRenYtsRCsXumE/w1s7AZwX/aPOjSHReRLyrw
8iFtOzxYR0HccGnK/lJA2FO0HK3qp+Hh1n8fnADwg7pUJ2cvHUVw33QhaBWXOVtl
7g3J7aiAsbErzqkyoDQySUqX1+N5Z72OQ80ezMtYXe9K6Wzai9ePPhigq9Kz1Ahj
cQAuNFP8StIeV9HOBngK/l49NC2Hc6w5eXA70fbJ/lTpynnnSa2e1jQekF2AeGlC
UBGXjVAHtJM1G/tOta+goLA25cKAQxg7+Si+wrypA9B0cW14gWh8ikhPTs0ds5jR
MK3qgKeAEl2jeJByir1auUxZkWl4Es29SfDiLV9G7aqXxcHy6vrleyNRF1Zdft3Q
g0RRCj10wQ3oQBkCG5fjOEfEUMJBIlJkFPISZDH4c0MdSVRkuz//EqYgrnQYb+wD
bDpQ0earh1FSdAXBkAgNIaEmw938hHu5hSih4uEBQ8OuoSXLaLMbtBbA5JweKqxJ
EJcHJA6xemZZd2R7KGSCO92bn4BXYT9XGakrVhjNKGr7QfnvaMj7DumUwRZYjHV5
t9e6zDpBuv1vEssEP4CsDAhoHloiFS4qEiZixVI0dfd7Xb7uaDALer3kO8KpjH1F
v9PpPZ5iio92/hhmAG8uACU0riYlhtcF9OGnRxHmlD1seR1ZW5tUYlI0imp1Ny5c
gxEnQHc6ClGIa9nyuwVcoS2OyYMqe2cLqA4mbewGcsKwMGTv5J47qEoNR84ehPPy
KqdvjMWQ4675YoxgFMGuUmc0/zx3qL+eKRdiuFgVTx95/PXbBfy+FxlL2ijXMoKx
WCeLkEpaUby2Z65XMelXIcYm6KLjavjrdCGrbNngE2cxMf6xZrlsZ9pOrCn3NFC+
buMiW2n1y1XTfDJpQqj4s0o+FKkxG55O9yRvuWwd1VW4HlOgE234gQkTXEFskeuN
R+6dV+A0u+JLimJlws+W8s68FSNp1qt0sge+WCDVVzYIHfiwHGMHGuz9PDjnX72v
qOMkCNLUF3aTovKygeo10KDhvtXE2a+xc1wjEnxWKSxRKpIdVSD7Fx/nymKAX3F+
tk995/NY9QdENRRU+ZmLRaOM7/UOtVeKsKBr86AiQ52FMz7/NNAb4Tf2FXl/2ZiC
`protect END_PROTECTED
