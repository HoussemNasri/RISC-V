`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PWly3mbxj0dwBoNLg/btkzbqUwBARMY9vQaaImfQNIgCssEh0f6lEXmS8/5rwTJJ
kzwB4h+dTk7xvXdfDyQLD0pZVZAO5dOsp0TGnMuTBRG0RMu2XC9hNe3AOu1GvMwm
fBMhBBhwhs4Pf4OV3KoA3pJkIw4ollKN9RzKkjlHkJXRbkMieQqyorvN5ppAEhwm
soPG6Xzkr5o9YQq/FPyru/p6+UgNLvtDpDwLN0iezFazXynG64bRMI3RRQxtKw5s
V2CY+PakbQ2EBa0UADaVivy6peHhTYUgsctl5p1KJKCvq9Sh6tk210mybDF+Wkmb
Brakf/dAz309EBHp1JtlNOUrSp0qI9EX3HcM5p7Ae0bw2Y7TR5mBCvzTl5Nsu/Rj
zgejtTZysmvIgHdRVaboO52Opatvsfe+dbO2hyCp1iwzXia3NUBFichn/+XoOZYp
+3CWchCqVWR5TSOVNW5qRI85AYEZskzrrgvKfMCfwpQH3Mvcj+1a0Kh0G9WRQxug
8yWR0f4Vp45IU8uc10qiKkLmLQgGghIZZp1jj2lFHQ3/pCLIMMvlXcGwhOxE6x32
iqmNgOPysxZSU5GEkhRbNA19edOkDufTvgt0lYs/lR6GJT6ZlyEXJlE4xh2yzQ4R
WqXhaXCxMuyizUCxvoZs1ASBrdu4IkOdzW6gfxQ2ei8hP6Gt9IDrO5FIH8bD0YiM
B0uOvMH5QzFZj2bnzXaMyMpirhxNJV2QdBHdGc3zk797YfGahbB5X3MrUD9nvNJQ
fT54d2gUBfvfeV2xJqkzQh1vabrjM0hXdGO4heURUHFLVNfMRuRXxZrC/nBhNzXD
9pXmKHjqfKrmW/+KPynPUpD5tDfh1QXv7WvYVD+AJgBClQp5aVt10BJiSROUH4Ys
rkKufErj7QzL5NSCN6tVegqzpGTIf9SjGkdUjS49RfFouo8RFtbOqWDcSbkpYFmN
7XNL8kXR2xPdWBiiu2CqiuzF9zdJyDgWcgnyp03RVdH5x8h/y2PUEWEqA1QfYIXt
fdmk2Y7SgD8xyIH4NLq4BN6wvMtc9MlZAlBF16KeCo+vHxp9VZ/3zBVXIjvD+Q8n
ua0WcsaHKGr3jQrOdx2z6seV65gLqRasM1eN1CkRgb2gix5Pas8ujUrB0pK9l0Oq
CEdfaLTVyBz6MvibWLK7mId0p0YyVAU6X6WzCy2bD2yL9M0+QBI8B7YUdd8DFVQT
Z9bNYqhQZj9Hgz3O1cBt5JeS8/EIsIpf6jmLT0vS41e8AblDMiWosNZYCo/ivZ6a
YKdUbPKJkM/go7laselQ26UT50+w/TGZVsypVv75ZadQNBCvIXjlruho7Sn9lvFU
C4OgAc9VS/6m4fT1GWI5IyfRfO6PUuQvFNwVpc0ZVhsUHHtNWcMHyoZEhptUDmBF
kgTNbfMliiIiLEMe5C+013dQ7JmdVROW4c6CRnaKPNtJZAXK2aamLV7TAZ/EyzFr
2U1G1GkeGKLZyTAxuAkjeYl0E0biBz5sKe9N9aze7iO6APt0WEFTgPoxBRijJCcG
vxwcn7OmULWH6IDvV5TgndtigMA28bjuLrRYlbE5R0rSpzsu4i0LI+ewo3m2KP8G
BcDQHIoylPT8iyFh4dwPGflf3C70SdHquTEuezdhyp4qn2WSELRwqrMenihE0yj6
zWEMeXmldwwheByJNjdN/sFIM/zmIgJ7srQfPy66Hj1DoDbz7EKVnOfwh0yLK14c
Jsw5i2p40tAj4TOHjvjVgq22x9DlwxrMzBpfKD8y0RKa0vvw//m8mbDIrbn7B2aK
VYktElhH6hCInT3lJW0T2Pa9hGshiaN8FsLezkbyC6HhNQb3Gw/qbHSZ/4qW2s2r
rKGM4E3h9r2sdopsCq05kOYsj+5LICMFUgu4d0g265p8sT2ApbNRLjti1CzTnsQW
jyvZBL6N9NdlveZoK498+rIdRMlZx/XOMBDW0oyrCzWyspH7TxuXfBZbc15Y503L
hXvdJhHulyJIi7EAlyqQsZLAdvfB2cYCUobJL4DKvX3q7RhE399ajj/qKCqlG3zA
nw6Gz2Ox4rP8vR7hBAdLSQvePPSp4IkMi2DG2Sawi6jyxMeKPOid1phgoZYQBvYf
C/JpE9rYvvLmc/7gY34O93p9yLT0RHGgw8QUY2wCrBplDCBM9m3/rbO/tIe3hc6Y
SOFhNXE522Xn9Wkk8SbmWZ6GaO7FjTu6b23QlLX3lK2Nze7r+9B4ONqanKKxk2qQ
7J52UUq0uUqf7eBhN8qR9jG8kAivhAm+4nCmoZ7FUvzhyGnBdCzEeIFMu/oXRXsK
PKe8zVOSm/a5v+9ZyWwt5FXCRLAVF9PhkueJHv91rTPgCAzv9Xvwy5r4Q7OctTbd
ReJgN6Eyfud67zs6MfunpxM45fP4dlDSB2VDWV9d5KNZaIgzs/GPw7XL6dR0lb0k
a7mdmspKAozR3CGj7a+MYcjkuOjlwrbFr6SkdS1JefMMK3LOX1INwJXwWWnUdySN
2rVCXkz1JD+gX0foVvCxvF+TQBt4K8FnF7glaqrBoz4NUbXW9/Qgl4iCC+Ac+woQ
XTQr/P8FuD0OZbBrPfypFf9k4wqgghiPXOze2WcGT+vbWYvLEz/qij3OWLODflLV
8a/G2oYZN2vbSxiMAN9Ui1iCxsgDn/PuLfoi7CGhOrkBUdren9ZGpAWkcOj0QKrD
3qazhq/+STXXUZ9nIj8eq+xkvhkEpcX9t3S2/oK/5VD0edlrm3IW5JnaO/9SKyDu
lwihXjFczHu/bqT2VxP0FL8UGVlcMCq8wO0e/h7Vl0KED+Kbr88xBP7kWMc162Jl
S0hwxX2+ZDsDx3HSLeb4AxUpRhasT8IvwZf2wnl9l1+yvwvWI8VEAFBLzIAniBwe
JVd4yo2hfC075ZflcEvEif2PkxBjLdkc2LV1+BGOpRwPbwNNI6fGstaIaSoSwGUQ
N/flgdxn6Ygl5jiNwM+mF2Vr0jYmEYFUpXgUhzFjpySn7xLY6wV6tXqRvQYJ3Rgj
r8DIk4Umtniz8sFQJN/sICd+VBqXDir56GfcNdsBkfj88j9qcE32PLCNY+avSYoG
zmobiGWytQbobq7XDcfbB779SLjilhBqFowGJ5WkrJAxExaisHsJpcL+s4fWotFM
8M4jsAC+rO6lC+pWIq8DUKQ6okmrEUe9LdVhFi2Fk7POmA5xxTkhNO5fiyfoHKOU
LxmoXqyEINJ79+FDQkRFdWroZj+gR45+TEEPftn2cHqxCTzMqq1LtLfTsFJu6Pk8
X4OcHtv3qmf+yZ4ecz82cp8kAlmrVe6PMZ5j08MULSMup9h1c98vanEJg2IW3cCo
Gz6vLUCmO5X1cD7h75kuOiD4Ygois7e/Zns0hZJWLVOUGdIM4tvsR0L0Ngu9ngmC
cNx7jrZuAmpKtuWsEo/4sCXnxP0YD8N0vCyVpUH8J5JS4oZcblumK8rntVt3+1hA
rgMUcTkaaemC/H5Zc2r12v7V7AfDzKkBi1Rk4T2hLzVmLl5ymNq0eBkz79NmhKWD
uV6cNZ8ieDI1z465pn4nzWShXDKcMlrryd7+OVTpYn1krhhJfgBlRhYkoUKhsjFE
zveobxgto9fhxl8A6LOBTyx4n465AJ3b5rAut6ZE82LUO8QsZxoOGVY/uy0adcS5
WUvDfVqMN2vholS0fEtNy6d0I3hxkIu7OyXP25sZdauctJ+mMr53YF674kmKo//V
0HXm4EtEMBsBYYzac3D3P2oumrJVL5HXvMeDczjqUyUyIdqyH7U0ckne4WkVy6t9
WeIzQ28C7okdMDnshO+CraautD20foSwT8yExB5Ift/lOyfIHlgPXeVg66w9+lU1
k7usqkCNDJwvvGNSdf4KPumg0qTVa28FScWsmCd3nHjcJr61LdBzLZcdPMIDa5k2
Xpra5HdflszGw1SOe4jdfHapwVx5NOJ1IxxTsD5Ddz6TFg+yxY5KyLghbRNZLnLT
xVL9notlm7ccXgjn10Gacg238/5A1YqnQ+hSU31xM5rWr1lrwayIMh4aJtKhkNmv
cujDF8yqbazzZHtvLTNCq36dD01lXwykvxVI7YgjfUflJpdySlxYoCzN9hdFt/Y7
3tYT5Az65pIXF0XxUaOnMolBxVjyxfISDAHXJxBgs8IXq27NKqEL7N4z4KedUlzP
b5M/BrZMHabecZMbUcaQY6M7sC/4urvhN7AoutpCWRhzFVEYHHAXCbAXEN9kpmWp
2axi3EbJirxrpWBovONGqdq+CNF/nApY9dy7cFS8npVS1PmGvfn6L1/nnCesKIcT
vdVFcLxdxDoNNBQRarMLu5fTvhHnXtgzeZ1v4cTLQmvdIugvzu12mQgzt3CZt3fz
xiU2cYwgnWTgGjn39Cj4PA05QyE3Gc97CU6VYxKgdxfk6ONnPmJ57gkQ0sqmnLIB
k9T4bytnXahoXORIbD9SxQ1j2Pb4TL0teWxBTjnCsXw211PagAhgzlCa5WvZbzSp
5/zQkeI4nMMkWwPmzwh5SCWn/qBXj9LZtgne0lM4S15VcFR/Z5ZL1siLIC/+v6tb
txpJU0VCWUmrHIeMPUKUfNR7FpKdvjYVf8t0zG9UudQDvnabk+Rwyo99Dw3Xwxrg
2GtyJPuCpRFj8dS3CipDF3zklInrTE/iLfSFWPK8SJCX3eI8U7xJNjkCxOxF5mB1
DAPzpGGRn4Hhlc1Vu2NAKidz+EFjVHpCVm65Hg6ErbrbNdgg9wSRMN6A6OYrj7X7
s9+AmCnJlmqHrSKfgZL/56KHNa6zvWHvo1Ko7NSOtS45xuPEjJF5cSdzysJrCUXD
aoRoI9ZuPlzphb2YG5MFh0JuIQHZzfUc3H792Aty1O1wusAJk9Uk2IWPpjc7MINf
WerlVlhmrZ8OY9vJsDDEgNA2JEAP4o+5OdpVKzqLPVDGIZIoP7OYEdL42FW9sd7G
AEDf3s4JwtVXhiWhxqTeQ5hdOoueIkW4yJkn2ZvCIOTRxSurBlyN0gUZf0lnE0Go
RAJiLn0+bxowfQ92HCAeKp4IJuATlrbbeQd7q6T1H0lv+a5ijQZMZzbk2ul8JCGE
842QGvJ6Qe1/SUEooXCi39eDHkWHuTRgJeRckTF9BB2SfQCu7XEsNJpvMc9WTncp
k9eJkrg/JEa1IwydEXhVHwqBLxkWweww9qCgtwjklcFe+q1FmpEGVHmMojVSGo1T
cvWbRD/8A8+pkhaT9kYWaNu3/BGGbiMYqu+SCutJOTVZXNo9n8gql3YRlDp92rNv
AoramxZeuK8BfRNKxoj+TCHUd9yGk7cX8la1bszd82FGMl/ZvxYLMJK3Hi9V9IbT
31T2WG7pgFGyQCkzjbVkQNvRQ74YSQ70YvBnwUx8sLS6POFwawDFOhuymPm+6ub1
swiVhXKZglWM5s41CCr7g+NdvSkvLkv0u40w6PloUpB2KsHQibAzNAXKp5B38Dw2
v57KucGhml4lwUoL1GzzUejUKl3+xAs8lFAS/iVtiV680fCac2nRFTVDH+dj9QsW
SqndSHHOPJHidEJrpJBbBDw1pFkdplsIuk04x8llrlLRUIKMxtfYKAxfL9TgWjXJ
DvD3Ty3Q2ys/ScBrjXavw+D2/TaPSC/6AZC5XjJlU4YnGr2Dtg+gaGI7MKVE/Uze
BP6rI0LELdSbin0rLS2ctmvD1DQaFg/diRRcFXzDCeqvrJBsbQuNWYr2HnTH1QAV
EG04jCt/km3tlxx1dy/SlT/dCtDiSoAkp+iq4iCFcr8yarP++rX1oN0JPjw4HFis
MyxvztCRbFzy80PXfbBK1XfqCYbXNeCTcCMVhF2FEhdVqXuZFD9w1GwZLNy8L8Ql
uj1pYsTbx7O/dhxLrbu0eAqku4KiKo7ClpSB2qvLZOV83LdfJDuhNOLj7C1NeMxJ
LvZlR1qAFOVYuY0JzX/2lQo1PPvBqVKF3wN2ACm5KKdI5s8DZ/S69xQg6xj8PZ2C
nxj1yaWs74A4mDkNtJ+3A/AsbDU0+wU0twXWiQw/YVeQDqzppij4kjV9Gd7LS5He
Zodk/zOOSDDfacLpPrfygkyVG7d0YSSPZkGDqymSwpdw1KHr74DjLbJHNhnlPGd4
H+rBjOKUdQqMdHQ22uTYm4g4CxmhDF1pcv4ou+/IyRnbXir3rzGjIMg8LnPvRe2D
2FyJ3wnL29pAQkypyAlru2qanINdc3GT97WxX8cFyn74d1+/DoKYjDZjmzG7kXcN
tUzvbOYjTz+W35itpKLrnkknw5bX6v2KCK51ZyqonC4N65SbPwr+G7dysyC59iZZ
dpl5WhgxDQCc4RLDGOZuveUR1/1HZwSCbE9XI/4QC3A4bbkOgBgR0VqLpSeBYhZs
yMr/+Uazzftbm6WRBKyt37MC2IaWqeek41XY8pJq8uihky7ZHU7Q2j/I8E+8xoE/
Adb0Ilgl4BfMSXDcGSXiml9cDpMP7O/mESGKrnmexODAZm8P8YyjOCJxit4IQzo2
6ivpXKWYYXudxpWW9EFXEAmsI2ECTXdgit0DaG01mk8cbYmWKWnibs+/8qpO0pEd
FUXztFHzh5wyndCLvnR2DbpYRFCEC6I1xPJau3fmsbRmamSXuoOP0ZnuYEOWRY7S
Mlr5JLbd7iFIy0UophP70qQMHckJdRJTn77+XXmvM7WwcAfMUHtzKn5AGFlXpYR/
ytlG7vGZZzutMfb2fRiihY10MRZ3uuZOJqQBqq8SDNTyYgWSrmt41GQXm0cHjuWa
88uxchgqzDSKPR7Pj0IBRh7yjrTSbaGayvcD5es2Z3rkg8Vw/U+It1e+sIkfLEiW
n5csksKB9E4vxrVNZHwXXhh5lWSY5cvtjICNWFbiYCW9lLnQv1MCPAl3f0J3DJi3
Hgk4GKozVKB+rnaMBVk6Y1OSQ6UeSqZl499av8nZ5wDwROvl4h7Vp5aQhPI098bM
xqW18IgSG6wp4zH9sJciGu19I1BCmgel6Coe4WNkiyrP4xhsMq26mNdP4Vj9bJrc
JUAo2zm4UjFAzt1Z4hENavGlxTxPm6Fi5Pu5VWtZUM/w/Nau2KTgLN8HWoDqu+qs
IcrY7yT48lcwi6QhL77pW/Rr5ToGe3A0tvy4f/5pYen9nu0kFbD/Y5goAvvINIC7
Uld/9U179kuqgGubg/MSh7RETi0S+y5X70X0L/PZPUn5rFWqyFPGdsBMuOf0LOLC
3hemp6L8D95og1O94rjdlpdboBjmhXUegbHzfW+rXj7FN7uS//ak3YNoWRco7TWg
cbgA1ufGTWWsp6FkQ8ldtNHWuXhKLsFcBGtQn+Mcc3laKgkj6X23u8WqWVoizwnM
P+J4aTD5e2fpS+10qaqN8civ6xZGmDdTJo6yzEjxFFPPfcOlnpbvfU9ObI08OEpb
rpHCBApo9NdERDXRLJ0fa2ptsLabKKwc7+PFukyKv9kMO4Q/P/brIiYH/YepwIOY
X/3ZvsLqomJCAS4hKM2gKo3FnU2eAsW1ThF9Z3+rDEUDL9+2O9ZX8WXY0ZAoqnL7
IttAajAt0nKseNDYs5DJQ5rKT8R1B/qZYVNDTXL+iMc8o4K8cou6Di13X4MBKtQh
UfYFTn0tPYG4EM3SACeve1iW48sVXOTpiL2pgQpyJ5yswg8AdsQg1HrxG7D/K0qm
aQtjGfNYoGFPGn34UAToj9cQxiUxIzNg1XnwHom/laYV6X1n4ySU8oeT2jLcPrnW
9msn3L5TONDGKPeLcJfdLqKUhSscoVuMHc/gAbEl8A0HU+Gn9b9pKCjYecNgd9lS
6tfUi+mQpNVxP7BSq80mqMyIhIz2aZFbS1JOWmemB4+xua3TzytpVqzfTlu2uSK/
KIPGHvC7L9+IW3UxlCNaXVmrP5ZhcQSE9KyQDCPI2jPpxzbx1r/kcstuRGDLVEDJ
121291i02Zj1UFo9Irz6B8aZjggQUdNH+WBcBgL8JJ2sQdUCcFMXuNBeVUbofVA5
SEcPlSzDWAsCGwZGI3sa/EM9OSdj3BARfAUe/lG+fM78IEdlt/HGTyjI+TF0ldw0
65hj2qCC9yfjvhB9pRL82M+uZdClE1qqsVDaxihCNNewyk40R07YDe9ATwFskulq
37RL4p61cPxC55/apVqcXIzOOwMmuLzcHxOYN8zub0bt/piA8Fa/GGk9cwYLdn+Q
LoycVUBB9kvdC6g0T8j7+ZHfxoGPPuKxx5hzaBiIxlT8FBdMazyq90+x4udwhPDJ
Jxsv+5YjgvqZcVsBUKkvVGteq9TD1Vv1FV74L850kELIRgk7BwolKHnK5sNZ/gWc
TNr3tpReP7zMhvFCwgthLTjoDmAnp7IfE0y05nKwKrRPXr/F4t+z3LYgcUqrVM1i
77mFFGIdnj8Sh/vxA6o3CYDDKD1Vonh5HqE2B29e31Og+HdTzLAF0vEo8LAMrBfD
9zVecHo6moj1RvUYSv7K1zW4pQlkfL4CHgpOsmdFUbpG8Cd14H7rNGQronep3uM3
vjlu0UGByTVrv48C9u19mKKtubmLPBrUohVSZ184KGDnof0kfFuFx2eKrASV5zu2
9aCygmm8si/GFIJNrrnPwTpJGsiQBGLLjozbC74Wegf5HTxE7UHSlWphZa1l49ze
JK8MKl+ZVuCWmah/mRtLpcaUqTQfVK8cDHbtScbrczvZKtccrOGAAz9yshGFxTXj
o8U4oLwDZvUAW7O//aXFFu1h0J5l++vq5kl3dxxRRTrJqVaZojXRABlQOku/E55O
+H55Ghb7otN34o6ViTy2LFkHtIsd8Q2auOFkHKcvY5TzJoHWWdv2uuyiyLThOiNI
ikGGGN+k0kDu7ARuNmdiZNv5IvqEjwaaZoAgiVhMFRPUEmjIFKS5zlxoORNdAKT4
B8oCQg+QY55tgokPKWbXtw+slOJz7Uz1zEwyITsfqI6UhkBmX33vGrYtf0hCnlzp
88DPadQVAeyHmVAIfYT2mK4kU8F2Utw42c56fmrq9VqDaM7asu6u+wkQRPrd9A2e
Lzw9WcKGolZT/fMwetsouqjTORIQN4oTqtFYwG8DKa4v2lExH0eeKmnu1wndOXYS
BGswKHYRrU3GA2tvTMplD80ZKb2N4/Ry2Pn2pe6r18/tCFJuyuxcMrfofNB1XeNx
AtTAYdBVOrOSRN2tcuukVuJMYiSZkR3cqaUGgglPTyIy7yrZPJhCZVyuQBVwb0tn
ROp+4Y2cqrud3dYTCgovho6l7Fk9so7paNxZ9jV1ZUe92KT/rvHVPQz5B101ttk8
REk+xINUjeNfo8ithsGVCnadoNXFEU9c5h2FSTXaODQDWEMrDNT3ebWTv6ZOSjJx
sQMheozCXyN/QhJ3eqhI9KjFQ8UiurCGUFodNy8yfe9SiczfjX0n9vz/HkNRIz1e
Pq+XZSkwIhv0c12V7mcxTMFMjaZQ2t05FpgGbO7WpfAsmmKlqdHx6y+3Y2O5le6B
KazBsg6BBPQ5PLWeh2IlonQ0dhbjEi2xPrshO9RRvjn7fVcJSs3wTlvN92PvHDJH
DfxPqjwMVvUtUuQXb4KznfkCBRo5Fjk6GccuBP/gGryEuS0sMBRQ4gu6HP8VqpA9
Dn1L+e8yWfrdlEHGoV8uYlpqX+AIajNXlcyJrR6M4ilOUyHBf9vl1X/9YKoOqNDW
WUgRxSKX4Wi/6dTGyu5CNRPqtzBQXF1dPPfJz+2XUh4e3wBU9wu3FbDBmK+IrXUK
dDCDfwykWQOoRQ2jyj69N9WrbU2o4A9huYTb/ezLMr2zKhi7wokXkgOgZ3FtchnE
PjDpWo281V09eW0HLhGnV5TFNhJZijoNLR0+LRCeqeWI7ltNUUyyeWebblbh0zi5
V1SHjp12jRP0HsMEk3bt1uG1SfoULhhNXb4VqMCCsImDKSSsPjgsdYs7rmVZ08pr
Px7+qxPdh66M2wTi5ddr/kkLOb3QNzO9oi25evZjRYAIt0MqqUSHRtRX8w4m/aeM
5PGL9AO3gW0Jpevvh/L0N1gBA3YuhLapEAB5tUqbX0hQNihCn6G7BMZ/st5t7b5Q
pxKOwUqTGFIMvqdEP8Sa+ZnzvdxPTH/GVmpcPfOsLBP3Rc5v84aFSVAZYpOik49i
BUyIIruovqgLiG1vHFAoNnintP28QVR1I/H3ZlGE2k9UKOq4YyYmO+ZCPoVDRj3Y
zjw8UKjjr2BimTr4rQk+SginsmC3ZGWKL8pGGhFqCBlS9m2dYuDsTY3SohejgnDu
S7G2jXwx2pSkwUrPjYHSWFhiHKWkugr1a9qPF6yXPsUEMKpwLftqAbCrSkeFeLjo
cHxnncZVDWSyCwe8iEv/JW+hWGyqgLL1hIXYq0LXo1OFvc2JJW34jPkQf8e+QJ10
YhldgNotc1bA96xTZjvQPfmhSjJg744ji9jpZ95uyxO/H2kdga+UrOL8IRnZ/WpD
bSlx17zgul6n1yqU8PpPeTiec5fpy+T+mWOQ5x7slTz8ReajXruNZWSx51Hx4ouq
emaoLRVfRDpy7ayBkYwxaMeWkKscC0aCAOtyAuF63u1uR3XTKoaR3TxgDSqHpKTg
b7P3AUR1rhpG6xLRpPKZ0FHlDIBcnPIWoLLSw7a+HtA9H5xxbCZoTYqQD7+YMhSf
ZJBaNcR/4WFLBSZACTjEeloKLkAiUKe5VMBdYH3/Z/nFeRVxNv0gG0PcNuBWk7+W
yrfQP/66FXI19d6FznGdrEA20dUaFabLg+Lt3GQlaIvcp6220XYQJVcMS86z1m0Q
ZZ43gEBf1KPz2cxWYIpxhtaBa2bNbu2XzqyB/Iy+v0lyB33dUyp+aM4B+NGiynz7
ZsjZ69mw5Qbzej7ul2o8c0IiQLNt8f/X1mngzCC4DS17KhJ00Sf4fL8Ko3Ht8bgd
Z/hBhZ3IgAtnbkstv0BRgpTWV9a9d+ClIfpAQW/QlvTDlkql5NCus55Dg8EkxDEB
+GeTrjW/8MCwV4csRP5myiJ5iOcYcB0EIejYoOm4gGEqvQ8tC3A5SAMPg4WD3VhC
kHk2L9Q+zrW/g7u2N1Fu7lpigb3TNUOOeHvTBuFiq5OyhC7glbCN4YizQWZsa2Gu
d32Y4nZDtCQGSb+sPi+iQBWkmBwASwVuHtKXi13e3CLFELpmsk0GKAzEJ2khPxeS
Smi+PNuZd4yaMWXFfKwvQV86V5fJUp6hXkK7SU1i5RrB3XW+ft/fa+Q00pnq4s2I
Zfsc9S0wLD3QMAUbuE+6DwZuKC4Go1kZmWlGJL8ulb07vr6Bb6u4bjad+sdSVItL
bpebhcHAB/jYT7la2uPhyxOm4qmwhG0aBXHryBymoFnLsXa+Gwy4XmDyaxb8Jhki
0ABvpT/NvInbff2s+jmyKIHLbiURsWB8p8GCYr6C+xWJnmKI7Gfusf3q5/SOtLZ8
fGagr0kI52I0F5tX6QtYCe21k5iYXHRVi8HTpIhef0oF+bot/Y88WDCoxzlFt62u
lLEukTCTMfMaXHJA85BXL8N9CpPZjGK8JRzxRdDLW0HsShkjvpwp7AkCkF6M1Z+5
oq8bqOh95qgnR1mPXYZWCBF45Gy8M9fb6HJvc0WRU8QNUNmtYwo3+rt9bKhO2lQG
c0V3rpYC8Dn7tSYUCTawC+tJco5C3TZn9MKb7suAs4r40yzJV0rgxUSIGRTG4Jlk
uWyEpT3CMAuzBPbVaA3nYVsc9N9KJXTOwUvkz7nDZNVJNC5fYOMD/Up/gTZgUR+/
0yX9ozELjP/TXRC0DaDL13zR6Sh9PBCOurrAz65e/q83VXk4TOyWBKDMEhFCOKea
nD6tMeoDOqjJLAQu6Di8ogosmGz5KEJOp4DuAsgLFkhPnX9J36cFAIvDicl6QV6i
+tsdm9IzV0AL/2grokkfNUjOcMaXYKF6bBJw6Y9cdb1J3zv0TTD4LBdx3dpPRpvr
qr1tligLhH/TePmSOooOc7k2eJrSC8F9lkJGtgrWirY9FMmN/gxdNbN2Y3EUtXgO
Kqga9GYK9OugYSmjPb72pLBeR6i1hlAgrF3sn3AoXQuoKygn0ageAMieTufdiEoq
DkAhtdiTz0Q4+anGxIRxmDIRrJYX1KTNnHrAgRmmxq8NRYU/XgGm7rgSAS7q/vtj
LMlBK6iN7uzHLs9BjfExVCq59N5+dsep6XVXJZ9Pr7p/DO/yb/ikBRfGkS1LtjU8
xRJzZMNcuayICWF50WV3de9oiNJI1nCdulTUrpD+rmLSiLlagD1oNvXjHMQXVUfo
SFY4+aJBlqJmBJmMKUbGXnLcSm/valgE3XWEbvIv+bv/4p6pXCP/UftZheWvvRzr
H4+UAkDoo9CzvZ40Ndbt/BJNbeOzALa/cLGrEGvqS7EQ4MtCY+tBaJ/cIxr/hGMd
kNhyk5xElg/5+u23TXjEPrW9DR7+dbo27zn1IItKi/0AgSznheXKBNc1NTAHeRep
uD+YLdXZKfwTDDnDUEiPE/UdcaCw6znNyRaB7fmgUPtxhmNSLvBPACLJcO7nQ/2i
FJqdx5wAVuPRcqSElh51oh3giEJcfBhD2O0KvsnNd0qGuqpf9M+5jVXBZXkuDuUj
KOvQJigMzZqUimBKyxJRGyoggcTe/pkY2JJvJAgcL1xeC4XRtMfIxTiiLuR9XGza
nmKtA/rhO3h2OlOmTOYCtBzGHW599h35kxv9lUuSeaVH/+h3IvveEwndZovT+eeP
xMxL4USxqF0TzO5rWWVoVL4qPxSyw7pg93PxYmw/jEVlUF056eqzigxaVm44L1BV
YD7pfJ5O7IrwCqFKoT5OXpJET9wF8/CqzDyNDn7mCbwJNPfbip3XI+xnQFMK0jro
6L/JOI/jmtiiV//BIbr3U09Qr9ti++P9ZWeBaYusCWx+Nq3lrds9nfK84CrfL3Vj
ZbH5KVaHLQl63MeCnH624DXNBrop3J37FIxrazNTD2oUBlj6St2Vtdjm7jx4uhrK
YAIXzUl7uOCAhr3mzdbUYHoKnh57Jn/Z5MrdVsrmXedyCZJfLHcfpsBgvcCjHwPe
7On0xh13pIBXEYG2dPfbHlNp6BYeDe0GZe/lGf9giM1fEOVLfgB0q8LscXxkD0I2
45jbJEQGzeBT7RF5NzwnYXwGibT/qUG4LMvvWKiXFF2Gq1G0G9/XFvkqbEuyy5bp
+hv10qgmagbnBNqMim355vMGK46m5eIRiysi3mKzl/Srkzxk3+/coOIgRPExCX3D
1hwIb5qS1romzwIRHCRWp6BeFB75iNYQjPuJJNJ1dNIbKDv0GqYqT0KclZvuBlUo
Urb175ppTx+Ur8Bprv6uY+eKiM4H8+J4rOmLiaFo+dWtD043lY7V0OZMfHW92EkK
aQtMvX7JNswDbAql8x9zUVnq4FtjZxgtWECUelU+DXI2PK+NP0XRrp88tX7+/ICl
DSqBQzE1Cxq87/Xx8DFa1dj9Sf3WBOEVHQDi2YlZDdeWJX5AjU0aoL/NU+y3+BRx
wazbwS/O16Amsi3EgMF1QELqxihtPzZoad0r9PG70BxGnGiYpXrwOo2JaGHizWHM
99exO2JGPkP92YLpM6ihxv9HlnO1VM9c4KqqAlTVFTpaXMzmc4bfQpTiie/e9Z9v
QwWkEUJJw2AqbnsOqkRKkVXXpZsNFhr3v/tK6LKJY4P57TVc8Y049OA3a2TSxsFx
rKVFSEtdhluswx3vQ+IZ2ZQlm1BSIg33gSyMQv8VwAzH/dO7MFDgy7To/YypQADM
8De9YZOAzzYu8ADKwy1tiibjXtBYOTPpWVCTtzuWx94VKnh3W66yIQdhJJnHKDxZ
mANwGgz6u+4Ecg+1bvqJLjwUuUbz24Tb+l43NGtmgCGRfcWEG7LEiioZyOF8FXsV
Z645rWZxFIkjOhlq7yANjjl/T8FFrNDZgHaECP5gzm4wAKaD8qy5ju9d57WhziHs
ezWt0D6bNWf0iSUgaE1Zo6cXTEulkEdTlpfEarWH+dI0KYnqoI3sH2t/NNyZKxO+
qvGbipJmqefwwEv4CxX5cfNA1p26SzH62Y4ampzk4V6i2Nhalp0ocZq0iTcGWG2k
z1u7oFPqn/KcT6KeU+kR/IbGqgflXloMLofFL6daR05GVfD3w6CUOXYEMAnRjNxG
3/AR41K3UPBj2XY/UdcWaaVH2kb/mJh7JVRiER4D3fTNwEVOoodN67+n51iJxbwa
x/4oA9s/mCUso5nn/wrTujH/ZpWyyFHOhdNCTP97BCmSz7MNvIMLhupIm0UrGx6z
lwbFRMgKO82SPTpwo4OA1r+5wChjawAL600O65J0jzys1VVS4XwFfsA8L0hSxW0Z
Kc+yyRLYl8qdiJPvdv9L2wlL6WG/kEdzkPv32ydISBuAduJq8SyOUl1iZ1neY/s8
7OsFcwb3OwXSRnB/bDisW3UTOW8Ft+yC2ZZBRwTzes/mRYrMM/F/kclKxJGaTOQf
RuU8abj9VbRGnCevigOrAnCdklSOa+SgC2GqZStb/eUhWH272O4vfgQLVOEglKrE
ldSbaBwlsHD+wygAB3uwh4b1ZeW9v+Oyjta/71iwvjvekvYjczFhv1GV3dyT+2c8
OTQ78WjT9mSh4Y5/f8hux/YC9J7KGtMIJHotOnyXrG/Z/AkvcXDtpF909/LaczH3
4aJ/T+Jw9Z1wdAA+kpOoYSMROnxByJRkLFM5uPbeyYMk+OBm31xCC82aG6Z5f9UC
bCuG2e0N2S/GFQwZrhz8H79eONkjfEg2UPh2u/oRh3jkveQaFr8jaJp8YuCcIgaO
lyOTag22W3N7fB6Mz3WVyyLAEvokM5pjMOBG698GaTRLYJhN+swYpbkApS5w9Juf
IVJ4czvTgJN4tQ6kpzMh0Of2XnbRluzPf2rD6/9Mq4oL7bjcoVk30HuS21C9CAr2
6pFt4fkbtO4fb0zo7/TJkBTc646DE2QkquWpQNIoXpDzxJrhyWZmfEFXqAngfhfQ
1Nnj6lCJIYFBPrZdaZ2EThDf23kqw6VQblohZy23woyEoaXLzEs+bgXnnzFhFfCx
sMqg8YnIf/TApwM5knvY9FuuVhj9gL1tyb2bp+ZiBgmYs3QXrhfduWlwzbz/UCIU
GXPNjqsy9js3ylKskymgYAUzBUd1XBslW1h2Be2Dbq8bJGf4wTV8ZcrmKc+HKBF9
AsWXr5NQqD9DEKfm9OzSTbakkA8K8CkbQ/uJhEt8/wsHJxRW2g7K4xZkuZobvdHt
5+QEWZY7x1pLO78RZBMwBoXZHaeMi+GIN+xXWMi59QBPDZQGDxDl9iF4Q6EIBRhp
W4l+Ojrm/JwGyZABmjJos4OF3aT+UlJXKYipIfy1yNfbGlN8woeQYTTLz7dnfNbR
xaDALL2e8+wipWHSyvUPFslLXwiq4YL/YAMQ3xFhbgtQsEqqptIK8OmPRwQ8a98C
ZLKOWgqjGZWPfhXdlisU0EIKyK/zaqTenkrqSax5ZNqX+/MkDGO8Md8qUy0yCBSj
hY9XidALvzTLaTt90k+eWuY0OP8tLTkQaNRMxBrC2gqdfzpx17hfq0fAgBUc/SeF
l8d1XsDrhB8M5j7C4a3/hJuFROHxj6qfRX6pGEZw9qsKkoAgMKdQma7tzL4fAsSg
i4A4JwaDJjQyv41K0xnp2XRBxd2yD9VTlkwnWJcEp1KpesNjoUUr8j5kltc0o26d
7hXtXcl8Kr3QZj5EHSJJLjI8ciHsB4ajjjF775GcRDIzMFkVYy7a9Vhtbx5uDIJ1
FyhPNsQ9y2fm61sFYcRwtjVK/xYBD0Ilxns8nP8f1iNTnkKLwpJSO4bM/IXq+JJ9
DXO1/6krV6WhOJ0NnNvMJCpyaTHVz88bMmWNdY7Oia5RmFLlkjF+1urrH1rxvB9S
gkwDDSVaj57xybZO2J9PYo4Xd7LtFPLWN7f2dMWDJUKXQ7w3RHbNgwuyHOQ2v7YE
LSKBWGTDUQ3uaVcV6W5IHxU1TZeh2tkm+mBu20X9rouVxydWhUC7HTmQaaLnBHME
0aV66qr5soe5l5SCpgnKq5V0zH0ix+wbC5y326R+fD9792TRzduetj3kTEPr9+dv
POPUiAL0SEA7cyFDrz6AQ53GA9r+UryTllcWIFlXYnZYBbsDg5lbrJ0Wxj/H7frc
2+n0R057oPxXlNxdrCOVcPVuYh9DHrI/+NSNYrxqrh3K/0yo8+JmIq7GyImm+eMc
tQ/9O67I7VZlHrwGFYAQmUBQb8J82wRxGlMEZ75+ilCl8L0XIiwILK3sAyVJF9wV
VrA8Mi//ouH3icg02NGhIXo55K+2uBs+bSD9TPbS4ldPlqMs04LyWQFd6X2izaJv
eZTZYSxMMioFVLxp81Ji0Eh/j6IWQ+etZmSwdfn7rDmgzxlukzH7cbnrxfM7DmJf
ZZosDxX4xDJbB2CY7Q3619olUeaqX/etYYtjve4jRtbRh9TPTqyADFAmY19PNmae
I6Ez0Mxlr+hisd8Y3HcewNmATKknuhnYUh0tHWcfTZsQNA5LWVsoBxr8kS+d71rQ
SupXrAE4ar15+0rllRcZ1S7bwaBb13J7j+fbknNUIxXEk9v/JsulJZaY6MEl85pt
uEN6pSW1bGxTCrlyVuzAalvqQh+mFwlC4urOIWY5126AVFaX12353ozmwzTF4ZxC
cT+zJhq4745Ffp5b698uZGrImaMxgtdok3UpBTKPuR23u+H4AlT+fBMQTUikchb1
3ba7K5WPudXzbPs9xmnEjWwWm9z2wmkWtYvYlF/YZUE6J5Z131Xt5aDdBjBaKtXU
N67tqOwK6koME/FPIZpHvwtb0b9v2P+IcuFa8Pz0h6P5wmIgB0EniDYxC74aXNsH
lV9OqYueFcooEdaPYXBeKWEjpspFIllkm8r0HIb1rJpWP6xN80qBRM0b/+vZAPot
ecdOQijtRY8D9RPMdzVgspRyJiCiA35AclnU1oUWWdvHlNywT/qP8y7Es5E7cHbT
QdNndsGYP+qnj4JT91kgtSZQDqj0fIG4Q7DsaoGshkcxVgUm1TOhe862QMQrRBGN
zLNC3Qrbn237eK8P+LcBq0PBUU6J8D7nNbLsMRA62GYSxiV/x7Dtu5vSDtYGcqet
Zo+e6uBYUhhtMldsRIW1HNwe/OSZcNIOJJ70lxevJ1xm2WCK9UbemSzxXPYm4n1s
8FGEujDuzyDzbyrq5D71HWmQg8vpztdzzTNnhRMcZFAEU84H/saCKZT6oR4oMyzL
y4B2Pp03GcN570m8U/DtYwgTQPmJKsf3RmX7z3/QHjFZ5FIeFfwpgvzf8eis1LxD
w0K41GFEvAoKagm2TPMV1jyz/6qcc2yPF3jHM136XQaJCoJ3FrrlE0wjWrl1qpai
0zSFuz4JHbRElQGgpVngs0KQUOS7/pD6SYghO5OC2dEKacxx6btguEenqrr3ZfTN
HiEDKryNFOB5/CZ39Lkaphh+SjM2+17BXw3ceXhepSgnentxzpCL1RiVIun3M1Lb
QauFJ+AT1hsznN+OKgp4137hxOg2OcJ+n8tt8bxFIfm49/1r64uZ3bSDSxFamYzq
LQcss17Utp3kU5Jdn1Y0+JWsqwAFtolC+LDxCuFI9+X9cpSJ+IplXmCa+Ov0F4fL
NmxD1n/wKmyLAzR0kk5O3cK711ly6jZ2D+SK7iFap1UwPSxAnzBn5jwIF8s45a5O
GbTnOpS/F3T5H1nTjnrLvEXk7fQquzhUn0wNp76i+fJ9mFE+p9exg/bCINpw9caT
TDpT5ZrhnidIb8VoTec0KTG8PtfjengAZRdsI3EL0zE2YZDzIhtgea5Y8eYbrcCf
TNG2aII23o4Y9H5h8Kf8dNvRFuRUuSrykM0lqrlrLzuoOeJZp16AeSAR+zVVxjJI
6EZ+6MFoE1ESxCQmxAF6+YS/WU01N6ycKl9vwRmPEUR1fKcwWEBN0pkR3ARHiGve
s751abqBwz41/cubTbRSh4c2yUrG9Qyqp0HZFSAsQvf1AIXA1yRPvdRAoXZ+at+G
EBgn45xoOovAyHsLptPb1IzpxpU7SfOperP1bt/xc0v8NWk2o0meF3XJporT2xA6
vv+IOvbDd5LUSWdB2l5tP2zvNXXYtBUVzMP0YFumEBvPbb2H3H2I06oR8s8gHJD4
HdP2AuO8yd/sCi/muYTJW6v58dZlb9S/a+ADFNVnOvLpjeoylm5aj7PsLGA9gyj8
lZ96VuMNVXv1DndSD8ZUl2oYNQE7rfeTCSyeDm5/vBomJgLFXALj+DufeE/367mG
tCMcsGxE50oCvSqAETx5O4/VqONK7xPxsXcepacUSQiabXBwKOhpWLzuyiMkCV6f
AdabRNCOLGeMlNRc6NGx16tCsq811vBnAB0i7xK06x/DSpuvCH4F08eO8rVAQIdl
dtElI8Z4BmXdRv5KFfiJckj0m9cTPcaZrEKKRf6PcGV46vTbm28/RnwCby7Zhadh
lRIk6bshh5oqndbC6eimaMwyY5xCEiPRSS0ZV/B1/bGxJeKshSQ53Wk7DSvW0uiX
a1PYqTUVYeSVZoV+LbzZ3rxeCBLqRQPcK4C1W3BE+gHcyzzCUcR4tfP9j0I49wQj
hIzmoRT1Dzr3tnNbYyH7m/ZcjpKaoKXHMt0OvkBtOdca+LJajysaFv8fvyIJFCCE
5o2c1KqAF8F1yYUwHXhIIpb3jc25uLSyRAWSnA+m8Ipq1pkwISg0/F/PnhmQc4xe
p5whjMdkmoxYLmzSKcE6qhqOT3qDrQejXK1M201sjtbVJUmRGaqT6miHk5Td7N2A
DlDbqROQodkKHUvAEzCjVhQR/MSQLP8/309KgZU/foBq3ufjhEdE7JlRIvUnv955
cs6lfDMjRZdWXj7GUcO9UyYw72b87e1420la6Bnka217FcafLTAOGfaKBmYssf3D
N2xf7SreEbRl4fMxemi8mVvS44axOro7TyrzWakGN8RSH5Sw8UOg+X8Wi1cKMLjx
MhA0lsn/pBP0BXnjT8ESPfrCqEQzIh5ASI047FIJQl5v2RI/9A7Jx4GfiOoF50+P
VKbmn99XPzUe9FMDeiTUR8L97upeYYXNJ9aXq5/YbB7xfljS/6vKyXdJhMZ6tKKF
UiawlDeuyQ57e7d1MzmUX69V0ASWWZQhDd1QqvHZ1s1mAvct7ds8R1f7t8tIjfGK
OKJ++F130y+OelxaG7SeBltbkqwqPAD1bPXi9dEoXT4reawbN3CXI4wIhPH8P13+
NrgNYLYOfvJyBn8MQTbDlRC9HbC1mtO6cbwzZoHWfyrsxSqwvbczJ8DqCwQOjiuU
UFY2auHOUSsj1bdXpvIrmfcXqGPTltkEAZia5OuDtU6iklRauO6EN/nHCD65Ff+R
SqdPpdoAQgHeCak2lKsB5o7VJ2XWk3LBbPInvceL+eaxdvCv4QDrp7U9hIIascL1
gf6704WTNC4QgqTqQogr0lrfC5W8pgHp6JQQxNdQ1Mr4WbDHqw0qMm/KXFOxnjwd
68/hmzcRnmT+8gft6Rg4+B8MiOz2n9/YNEBVE3DGDgqJeDmdoNuoRxqhlGYfvSyk
19tyR06HGLDK1mQt87edFGdW0XJeajwFuCr7yMTeIOvS5pFuW72VJc+KtNjO8qDm
YXMZ4AsRmHXYxMXsIJqKHF/E3uppJRegwq/igy8PEt9QvhSsJ9iRCYfhTj4FluKy
NjGsawaG6F5y7SCuZXwzhLlwKrTdHLou+i8HsJbB9y9pePHMHvqlEW0M5EYiGwjr
iT7MIDFgygNxTiGQCVUH9blxEwcChJY2SrnKP2K2bElBKp4B5ZhSBctrbpqEZ3Cg
g5UZDS5KDQ19g0YCr99YA5hWCSo7HqZ53wN5/jHCUZtUabjrKWI13ZULRulaQRPB
qm4Jx9Dn4vNSFMNcJEfyQGsWLD9Q0EU9JHQ3ByWwQOIMAvQI4rMzNHrpbHQjM4ZM
0QVyez2OB5WAaeP6ZOD8hSovN8koLMf0DcNVpLD3FKpI4b9qJgB/ivT0z5m3LP7C
jMC/Pi3OXQYdjse92SJ3Fty9frmmxuikWDUEj3nVE4RxPc5zMQ1tGqxuvI7iIWzM
F534+BC2IvEKxH+ZAqfqlIuw99MMWl8hmSPkgKm5Qho0/Kk6L9X9ZZGaORzs4HY6
o59dvp5XEVqf1dlGmc6iKzOh2FUQH/3LEiitUUp6B2U05Rf3pPYUQRuWC3ejKGT2
D3GUnb1N3CCb2puNJXT95tRlDYtXDMVcMlF4BCEZu2mJU7P8EbdWuqbcPaP4hGDL
/xSWlFd/Ii0olvp9+LMoXMbCAB4OKr6NXumdHLLBs+MFIjQsjiGDlt/sQ1yVyR5I
TWGlX/KjAKYeNUT49j18OR5MZdI1NzL4F7/h3mlCYFqZz9qw6KsGpYDZwrStpeLz
fIaHUExsROHEDYb0EH/5qtjwDZEMu6omCduHERJmt+SfqdpyCP7wmBrIJTKEgD35
n7UrF3qYjIyBAu51dXmIAc54vfACkPUM05I6buu8cLKdQLWScXaW/5uTMM3UpTYp
8YuEAMKpuppcdf2wTB6hO4zmio/QnJKD+CsuQJa6Lz5jOeu/ei/UffS2cHkBZbwo
WV4DaiJSlOzeBMrjXkJVNkS/2bp0CQgUYHqK9rbUtYZwexJvMiIgH5EeS3/CqTBl
vjWoAgqd54C/RiaeoBP+xNPcR8ziINjxUYTAvck3vSbFJSyIBT6sy46oROTl6vGV
0UUUMc9YVUk7GfwrfzRn/trvg+ZNDei/zz+dEjIqFmh21jdvR7bqLMWzKWDfoZ3h
sFIXP2rnC40prH3Yqn62YNdY6dzAb4egnSC7sAqXaeNAVMHJV8djiK4XeX0Ct9BV
FISXmZByCb3Uls48Vfb2GD08KNGcCgHFpq/J53qWZVEAoPW3VcxD9U5EY7I0blR5
F2F8n3U0i2av0ANe+rH/R2CmXxjicCUa4bQAoNW+uOdwGXsc9NoPo2IzpUsY7KlH
rDtEiXFFxjM58yHPr9C08h7S7/rD9y3R5PfaiNZ6SpsBZyajBlxbViYgrIXyxjhT
LufIlGyGppg0uAXeFXAssgyHxVdD0JBkXgwcENAS+lAyF9DQcVDYzeLBOV7w1Qo1
JFbjZY+dtsBNI/QGmRRkHuHecXtNfB0VFBnutWFUb9ihOEEOHNbcph5Gv4QQRSNd
JkEcmtEAc2+DfQU0kE5gAkMx71MdBJRIdNXEflQQngT6bGPigBTWlCowcds5QguV
DJqLpDq6ulxlqkRzvV5tjPcSW7dU8+HbHeZOo3GsjPs9jcVIGdNTiFY8XzP7LesS
BSy7W70ixhtr4cQ2JpFYwC8oI7FLY3ZXyGvSahC0AbHudwOMHU6J9dgfSLuM4Etl
wgmoIhVq+2JtQ3uP9myDj3GVUXGFG9Csk8FyvD4iUvsoqOd/6mCvTqleRMT4bNya
APcQe2E7cH8PofGsqorauxPONXVCqsAa/tRVAnaHCaVYURahqAMUikLtw62dhFfU
+mECUFX9cD2BaAR6kFgeA0L4YzgaPqxwMHUWTQk+wvH049aI7zQKt7ggSDm+3nP1
h5TjLOg8Pl2XpXQTqx5qyVEFvx6Ij6Q7KtlmeHGEyigSaODgcYoZhWgNx+sFW6qN
WEftqiulrbNSEWnZD98DyN0ZBeBVEwv5QJ+sootgUyqJmuOP7Gz+jb1+3EyBL8MV
2KweR5uSvgsijxT3QYoLnOGf7GTwMpazJjIN9uGLDiv88CkID0zK7f7bREuR2xnU
7Cj3v5/TOCiSd6mh7UnfeYX90dBz/hZGY1WIoI/kW3XZVXhPUO4WySxnEcV3A6EO
cRULpxH9vClAmQUI+Zre4j9eeDIXlXNy9x/ko+PlAPEdIGXPFUdLvgDDjKUwBrP5
4qNRvB+HRNB4oEObLKabgOLpYkhCMRj8xf1V44i2dbvCTOeH6X89xQa8CJtkv5jE
82sVBbBVb0nyAaUR5emKbZUE0VNbhSi5fBKnqYO/Ohy7iEzA9KE05lvZIBRbOQbI
kbgB3H9KnoTVmqTr9V4eoadmNSQvkHIJ7BkDRGeYhxW+Zofg4hDKrTCP7zxau+iA
uUqNVpYj+am0TGN1MMK4IbAEQ03OuXlLaqI0vlv3BUBMP0EeJDdkGbaSDVHB4aLV
FqnYy8yzYtINwLwQiGWWFk6JeDx/6yCEch9dZCDGSw9tvkwbYzyDYHAsoMu3TPZD
zeKucrm/NkZFTg0y08SK4xpwDB+uD1h798RUTcAFqVmGPZVvSKMIfdyPZ1xdcWtg
XOJ7heT84/FmYCtajI2e9e3huTKBpFzRELUn/sefwbXMOS+DVIpovOVOdJm2cqvc
kYul5qc/yxfENSRfxOE6JRVHK5oNvI/OCjg3quLkqyK+fQYEU9oJO8oS13HEt1se
KIZO2IF44fyVXuomlZgQFRnTk/sIpLlBQCHbfzC6K0Tb9oP8B9o7bq9dP/bUMWv9
XGpOo4+c9yWmhPbR722rc9K89d/RE9w/2b7UJjOVmUaofu4aR+TsoVpPoYcowTJn
8DhVIBaGpXIQn3Ep54FgCb8ir8JdczlQWL1G3rwNwVI8nlYaDyU0cR+Gj8mHXRPg
afDmzrVoYMAooMVX2G04Qn539HEHh+gODOQO6FDnErofDSG5aT/fP51YlOBwLy1c
iJ7Kiv04NiIl5iEmvL7+aHOHwyt7eIf/VXx/zn6l9EjfXwzePbJm55Xz8xs7gL23
Rgfy2YI2+IVlkzWAsu0BL748BwaNf3aIZOzl004djTYozv24lDntfEoAOpbmmaKW
SiHX7yw0qySP2fcS3GO0bu25YvlZhStjid7gX5idSigRrTXAjfAzUL3FlAc+UlPK
5mCrMLy516/0SbFMsN7YBzgcKWtJBEpgs8GYbqO+AFhPBkrBmYwoWIwE9PFylpoM
qLl2KRyvJzVMo1BHxNnAkhFqHGHmuVtCmuubraK1mhnmRzsNYF0I6OYu4jAZ97R4
C2xm+i0wvDVj9rfHsPfsXkgt77zjn/8JfG0Snaa1cZMm7iLRneTmwXXLf235tmDu
f0TdG5+4FwkhsOHe5+EQ55+FGuEl6q6BRUKMWB9pXZ81DuJOZdk3E+kVdK5VqEII
GSQyjbKEfBwTpmP7u5wXb/URlQsdJ+/NV7WZyVZIinM3v8Gf/FoxG+5HegryodCp
0M1vQgN7fejPm3Zcq2UxtcP0FwTGPTUYkx9u+o2qzIMC3QzICuovYmD4dOcKHPNE
JPe6DYRnWdAOqTGnREYS88BjvWuacyIySRJ69ZjeDFihdTPiXyVnM893ANAjJX6o
qhkW2wPgc3xRBEQWsATRU4IBXe4hd3Nf5raZbj3JCQRsFzONaC+H9veWQQhEdNuw
W0GghuKFm0OAqlurDa2T6gHeOmsiLoWBVkGC6BH+cnzjyDbpiCxgr5cb5N/ygob6
wR1w1ofCYNDqWcxwOzloEEGSq6idSl+qo74O0Fyc/DsVs9SbkWFrPuV3AnHCx7Jf
ssunSSqdsvdAN9aZ241Ap0oG9xQfLKx2q8k44rFxdNQoSxPxbnvNkH+Baq2rpy2a
EdCSkJzaml4hMkYyU8Zpi3dqXew/M33s4CXASIZ2bZCn9a2N19lb/7gp+aYb0TiZ
3mRFzsWi7Mp5kmnAR4bKWhYy9CW4GY/qT7uR3SkqYgDnbKsY1qurDZQrl0ATbPRm
PBt19oSVPVedwJFnU5FhHxS2PKQJv9Y06D6Go5LWRMFmOQDjg4Bd8bGmVM0/vXG8
HSe/AJMQk+kuECpJhH7+0dFQzIO8Rb5pqLZlN5NZ2qEUJO+p6l4fztjqMi8tM+aQ
VwZgNcH107WjEX/JR+BeOVjZkVjPPJNbzRp+oNhYgT8TAxk6YEInXmCvqMniBER/
XFhLfWQSvZNtYO6dcMQf9Ahn+ujQjgXSdg4jdYyS2H2oc5zZ75xVBmNX8vVSPUT4
4+082bSgV0JNq4FXRkUJJUg+zR+hFKVO44Ed4Ei60sM1JvmfTIj+oGKApcmLr9JF
sju2gsTPAO32LXORleuzNEETKTLz0vhvDNERtdEV2Nkr2kyiLcGK9TYi1Ar0ZeQn
FBsoAx1NXicZhsPoplY/tvpuiX7wDS4lHwXQtDws46jfWyNXy3bsI7n8cQGIyU4R
s29M50ko8jIw3UEmI2/GAxvoTcPxDQqBA9D7an6n5s2Q0hmQTuNis2YzJHhNXkXC
7JuDJWNpetHfwhbgvfLmPkIxMBbMwjqeuOsL8sUuD7NLO2S0wYCe44nyvCJpZIRa
G0V7ULSq2wQEsMwPHznifVcljkn5kgumiPsbiw7tgXXPxuzp7fucoKKFS/W2ZIPx
PObVfb9sqCLlL1lhbtOIwaKwQSzb7cLJrlcwb9gf9t8GOUOrBaIMf3fcq4BMGdZv
N7kfEXHc9l3YCbi/mm2YXD9Ko7Ij4EJH/Fzqemt0dvOepuGck4a0av40gRGGrX9S
w9NZjvYFxxS26bNXxNM8Mcw8nUMKRXTvffR9PAV1r1g+PaaZHZPjfqSS7eACLmBy
H6VekfZBEnySAO76Fd3MAAVD7OcDSTDwNAOjPcLBrE24W6/XypU0XPJ5r9NcUFQT
N5mzyfCrP1EX2Jxx2FhZhBabln4id+V2RWy6sJ9Owj8CGIOLR8D/YgDaGnqdsbB0
0U1GDd851UO7CgbpzkjYtnzBSnzoT1UvqnMIyADhG9Un7Lp4bVGYlueLkfI7WCVg
CaU1XQnQX5s51uWikhCyUXEtuthwYDRM8ef8BGFL9UvXXViHPnDFDS3X97lE0np6
HWlODTL5Yjc5/FUgsd88EqmWaFu6c6a4kioQ64nxMiArJHGWJmkFlpOIfdYAIbj5
ttRdVYc9PbxdfnWEEpklzhoMligAbiZdcL8HmsH0//8oi64JecztueJ6NOjV0Y/U
qWXNbzjfvEuJuLAg85SWauy1uKfj17diV4k8ironF6S+aYr5TgTMXepYhhyGECyk
X1gMXBQCw+gXr++9c5LRYuED7UQB2G19eTsDlSvr8qs5gkUYjpTG2J8iGq0kIJZj
GMod2guE3VSRswrdmHFBvLr24XkiQfawUpES7Y2fpHax4g86fbXDxmu0au/ltI9A
JlRCEpqyBqx12dezKr/OxeO0IjfcojVwxL5B7NEU0GQjuh2aii9AgDNXej2tFUDM
cXFCT5XSTwU6FHOevDO84/zximtDvuXJyrYZgEifLRUjKLK6zXGv27NxfMZ1odgi
9b2qgYgfKPQnciW96UlgoOTYS9ubfSsoO2s6PwlGX+a6h97iixPLRz3ZCY/HSmso
fKuZuDhVt++Jx3q1bYEfqTEl1tMkpF4VGVeZFWjkwoiiXCAAGhoZAsmA2v6ausG4
KTwWrc5Yygs626VQ+mEy+BOdjedDl4WIxqyZj9iUTKNbs4F2Q4rYSNcHmDmKwf6Z
ottzwcl61OR1JTcItEjzgag0J6Scbl+ySN2V2oB0q2qkfTCL3jSokTFP/+wa3SpO
fqVkBVYq9zVd9McEvvx5U+BTCXgp0/tq9od/mFKg38L/kY1wTUc06QW9PeeJqlJG
M/OE4Aty8W6oKpZu8LxH6Tgz/au776emoGD9ut5f/53+1nv1beLxMxEZ6+mGD2SH
kswlNcaKENZF8LmbEnuqa3FL0hXzK/9a1rakOmhKTwwYnFvHLSuLBwM49hHFNVnH
m2hIb5xJT2wX/TEfpRtlBsiOygMf/J+b2+AKLUi25Oc8KepbaZBZFYNsKVwPMhGT
gg+BqDZr8aiLr3//4c1/P3/7iEKmA9IAIMY9HKOsoYjL9DEUhg+rYeGorKj2kalv
sf0lo+yjE0ASCULPvxTaEADAamNNOV6bp8Y2cwgqFj1Zzt3XqkEI2jzXpNyAidT+
XYbfTZujZ+NcPeN6NxGeUXLu9vAqoHTJrATx+J9UG9iiSOyuKSPJdnGW0T9QBb30
9qtPRKLOTrLrBWEZRGcqB2k2yqrQ7rQiPSjBz/8WqWWHZWgY3esvlBEyDLX5JP5Z
SZjQyolkVJGYBa8QpTMQxk/05Lof4ud9dWZRPd/PtEyGLarqGGu9THmrHqY9Brny
iPOCIyGn+BX+B0YU0tFwzcWdqMUwyuEM8gpCfFrZGqviF3BvfEG6XK4j9grtIA2M
ln/X/uSvE4iZOcMwT5AvcnjK/s0kJi3pC7ahLLFvvJMAAXKb22tFrKpk9Q/BMmIU
IkupgcPeKawjhGhASTUQjZN27+ui7CKoT/oiDFD47LmEcxVGxJoE3rkIvfHijChB
lk4vU5jbT6k38s269gl6+Jfc02bvX04cwR+E29my7Oc8n1mKbVTh26pJwAKndNpI
qqlq4geGFcBHLAXxDLsCPGkBI66w4F+IKEvabfcLjqz/Ts3hN0wdoC4E3AH1n5tl
CZRfCehADbxabiPOf8aTu/l3zJJ4dlZei++lUmUtvWpm0BUD5VcE8Agd/r1PfTFS
+kRDFr2KwugynTCejMn+QHzmiUzXx/mf8vejn/PE0oO/AYUciLiPvq0VsKw3yxiv
Qj2N5P/qALOkHwGcz6kArVVoMploGfzPckETdJh/hcGHQWrJERFRZtj2mVMDwyD7
RY/Kz1NlA57ZfTbjJYeV37X07mJTCo9df7xWdnJy+LlBsTaefpnSyXH/dfPAifBy
V3ja9mBVMakL1yIgT8FuLJ+cvW0rOowDUFxzsIAH3++cPk1FMlnyluf+EfDJQgwA
un5VuC7nZwkMcjp1Jjnc97T/Ey63bCJb/b++Gxbpys4nV993+1kmz0BORMHNerDr
yVpTzBfMo6dvFOH3gQAl5zK4a8pnj3uWxyMR4hALCM3fLX2ANbsW+ilq++I+gHE6
XFKVR38FhiR8pKft2irDL0+K+Ti6uOVyU0rhvvr+We3wHueRITlY3HAQOruh6UKJ
XhgKXuT/nULRY3x0rR2uBd+Jv30M33H8lJxPbGdT0m/R6KqOcT7PO2O80axNStvf
Bo8snIxG85Xqt8oWzpWJOnv5c4ijZLTW2Sxxy6nQLOQWmNU+o22wEfpPIsBSUIHe
Gn1YOa/Wka/+oWFIJyadu6DLzHbNJ4n7MeXpV8JGiE5WMe3zvSgFDgwm7H9J0oAX
UCt4kFiNkdr6z1xVsQPF9xv0ViBvfe/Xa57u/dQmpmz3ZH5NQKT18gsfGdQzyQHV
QJ+hppJhKniakCpcp540Wbv+3ituA9RsFYPY7JUy78Ia4rLPH0JiRCWHLTMCrDQU
7kIUD01y4zAD92ACSV9NNwprenlxb6vsCZuvolWaUFuze9DawYQi1cupp3g+9zfl
VsAN/6W71UG4w4fYjfpJUPmwImi8SArlXug1dolY7lEYEaq6zQCpSl+HcN4e+wRz
lj9vtU4QE9+7qC5L++eU5Bm4x6f3/Dqk+coZr7KII+7Dkt9EHyfSO0rgatlLMTJi
4f1yuW3ghRDjILr2HfsdewjfW68WvSV/N4EbKo2HIXcBNue4Ajfr0Xdyz1d7GFTt
lPN8qFUTo4j1mTcQTioMViyauLaeFMiPpLqPFyZXhoQLuvqVrEhNKIxhtVPO/2YY
AsQ1hy9bCp4Ycg+VJdxifWzlfDws9GfddU1q6tq4IFviQSlfHRkWVOaJXwHWqfbZ
veA4xYHMTObzS8Bfh1+FO0+pBSYQVINnNq1UKxf1hb2H59djcdtKQMYuqsT8SElb
EVGK6Qr+I/zOkahNYK8XwQelGbh+9j/1HXA5F5cBW5lXcw5hYKwBsLZ2mrthwgOr
V2ublcxUhg2iwVPlIU0lWrKVPo+ocuq+Vuu/WvyUQ6nW646AxlIgnLrcje6QvwuR
bZjfecS4YF3nXA7IcZ/Sy3Zaf8vymqG/lYlu92LNE2ocviDjx7iOLEgadzPAfYZs
0E5YxoCVOKNwdNvJ5cUNwHdPVYfGy3xlFQPdYRS044q4ZvNmGJXdXNUvFnbMo1LS
+zjT9WcwQaMbVwPthkeuJjmnwJ2L6ixoGYIrWY/el9TDUw4jz7wox/iibIkwsXGO
VMpeNhm4buOcMtUBtH61d/xeloSCwuI89jQBMB4Q01wYAFAmjjIYpF0PQOEF7iz5
OMDFMweRTuu28s+bjgG9y5V8SW8Bh3b3tKYrdkPIXKCzQr8FWVRFLfAlnkxyPzMy
g+EYvvUDbT2ujdl9M7jteN+ypiZ7Tl3unQGYgGwprmzYiWvBkVsBRI7tnfYnoKw8
iMltZBzcoNHuemtQfhOvHGnvSzXK7godG/Ry0O/DTWzS4ZAU9qWL3EkfeLvyYRN5
/XXeQB1mqXO1bq8HBAemfBQsY6JSovxeXvjWYIflXn2P1AqMrKpOkyk96ADlHEaw
GAN1r7oMMAwCESICqCPkzz+PHgS77+KTjctrBKroFVpHr/qlH637FZUuAx7UcA4l
QYyyF/7WY157s/acvhc+p4a/o0xDBUA0ELqCIaJ/8R2r2VG5BW9sv/dQ7/iJ7yHS
23Z2TeiaXBIZPty6hoQE8M3Yd5XDFqkFO6EVluwZ0nqNl4KfMFMyIj+ZkEEeTptS
bnhM7w8fpAYb/O8Bqymea56W/bL8vvjm6SNM529jC0QuLa55Jwya7JShnwOfl4Cf
SCG5agR9q0/9KuAFelFvRYopB42jVXN3zulBI3UiwXBAmhBx9thnnl4G9ZHkyEJF
BoGY2DU0lwIHYUiwgTLxXsifOLvwGM+1vxO27bhpfh2zM8t/gB84jMAKDbOun5if
E6LmLAOxertuhfnLHTWef7MXfNjWYt1VfBDLmU8qjxelUl4qShUc69teiFBwXSzZ
FAXEa0xBqbnUFcq87riaSbx1YjARSky9m2WHUBdUC035IqBXbxiEIDcEgF/KxDUC
dKQQaW8oPCd4Y0AQb7CbjD1svj87MYt8g+TzU0ThZvEbigWSIW5+vxE/i2gt8pLO
xdKoQTVt1QUIJNFTJO89Ghd7vhrilmHaacqX08OMOvS85+nXy3raFGb+XMiZ1WZh
GpE/17jFa+6XzzPow1wujBhoK+oQXurq0CtZX/dZLz5cbtAJMvIIN7MrDdouaGrg
srqbE3bg4D1+9YkLjlj1LTczKVxEXrHy6LvW+pIWr6En9mAstdstU/m8QUb8uLfL
Jlqk/GRwICPUTaVjWW6HqzZYuhINDAGj7mh8QwjRBuyw7Zm0DjlC3zE4HCqKusGi
DsTGa76Ok7a15fB+DLMqMn12eyFHTQH9EuTXeZJxvC6QdB98dtjD1OlxQUCtOZEj
Sg3YFQxnv3PfbY89I97vOhKYht7sm3EOukj9YwH24CPpzXGh9NMCL9lUFVr7Xcgz
PihqhU8NOvxKHnzFXEWzhEngX486vP9J//D1IC3xr9JFygBYBatwyTxgaLUSUKQl
B4cYnhYZiMRrteFEI5TtyJLiQ+LAUwAVr2OKN/F2HHeqEmdDYrn/oCG2ipoqZU/m
/he0N9/ZasV/sDQz6xV3rZ+drmPTfyFeKtyMKT5CJGHe8/qkmXJ6m1+/+qOa8YPQ
m4HTmrditj5Aky6Dl/frWJxDM1f58bHMZvs+LWUrWKlsE+1YBSZtyNTI9XkGv19u
c/qc4I6iS+1qKQ3W2a0H+WcsHt67u1YcVfBOQpbNPF/obMz0DDHAyyHCVjMHu4W3
SJYX6MC/He89GuDf1Bk3/brZoux9zhhpiqTt4XY3xZ1P6W3p6Tple23aqWQCu/rT
h830SDmJSJXladO2W5sywMKXPj4z0Tz+eA/R/6nQxc/2QGT7Mge3JozRbqPl9DTM
9sbHNZGMRjk8YBnc9kjcpAuEAAq4h+N6eX/bhDyyO+pwK6Sgi5gaJMesb7F04Q+A
9EnM/Hwhv5VlEDzaMpoAl6BUSe+pB6xVQ44T/qS36b0ZNIeygSOjDJRxChAjx7be
XjWb+5TWBzGbMgSeu0oMFx5Tl+NtWf+he8YUDrx8no0VNoxYh+O5JdVVblA1I57J
+17OjMoplmS7MEhoJQfJhScY3zGCwAXPAD249onYb3VmO2BlW/QmZgTusEw+AhlV
KoZLedQfez+53W2hlFM1Mr4wZZ1k+pkElTULD8XmG4Le3McDdoScxty06FQI2udh
ev+IA7+ZuCIBIvEDdo2nEHeRDks+imrL9lVoIkV+R4ZNajQmHEoEmUcenzOLbZgY
ZhF6Vg3Z5rRgqEaKxlzuSN8tBPhDs8Js8823nBlThmlSul0SMYlssjpnaMtJP8+U
T4IvDlTqoK7sbVA8VwvWxDX1x7iP+Nb/q2QZCgUtkQiZRyLIuNlIIbbQdN57aNyo
P8pNkb1XLMwbRyMa3woEinZ93Bdb4Op5afLSnQ3giKm18efUkFPPtt2fBOq9nwo1
CjkPArsy/07t9Wt9Eu68erO3+taZM2LGtdbJ1gZRIjFP9btVd0uum5Pz1458cItF
hXvLfX5lueMEP4tTH678TSrzoFk6QAlkUiN0ONb4JFOn2TxHQGnTtkBQzmE5vPFk
sdS1PMA/T6+AUvVJ0kD5y+wPabd6npnlOf/3se4n2duvRfHOx5et46pTeDXZJfL3
SNtA5iTpC74aVI1SmjELgvWxz6Vn3Emqd8jJBuS7U9L5LWcH0Jtty/n/bi6z6W0r
0u1/tg1+fJeb53+jEJQHWJngvNZjPC4r2p+a+OeCzfHtcL9UaBhDCddIC5YERaRu
JPjfi1fBla/+4ek+ASHvJ/giuybbeK6aHU8oEEiX8KFsmppm2XSwcgvIbCwcwpQZ
4UHWr2rpJvNtUBIRy0yx+gM/1c4FD3n3GjchPwi3E6YF3IIXQsMNna2VzkPIb+mT
jikkBr9dTxYrkJTpsdIFlIYS4ZGjRkyDjPzCq0O5uaYvg6cHjeajtEt8JJIebaC6
8TPyYJnRyt4B/XnyQjfRFGq52J243DbHUg9u+L2jyMSpkoOiq7n7erYH5jk28xVJ
RmC6b51kjS/h2WEGwIFCsyQc6T2yHl2PKTEiuJrM0TD6ZqNfbGxDUU9KWz3qkwEF
iBj7ga5pOumlu7ewxAyF2qzfAfxIiRAewKi41PqOLumQn/5vgwXB+dU5wII3vl1q
Pev+QVwQqmV6p+prjBqQU7L8cyPisOGo+fGA908EM95TDyp9zA/oLfcCAoOOx/rJ
SEQJ0ROnyebS/uq0i9ARoUTLoJdy3rFglNoc54xay6lgonQKeQIkhMp0DWDV4hPr
vijdHjzJP+OGeZHaqtlJtFT1a81ebRhfBjhFvNuIP8MK717XOT76sy1cgSxurQhQ
js31Lcj/cZONzgd2d+faZ1aYPngxeqFCE+NafnkYFK6QvSyQVHb1Y9P4jdYvsucW
OkToq/W8izviSsKxoQRkU8mMEkqoo36HDOINIHO2o/mwHUv5/HD7kpUrYWd/gYN/
7ngzWPfWmVfIDPIzIOQBaMjwWBpzHLlVxqVUuov19r3mT7+X9jbGPliAhxoCNoq3
TaUARDBa0SAhGFovhWFI+gWp8yTNEvx1e+jVvv2mx2Tzg8EeBf2j3Ip52YpptUbF
dr5+gBGwy2xUQn1VOMeIUEsnQOUFtfgBBLpCwVA/paxuabfzBikDFWyRjTMTwFPu
Gmv6f9AKlxTqpSXfgSAl4oSKZh71VMxkFapMU/6Q2e/yLR99LNehJd5QvP+Z1A1x
cpHe9Zt8RaZvWFI4iVk8ytk8bWx/o+YMsSuWECI38NxXdTbUJX8x/lWQwnG7QkvJ
HcUfUOtlmiWaOWXntt6GLCSV+6S94K7Y+KVeQbslma0/Ht7oNaVZlRt+dYeEXz5N
7uSOMjsUa0mA70wsoa0sgtjgglTu3tDPdoqIFnEkKtWnZJUp3YOVSHDM8h8msTe8
u2+4xZQfn+IQKtSOQP3OnjZ/NzEiGuzcTKa7r9ZAruyAhjN/ismiMHw/Unt2eT9c
1AqHuqXPWQYd/Tb9JY8c/XSZod5gAgtGzDlw238qS/eDO1//SgHJo91+xp2ujSwM
6DXNT8k/pF3+NWr/Au1f4GgjAwJRp9y4rVHocqoDgDntKAbib0wUDpFBbgmBBB22
/WJ0YBi7nq4PApDQuGVQbbXRqqLHRG6IL2tn0qtw88yVQ0mKyChbfY+U7uysyi4H
tvFcMJUvqMWsoS7ZOig/1mvfv3tHY6iskOtSDbSuEl8FaNIfjXNYrKJ0bTfr8oZw
fEpo2uhOLrjcP31caN7RHbwIo/uvU6C6btkYWoUgDWHbekwfWZGIjPYkSubvWhaS
Nn+vt0wcmIgmceJ0K0CSM8gqA4I2FEw7uVZTbFAI6/5RbNR3iECAO+R2pdhIDPwt
ZKbGYMlwQmDxMeuK0jfz1ph93xkJHH0CV4Q0gXEqOh/UMHL8Rv7GnVdSY92d9qXb
7TM1RWjwIyPfQb4uBu9xQOGAIrFKiDJ0j47qG+J1ZcxoF2RF2BS63Z+SurzXdpVm
cuVS3wxDgGRvewMTk/k9PTTBFui2C3W3rdgnD9lD+x60f7UfkixgtDBkY8c/XDqa
gTkCtu8opsdnOvdTHrs5itx5hErMTINxU0xb0DGUWX7fq1hKlSg+WxUNbSZLbCYi
UryyRqsHmSFzYtsuNb9jm7SVeRLchCpl2+wRspKWuY2nf6EhEvhDkY68dIgDtE2K
gJ129zCAsTY1eYgdBnGkQ/FXPQY2J/+B/9k9eIj1n/hPZhJuumpZFfMfvRhVi92j
noNDTRBn8ipCQmrL97bKYbyzwYhMD5+tsujOsMfyEF8Lg9f0G3akictAWuZBXk3p
D874gBCLGxydGDUA869K91dQDC2rNs+Mdc+USS7WJVyABaM9fsbx1D0D5J2PczjP
Txixhoy5uxEaRKdpTfLP682IHQGykIa7N9VltLUgp9hwvC4cTDUciFDrjCQ6SjOH
giIOqLVk/JeCSKC+q0eTE6suopNH8XCvqgtuFXRh4oLaHRJCw+NeJMTNgK4DoRfd
oWLMTugbxBZfPeU3vvPyaikfGVDKQoS00RSdTt/zU+NEdKCWjmcRCDMBrGFIcj6b
gX7vnNy49ZJSvJAw1G7J2Ap29TQlg+R2O5P2fsq2aTaslE5LVbe53r73L0bUEmTp
0fTolTkqss+ZCPP/kkMnk/rdjlRsCJYMRdR+JxMjtr/3Ufx6sUv3tXyHfT8fyE7H
Y/BUeVgvKKaPJcEfHPpeu1EJw4M/BSkYO7xT+htd/PAPezchJ6Gq0OudTqfFMQmO
4G4yTXbyUBUguUBZitNEy3co8JD2HCrrwOl46dN6cbSXEYkdu4i6GBh3xxSB2Jey
UNW3cOic81R57vPkfkbEpSmk1tW6DnwkzkUec7iu22gxwt65J5rkTqrAy8IEav9S
4xAYXuKDU0k5HcF+zvXG3mcXawJ9JF6Z4TnPSMR5WVGUmASLtYbiJcCKmx3lWl6z
MnBoKDIKPgsQztl05kIzCEJH85xodP+2fDK9wysfHHP+qFi2odW/XoCAW8WnVyCL
XkJI8NCx2PSRh+jobm1dr59tc1s0tFxYFvqyHWXz4Q8MgUKQ/yfdzn3kCTuJlUTf
94tJaPWtAvwE04ZyZeyNbtSkS8DxT7t6lx0qcQlbhg+HrHQNYjF07Mpwmvv+6tEG
8ih33uRFmNEE/abukvYbi6MKHWuFpTgQqjBfeBw9hmPQ0kn/UJLXEepaeJKcQjdM
rhfA1KygwPbSZkhgsVrSGaNdYbld+p5qDUMi9MI6kSMy47CzLkus8lSWqf+zM3zJ
0VIWunTJCGCxnlzvEWaA8po+5ipelE5pdXVTFPtsG7GWGVPHu1SZi0P8oO3ABBRb
cAbjxGD3nBlmFdcelJDmXB9uE8dCmh5qGrsPpB/tbQO4WSX/OPQI9vs72YILJREZ
FXOJdxEX3cVLgFXpWHF1tLhVpZ2PTaPpUKxLfMdkSFP0h1w+twOKanEiL6USSwiX
8sl+Emeqzvz7JJi01Q33JzoVFpOoiaeVXMjoPBHxoyYubBRPPz05XajvrrKdc+u9
Zwrc9/BCzHpb/JWO7g/rcOJVdwJslTl8xBJLOszvFQsJBDUwGXeJmbpI4zHi1GNA
JFL+ek+JeuiKoN7QEy4+DPBV8jsDgWHtJbRNOHx/DpqsqpZyMAq34fT48XB55o2n
oHvG/dQUsujhaYWYOj8Xn8yTNyNf0BDzb46B5307LZg3EU7QvSnhKKcxdOcEApad
KobGfIIg4ZNMYEZ972kMQUDrBLgmyV+LGtrOt6QrGMfDp99nwsJ8R7i0Mo7y7N3L
PrVisAVcVFiVWQy6Jf7OG56/7liO6Y08WAPZPHUWa5tAmd85VNgNAhAZWcOCqOtZ
O5+S3/+/TqXR6IG8KL9ZgRANwxhKHkMPwCmuFOoLGZjbreIp/OEWqBjDE6Mymo8H
x7LmRlShnpOBRDCeQGSIMz0g0pecEmBglDbbYePCEhVbf9nan7a+j2FkQnXPkFsy
a/gfBZu76AbBlT7ghjBTyj1u36wEMERQrqO3M/H9ZX9JebLIZeIbeSUFziTgmPeO
FbmTsyfTMsv9tZcYygORHyVY/tKTpIiW6p4x2U37LzRLpLdvphK1x7pXsRYUyhFN
8qNcFZCWX4n4rlRoEElbQNUFt8hw3/huq7ipr7DYqiP0QXnkHK/0mVrWGcZHeHJT
FGn5gLEFcP+1/rCCtttVBNJJSxYGZHyq1zTAimBlZwBCdcDABej7icY+K0m+EoAT
5IL99K4Wezly6dMfZ5MlgcNEfCdnnHqrXoh+q/PcctsOdP3qM4+npAyVozNHr/x0
k5xpkn0EB+lTOc4goZCvGEIbPfurV+Axa6SC3bYz/4NHak2hlimf4W3jh8TIUdLM
Uv+TywWMVCZMfMrSGBEZ94JEulfJ3Q7Z0ybFixBAMvCDkGwc4ZBAylIq4fWGHRLn
vJfY4aieZnrXUD1TadIBvHhbMfc7+dQ6NDlMLHLwHYePuk1ktK/wst0YfP5Dyw7b
RcwR7sZR5pnm37/9nKqJik3o1dv6ckCK/ijK5/3BbyZZiVY03gRQl1yfYJtR7q9/
rNfP0RQA0ZI6FTbjJSGUiwnXpircpX6ouXH9wVi0nct6888ZPzxXlM3x7YpBwcAo
a4AifqfQaBAtDVu/Vid9twIlaOZ/wriU1t0smJOtnIG5rmzjqwZOi8mF5uWPoo+A
2fD1pDwaDm4R5k9BwDvpbqBK7XWdM15h54+NDvfJcfUEAya7NYZuZ8R4RKbzdiYY
1GekrUA93BSCeiCKoqzUWoOVSYtt4YchorNB1GMhNBPkR+a6g+EM1MDxDFUUlzvt
Hlzs++HcCPaBdStQeIlKMYVr/CanBNmFYTNG9Yr6krSIelCRSl1Ow/V2sxCX7yY8
n2HfCmpwzhZz6h7WJxPeXZnr0uV8yVBMM0BgWN5f/7henaeiXlaQ/XGs21gJQ3oT
lDBiITVIY3CBOcn9VV3zhe3OQ1Gv/mA/eKOiaVasNmhzZOCByVcynqQRmcPLMkXn
iGdkLR8WM+THl4v51c1kIcUvuLinKLCpgzG06R7IfcrgePH/afIyY3SmPFWmH76Q
BMua6xikSCsOORoOeujHOo4YX0KCx4Zqjq76VKwem/Spu8rPTA5c7brx0tWV3LeL
TDKds6RNZRr8mJoLQcShlEdYqiNP8lA6Wo1n7ndhCNNcAvMHTzIFeGQAQ/MdJI7d
BN7kskOgHzOudlRdckIbhx3n1Zh17YVpcG8xls3oQj/0GDodF3cswR2O8wWWwwBN
gFrLFc/afaIA+xnurd1LvOin370WvLZkZDfisgxCzPb1Qfp7OY3vl8UJQkqofOuk
vYKnyvqE9aT1od8t9Awwc8vAAhpMGA2gxcy17t6s1KmfSOsyEg31bZQhAFJ8kgZY
w5EB3Q1namP1cCoWsnbHghqAw5D/JSKwvlkp9GIB8Yc1am/XgsJxE3mJcSvnA6wM
uX6jSRreG4Mp77onZ4UEasqUCZpzhYZvsFxTIe69HoVwha4zOJfzsR80PZdIWARA
zMoFU4OyGEGNmoHJXRu1QtSeYPVJduFKiR3JuGyAJ0EeQMSAXCGTOY1sDuFGU0r6
lB15W9PlSzkOXGXFJhaeO+d+8EKwiuOCuwYrsLfBFDuFLdWQFgIP8TxQ2i+k3BUz
FD/x5uN/4sERQc0fFg8xLIoH7VTUGdtlpclck3ntq7LQhGWNAag84JLqxKgFKF77
GqPKh4TnULGuJvg6FVS1C2HedAisOcICs7U6pIEoWyzL4RKy3NQVwM4iTjEkTZUG
AG0ZLgP0V492ZaZsCgvJ9oiD+OV5alxPAKCSJBUgJnhBvY5HWTovBF6dgeLt9tAQ
+4KK6eU4Yb4q9jwEWbsFu7ffKvlz+dxhUx/BbllZL+SOzPP00Ewt8PK8C0kTsDOQ
K/QdRurl35YLiHPRuCY5aAavnAEUAWClUTHnSd+2uvX1DHJeT/NwwkmQ4FiI3ruV
1l7J8CbNAYiDmdPSIPfx/ViwKXbeoSlciZiAhOPh7F5Tzedk/maP2bM8KnpVUWM4
AGuK4AeSPwdOwpWcwe8siLaBN5RlyPBU3JJglDkz3PkxnYZQOWUxmlVhYo8l56d4
A7gPJH+mNwmhZcKxXLtZIGhYK4r7rnpbW1wSE90nMUmDGaxf4j9O3vEVYy24fGcX
0hoMJnwC1+fycohC4Ycwf9/yDzUmDpBrGMRr62vWn2bEnfLkiZ8HQ2hqGlZ011vP
n6XhouTToym5gFanLtJTnNx5Bm3FR1K37xeV9YFatH2iqxjyBE9ZJO4LN12nybGY
pEc9Uc/GuF+vfWnsjwHYnClaE+U1Wew3jVRHhV0t7XAreJ3Syoy9W3e8m1v7UOJj
uLWH5RlwKqPPiOmomJQS9wZVrePyE1DdTBYJKMn5icevlvRifQ33Lwm8kqt02WBP
9BvKxuBlVBjh1u8uZ7+wj+PHgu/i49oHjIvYwDlQ8/bKBk43B7FK8lxEmkvIg+/l
DH4W8jUd3OWgBnHDyzZZeHc6zyp0SxSKahjtUknvlA6Db3SZ7yHMHiitniKa1/Y0
SuSAImqSLT5laWeBH8xdP21V7JBCM54clpPDGvWIxRSKCP3OnCbjp8NoPHOZl/Vg
mQF6uzQQrDGg8gIQ0fgy5sa2v9+lhP7uN1gmkov1bNxesahO7siKDrERR+Cl+2dS
kaXXEmJWP1Qaq1HpfJ7cH33V8DRo9QmcVCbuX5+TgY7O1BFWrgtjDo2NvonX/zlv
6XmklWb35WAYLAY/uF4bBaC2lqC95WKS4K/88gY6/GSzE31wL0we0Rtdj1AApLjX
A9KDsBIpFmo05RTM0rajizZaCLGfB6E3DnBq2+R8jpv1FsJpGWLCyl6vmGx2jLM3
7HKj/rOfz+OgdRj08JMaCeg5XfJIm4EsyCW3zurH+lKhPHT5n+tWChdZzbt9VXQ1
ncNUk0uLODzUlMZnniYTN0dbGyVdEiFm9JuywShDV6Pt63vRN06q4zRfea9ASc+S
IfgRaiifmWM/05T553bIbByeVZYy3AT6nEXwwQ0iQwxDJ5BIGtkGdghgAoPiHVzZ
feiRVQg6PTdwMe88ncnQokTciomFNUOtYeMiJRXT4j1NXyJHD/yuS/HJp2M9V4mS
hb+8dHlTP2K5hOWSkUJXDi63BgfS/FOBpwG7AenKe0DeI/7XOsJ5NXbIBdRWdY4w
dKvTe2IUmD3+fAxzdtTU8rTTo+kxpFkKsz8jW9EQAkoKywUXCFkYSyYLW75yc0h3
4DV6uFP3Ch14vO2VXke8uBbBQDj5wldwSIZw0bKYWEuFriIBHMKcrHg8qP19roWz
etATs43NToRMof4BMeeYiSBJNeFppZeBKu2TJFK5N/OIuBAVsMQ1grvCxMvpPul8
itb2wXXRXsCCgNyYWSbSF/+JaXKvoQ/K0eFaJeKtxYk68vwdpViO2Dtfy4Ryext6
1JNNyKO16JbMmm6MC89YtJTviIjHi578f8G2bMTC+tCO+BvLfAEXRzexBAu0iFuP
RqUmZXSej52rtu0HOt+whjcXxlm190Q5hMYyzIYog0kZOi6bsPMajyjkesl0T83K
MxjWk6sQbrb7QzWRqEqHRj3dD9MJoWqgZBLix/ieYawQjjMsmqYV9Cl1K4z02PA+
OP2HQlhrTyoqwNybmE1WghLPsL7f4qIwcoMzI/jbGLe3LgxSz8+8wpnadZraaE7B
GRTWRHXCmpAWE3FH3JQ2d46gAv+zHTSx1EgPIaM+TlcTeFEeUg8s0ZkdvM8ncMP3
mm5YevxEkAqi/nZONBjQD0e0jVM1DScEKbxikuK74ujWw2wTjcThaiRFehKLnBqp
Tq/8lzou9oPA3h6cA/s/pw9KeijMeO7voPsjUHcWrc+pZ/zu7ulpTtBM4dI5LkvQ
QV/dMChYSlp9mFFzg6AlJL5mMVL6BFwbd9RV0AtG5JE8raS15HDVlhU3o3c2wmlw
dIbDGZ5xqOpTA3nn43kC6M8tRH6M/ptfFhrcN5F/Vtc0h5dtr3CxnsMG1NsdIiKu
u1UBYvi/PRbcYMw3XazMEqOsN33+w1uhgVvuxCsoVvpNAx6gI5MXfcqU08gaMwNj
l1kLZwcv8gSMZ8xGOUhQcJ1nA8hKEOr6GUoNbhJ7LdEi1VPIwEfK/6/l+vQsima7
7XkhO/J3vipcWDGRHZpnoWExeQP2/ysh/kB7kYPB0VjNA2L9aNiWMc1AnOwTIyQY
RVwMCgkt31dQbheNnDBOZ4QpwZr8IMOLVVsURf8ifnYfduqQBQb5ImhSCntxiTad
fcuJMpg7sXTUpmlOMhz93rm8rRzFnN3XBpp9PZ9tp/jlvWPLoXCZ9ltXoETqU1p+
mu6EH/x9R1VYAsFDtgaLN6bLyPc+z4tMjlrg3jkDzZuPkH9uv3uzRSOhwyb9atkH
oql7JeXALX42S/+pZXoVmRIPu3Q5V7h36oziKm/n7Ygcr2LhAtkdkYuN8s8y1YVJ
u4STHESOeDcddeNfrO8e+H5aIXCBhCe3bbtnWEIDiJd9Cs1DoyjcZQe0mvmIQ2KQ
kCNKBD2CV6oaKrZ4QFywQnX6/YOWl2pj62T/ZxOD5Vn1uOX2zYfMjJq0lBuprzw+
8ILpZtbpJo8cYVItca2QH7bQq9jJkH95UtJ3Sts+ZJsM6lZuKN2J6jR1nGRUS6Vk
/ikD8GjjDr/lQVkHiQSQ6uVzF01fWCeISrnngq69Bq01lpZPdkfokiOwORw4hJfG
XF1Jwgz3uXHpcUZDQ+Gev0QG6HCUwkZ1A7gPidlaDMwijin9SwUeRoqRW+I3eYTm
D+3latSfhBPQJkyTTBiLx1DiGfMITH0L/FCsL0ntsA/8dKoN8to7PHxuDbImGyNJ
hLUvkfWrdevzW/eQNNWwFH2m1M6bToNIW+5JT9MhTal0ouwUPT8bbPw2Lz7QEbwh
Dv8ZKcz4E4K8RfaAXPGmNARU7lTa6CHIbYPhd38TDmTM3G67nKX+lc64HY4N0wCf
itcr/gEkEGSTY7wn5aYrLXVHyLbMLyWveHogTLCLVhXWAnFt6U1JkD6V7IYOI80a
sgf2+25MchlIShEL56C8ujcy463owbaYgjqYt1Ty2KCiPWqXFRhpD9H5/jAtrwM0
8SzYvNYEV+UpS+o39vc0KGPTRK65uUfamDkOcOZi0dos8S126Hvo6S8O4UpDaBTu
LEL+THYSqcPXJ26r1dWiSoOG1bbTGZxGYWOwbpJExhuqqkIR/4Cygs2fKTlJwLvv
dpJrs5sqD63Iok2+TuwUNmAax9Ljyg6qod5kA4VuQfC55sKAnx1mLmQASTLRs4ax
JYHHLYHfc21vTG+2hkdf56TA2gWwA0/+Snn8L1hTfSz34LUz2fdjCHh2t0gaZE9Z
`protect END_PROTECTED
