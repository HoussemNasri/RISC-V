`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RaC2EfMcqdPk77cIQ+81C/cUYugB9I2IAplUA+w3ZNzmOwneRhCSJTOu8mV4+SQh
yONmKCE6+D+WweLM2bxkGsS1rBzmuMzXc0v9TEGEdMePxD+ol5gLtHukWl0mJaew
/1u5ry4ck5Gg9Kzecvta86/SMEzkNJ6lFbMFbz0aa0TlpWnan4L7oc/23rC08QgE
RZS6sQPex+7HCimdT5H8HFkCL13VcVIeIxEyrqGyRNfg8OSDirYp2Hdc3wBWn2He
FhVGqgOdlOd99fkkB2oeuvvpVQlLH/yf1klK97witT5bCzC619OplxBGsEL6QzfT
eD6cz3jSeoB2I05sPKHt8/dh3hdeFW56hxNkkli9OoxD2ikIgBOmEnAgyp8RqLd1
5Th0anOnu5BCegRike7bQo8EgbF3FFtPW30tzhSvU3AZzzfuydYh+566DNwR11oQ
aNB7VAaPGl8jlJ57mAzv5yHRWvicvtw0QbNk0Nz4m2NfjVvYMRxj58vwZrwFSW+J
gwXEFBn1dAjm0xI84LKpG6yruOjj+7d47BH7ZYPuxCc3jcPOZ5uFUZNZYAratWiw
MRA+adWEhHF+YA0tOsXOxGvdmawgGcLgDcv/ZivVlGKP+CvSY7wSblvYYDNv5yp2
5OZm9IMG7A48XwhZ4NKsJLl5qkCr+T0HQeqyPsVfLoGXh6iYpV7PXfMq10HvRIfB
uFbky08+vz39BbMcUVDD6tXne1Cj9wj22QpRe0C2avJq0iJ+vWrngDHnDpwYsUFn
e0VpGPmIQQV8H0bU93TaBaxMqUbFaeiTM+0ZJnAZT+e7g5YqcdJC7OCnXKWjmK2/
QegEFP/Ym8ONw+wz8d80/mEul3kpwUDGm2F6RJSBtF5fyLJtLUtFvxDqvc3M5NNy
YbjOL0tOGIRLatEPGv3G2H9oOBEQhnjFMXEQ9eFUSEUyTnhp8rzWAAmrtvIWqy5C
Te8iYEjaZZ7CeVdjHTA1uECT7vvQWOF/Ftd8XEDu5pcW5ETXtIx5yZMTlWkq0EnU
cFsZuuSKQ8iTp4svA+kSfVK8sy95vOyjU/BBEHvYtiYHPMCj5qaifI4Ddl4l5Snj
ioyeDgnaSVb1oTHwvBM6YG1ZfOlQyIyoHmMZYLdXULqsaaq6NkQKqorwkjzqW3d4
wt7y0cviTbCLQwfa8HxsX4NQIVCZZtHfIqzWoFO/6nwn6TEFJYuVjvNCN7xarSHW
EcolHtPSB1RZWrB+BAGF2qaPNPXcj+UWuZtuJDKsfcVsGNDeDc1TtTA+z+5zZGvg
KpzX45edUIp3T7NqutwL18ha/XJ0p/Wh/HxYAnQUPp8j1+bLrlTiJzxq0kkAyKtS
tGwb6dXRQ2UITfF9aTG6fTcBu1nu9xiF4mMxmUaT6IRQB6+wSylNMQn7wacHcTIn
OldVamedwMXeJlhV72U1qRcNcwPsm3Y14AJP0Jb4zl1XxAaYGVGzlo1WFxNdS5Jl
5pBpN043o2AU27DoH0ORfFf7e7iBh/i/tWTCAVsF1c505KcyTnlW1jJgdYEKd2Tc
9dwOmRMfsIdnJ45bQUEOk5De3t8fQykpCW4vlOqUiYR5wBVn3DyuU38DKmYo1wov
nY1JN7ImQKNKXYmFPf9yXIdVsenQET7nz4z01mI/0fzwKwXU1jcyQDG2ij+XRs/d
Z1VrY1Vhes4GLh0ZtHGyhUdVxYtR9zxRUozICzE7Q5PrnnHp5EiJezOTAxVhMby9
dRorW4AwjQ7JZbV8fmoWepiaPpSvG8oih9okI/0o5y1QAP3WIRObDiBY03qVets+
dGQdgVRQJRc4zql5j0jjpZfMoy0ffgt7fneluTRuH0rIcAd1VmqM4TGIt8P4EgsX
2JuFRMYqo0j8cyPj7mrlvYAZfv9PCIVja6pYWddvMaxv5oOWMKF3JG+xS5az823K
YHwIk70t6tJNhH6PPZjNz4PoOYmEpealVyC4rFQ4v82zjVKMG8e9hPvjNwjiZMBK
yBA+BKcyCtlt3HshdAFuQ3BXl1nb3ddTrvEB3Icnbj56JDtSOnbCe6JFAM89DJCi
PTbDzud0Gls21Ol7n9z/ESoHIyjLqYvUKyYlATOgNF8yVnlfI/q/cabvWLXKrKyz
J7Qz/Hrs1DH2czsiguhJ+Y+tQC1BNm+YYys/PEaVqRFiOGxHeR0/ZpVhXFLGPdW1
lBErGOGpuLEqWrXLK6nBom4kDao7mKei5n8qhXTqs53yd/IzW2pKml54YYfP9KF+
Mk52QvUJ7AXnfXa5VVvnvnDrCVXxeijbMqwoxHWbh/znGQTs/nrV5r/iEEkANZkc
UUMGIWU5IQTOKYMQsWZYVto9Rf9XH89YJq8TGcWVSGVYqpiJnEG3tfF9WRYFNaJi
`protect END_PROTECTED
