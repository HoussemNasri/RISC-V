`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4QX7n6jq48iBq+XUJMwqSzEAOxtcj4acJa1dg17m433Si4u8zQvdmWjwxckz6Mf5
ixc4+hd0JNOpJBKW17q4bNobRtp1BZRTCAt8F4pkOu7czwHuPSvivzb9NwvMkSrX
tqpqOpfKwuw+vaa6AvWstAdN6wOOtWc00nChK/2Zi+sRblrya+7B0y9Gkm4RHmin
mDpA9+e/X4m6iff00l8yhJmQqtLgcFA+u2MgELH1zm9w6hcg3ZTBUy703k40fUdi
3rsRItWpPm2vx8MS1mzq658aiFlg8/+AX4Db8P8x9vsRxBLGFCVpZScztL9sxCxd
C+Sub5KMh2H4jQwcxQvolDKaZ1XhY8ifi3JJN8Nuj+9QqCTHv4NrdH8QC6Gc9Ium
UB/JpEiv1wXF77k/DUxgtqBvnVK2NiGz0NoBiZk6XAmJSQTo/JtUSnvn04S15/hn
Da1cl1y+9MPduq3GU52HNNOXnJF/oju8L4zwe/thYK0gf+6O6hX5a3QpQBNeyE7j
ns26PoRPfBdcK0d+bRQTk9BtOM+eQhK4aBnPdaFlSSvf6RAs280ITJs98ak0zfr+
UWkszfBu3kxKaxJEsc0xoTY2u4t+HpXEAfK5E1PVVcfNk667x2mE3Pmp8pL0pElS
h9P9HYDGXQ/0VAhO5pqhiBuPesJ0wd+Vn5zTO0XVADZIkGgHzRfrvfLZ1A9Q5mxA
Smv3tJocLAloH6bHx0VIieuYJSoRTCXsP+YAXoStMnehmCs83LZbDkW6AQ7yHCZL
tWqNKiHGpAarmFkNZHPcMee4SEpcAtWPJWHQxMO2d+3b6XlJnHAvLwTvdgF3pfNe
iDZGgGpfRrv3UHvgfU/z6wfXhEcoNJNR66jNEmtg8zQfHOvIvs0OsCByYLczv1Ol
`protect END_PROTECTED
