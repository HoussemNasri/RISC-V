`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Y9cRyU2f7NgIbkqoCCvAIB6M7nKYa3mfE3is44/auWn6bnBdqDmcTQTJJ79uJwd
OdqE0SODosTjCBotEhCoMtitIyzbgGQwdnWfzn5KULbGDfj6AU19P0zugHtxeqUM
LAON7iQj0nojkXX5ou0YKoUHfv+3ZwnIjQfmzlkFNSBcFfWwI638Fe3v774ldHl+
MJNV1nXGlhtAD2dMuQSbZzuEGxHMZK1DGjLOyCb+ffSjZPyFOScusHJOA07J3mBD
M8syaWP+XhUhFSiZB6rZDh089Gg9f+n2aa/5zTxeoHf4yPWOOw1rclNJO8jSotwM
IHPiveNoX/TWy7K6+70UwdbY8MQR/6Yyx+SnUYH9LWmK7gHrNulD4merKF0R82f0
KgelVLcb3q/PrTDxr7JEp7WYSekvi4aaHgkbwyOT8m29hg4Y3tWRg9vgTV3UtBY0
YUK4xbSrqMHkP4vkTp3050nWrlAVfRq0rXfW1MMVrN43ycqwFslVtPYAoyaZEVVA
OSk2y+iXuk3q+i/Y3420AmgCmr5gKlP3on+Cd5PYcWxQSUvM6BOiAp4pC9FIybzl
f+vRvemmdnrONpW94WbbYEhFOc5hArU548rPz25hoe2s479ISFoNzrkw8d1kzKZZ
Aermqv3kUsqPpY5eiVFst5gB5GA0vgzs+U3gLQ8ZaxrOL0JUKzn2nABtqoFGkugZ
ZqHUxDT3a9vPjuWDcZBhdkFOt2E56mVPh/XfPTWmRdF6uuoFVO4Zzep+7W+oZfKn
5bQhU7gIiIMRX9quLobFAD7odUxkd4tvzvd0XwMnMv3GS9Q/wRDx44jKXkYPjRSX
cPvrWhhr+rVd6xHT8KTnwy5yw7jfMwgRyIApkjzdjrihLDp+Dnoi1OJuT7lY05Ah
PoBDy3bMtKpbhxJQYhicW7roHTrRUi6VZ7iKunSJpOLX/cIz19jgePTTjL0Lo3sy
R1lAk2SffMYU3tIhw+o1yVznR2TszHi3yXDjvABJVu8EmrkF5xgDf5CEC9Of8yrx
iXmmDYX2CD5MO/QAhxZbj5n+Ugzpkc6LE6ZGtRDF8je6AH/1J8u2BibBUQQk0ydB
KqS3cPM2SLawfGRnqoCn4EdG0+DQoQsHHgDiOC8k0XEvbRj9hHXGsUELT4vwiq9+
GvdPoHzrqNmWnJqYqQtA+Fyv3PcUPM5Y59BHQ+v42EQZR6uIyUFdXfcRCC/rGiyd
Mu6tr9qXywX9ArP8FPPD1ZP6REAyB+c3zjEQwB40G2aHKInOvhcNAUwDBSpUJWbR
JaVCG2+U8LsAVnQOdnp2I5nt2skg7EQWFLRNGgDhnX2d4dn4BnmAu9cy9K5duyIU
/xDPAida63EQMeAFt2xvBf54/gIBWrKtiKv5OSxVFa0Plf5x2Ds53RIN6qDGsteu
vHVe/thOQhX0GeNkim9Rg+YfZIJ8ETikE80fJOLQ3MWU535/3jsS9cZXswjEGsbm
CTrPnXcz7yhHhWrr3SzknI4L9LJsR7b6V0WfHgAthLi9ngWbGNj+kLz85mkpMitf
pTZx3zYj8wq9yIzQ+YeKqxAsSkxUT/daCrA/aR02pFTiYrd76S+0ohVrbMUUhgKg
8uwUIRGVok2B051TsGSd3UxfARVkHpB4dL6UQxh0N3LjCtZENBJjg4NNEliSiEkU
4TBYDwCPJmLKV/13aRH06ulG8IjQcW7BKDs6i2lIB4WuGKdkVI72c+u/ESOzLoi8
g3K0FYJMadfY/JU7buBE+Lp4vn3mpRzyW0JPJJD/Nbnu6kjOu4cEziHNquG+SxkY
fsxkyBtWP0QvRbo8HfLLw9TQRcaJEumYOf1fS8SgM46+pZ7HWfAP0Ah2GKAYzCTC
TDW+TkK6zOtjsj0Es/UcEEjbSNtp4c2r6JYLuTA4z5d1ryCeS6Ngoo+ZXdwuOUED
VSGWrFw5Qz714oRIuLxEF7FV3YKJb4wkpCp8Im4eQ/ADQn0BmIJ+f3c07joSZSTY
XNmHuZJmgr+j8Lrl6Z+jESylPVOJ+O+YEZ7zKGtlFA/uTnmNJHrzDseVMBE0tRu/
HfEPJZpOFSn4AhdeOCW9nCVQfKhL0McZeCXHqrdlZVI6DOH5deompYaCxwG07E//
IB0O2HzlER/ClcpI6k0fem91/6loZsxVRUTBNYQT/T05xOI9ZG4AY31zwcjy42s4
Yy1SigQZ1n4IRttcTsR/XPKTpp/44z5p49Qmc5XL6kDxkQWT7EeHTjeiI4Jm9JCs
BA/npltREE0gMM9skFpXFcR7mLLMRAxfcZKlgEDKYkaqIs/AT27/w5c1PSajAqyc
Zd5Pbh2d9DCV6r9HGf/hJx5iKqUfMtRx+T4vYlAleA0XLUn1ifuTOMaNIv0WWQdj
zQejb1pu4cMQ+c1xdOHmEZJNNAVKg27YQhfx3VfM1+hTkriWPfTgjbkisvgmwOsI
GTbj/Qg2PRltMT5LBm+FNsf/Mu/xLACIQZ1b55xCG79HYx0k4l+1XhTupju/CXQw
oSYUUF2tlEbg58G0U/XyFC7pvgIJ5/ymuI5m8Gyvybv331mZEsKNclPjc3MnaiiN
foHgRqEGftCquBuugJErR34pQzv//bZbL/vL+zeqnKqqO/MrLXEXTWphTVM9xvqF
INt473csk5HCTgwkuUpdQGcmbc7AC7DgYTNawNN5oCta5mFMu+5gti7mziKzTqAu
sXyVkuBmWNyQnJmiX/rIHVzVrD/N12vQpbAjBp4d1d/WfUA7Bq5llWoO07E8xsSN
ud/zMnwpAubrJs0ZMM446Vah+COWjwVQ9mwSOMgu0eukIU9HZGkokTNPKVk512PO
1HEeFbZJNlL5j3z6jRMa7JigRBcmvClsYaHhwQnJ5II7RDqrgNPLim+m+XwHm1Fb
9SztqvgfpvULLgTvV+dBtOOdbExLIaY1+1LApqnZ338dp7UrqUgyBumve5NdIs/e
zSoN+HnyESfI7WMc/rk9qbpT2uAxQJitbJwANGg4V6+IQNioQCBWZgfddtsTq2En
JmJzJ/2EHIgFvfYqGG2OeaA68tPpFcwpA5RaUMaP7lx0KqM0fG5bhi2lGJZ9xQ53
KVB+G8ZfGcq7W0N9GEH+a9n5h2VnAmpYx4/zJyCG59yr15uJQKqEM3muJ+vz9dLZ
zZxWyvvmHv8Jl0Ec0dIJYqaVNo6/mhi6o/pQSiBwzJPMofolrOYJUMBx5pJ+t9Mh
otDRELEi+wv9DlGJ6M/UtWw5bo6gqVNzaytGttpzqfjTNLKuvo2Ty4/ZTteonKmb
gkkJHSI+v2OAJxeq8GUdK92/Y6aP5EjLKTWoO6u7B0YfmaC0m5mtiuDVSslLSdSz
wkuz+cgSRS8bWyNt09lQXdr5baCMtR7THRzUKwVzxs6ORQhpJ+4e+NtiEhUEZ9SR
V7lrWkC3lwnuFnNwlgKt7vdiCBGomPFFc6ZpLrO1CRbBr4sFaNBmRBARCzUGZeSS
KCw3muJj5qZ1WJJ6IjG1PFGUdDI4asCDvhYpnaGQmk7FIe9c/q8SRm9PCh2MYrwI
F2SzuThtkqMZgT2yMZ2E/TE/aSzZx1UkNPPysZy9ncgnLUenJwdgwm1qoHXO5jI6
ip08HULRC6uefVXXy4zJvpXm0tvngmnZi2m0I9gARCj4tf8PCClNKsDO37s6jjyu
W+9zJgeyHAnsHOLF9msKZAoE0PBao4PP5Fai3VzPgJK5d0W8lInIVyEWVY+LwdLg
cObt5JSB8pCijERAnyyttg==
`protect END_PROTECTED
