`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nbi+ym+MKb8mbbVTjS8F/kUX0qTEFVFaksK0ySGCBcoqkPhRtAgVeIjOG5+B5DM7
zW4j70TO1KrBa4AyhMhnsTLE83Dz6KVlu+gXqsJ7nx2I22acmsnkBZcyLjjDPRQX
0zbnppmYzSpQW8F69H7u1IZVAEDoCwDx6+5oB1qouLyv6hwIHC565vf73cSaGlZz
RRkte6sUgnaYgP6rgQNNLrtsmPSPgCoi3CdHeA3BF6PiwDXuF8/1fk7k2e7Jx7qr
TVPT175oVMWcpVBqcS7rs3N9IcdxQamWZCNqfsHdWn6ftf131KSnHKwXOFgbELWy
pwEWnsoKyzuyATHlXFx0uZar/yZYrdnbJn09lp9zb2DVmDINTd5NNLyAgqRiG+Io
BFqV7oqkG1rD7u2zsYiM3T32KvkPfxYFQE5ebfflz6Za6lMm9lnL7OZ1VwMQj+4S
gaEvt4CJWAQHJ9Sk0W/Be/whEVmZBZBevC2Y029d1SQSdPwkQERriYnkdtIX3h4K
uOTW1EJRCgt+chHqv3xfTHaogxYSIZHtADruaZu8i4EBMO39IR1v34X4QKjM3ZTY
wom3Xs6QHcHcvaJY/3IQxgd2As2C5wQ3QQtBvCsm/h/3OpsrfmJrFA/BSPUHWXQG
A7Fe/7a2GGaA9dQ5tJ+Ltb1AX/wfVJR/cKZh+ICf/ZhSilT0HeGUl08Hbk4bCEBD
DASfLF63/tPDvMR1qpIytVMBbc4buhd9XaIY4ZmhhlyG42ad5ZqgscyL04SR062u
7B3N35I8Oz4SiMBZTAn0U37HlpPCTsb4RHCdN06pp71jkkP6DY/r5HQgei53t9L5
2wqhEQ7zjfSbaX/p0yUguNNNb8NprFrQO2nqGmXNRRnhnPzrClCzGQyvh0IZDeHB
V8PoTLAcJJYplARbcdhkXQC889iAHHuk+q8LbWNmXhTYzv2KkA2lvNDTGiXHogsr
Zj4ZOAK1CEtD1lOL0QBFv0ov16m7+Vr6p7MR80iM4vRRcNQ9GOLW3WrayC5fiRvR
vbCI0J7xDgT94xVfUe3YGyVm7RRVFNa7tXUr8Kcvm9oj7Q2NjaO99rLZ51oOCcZW
xJkVyzYKhCVPl1tFpBwQJ9FuSWHKVm9V8kL5/MCy22e0/PDcoy2L6egO284hPFMk
dsCOZoh9M07eOGZOpPacfuNVUtUpsVAY+DciSL2ZwHL5GZW+Sg1mIJoDV+kHZlXi
v9OrQcuIOWkcIcLH4VFZHkUi+67qUmzUoNgSr+ZPJJRVqX7Iq7o43sBi0ZMfPUOr
wFmqA6m8A50s4aanlcuir5Dhg2WwAUomZwQ4xiebm6yPcpjqH2YNAKXG5i7U5ptI
BRBAJ88HuSlV+B/jZzIZ4uxDPIyljTvj8BLAYp6z4H9SlwcB0fs7X6BYbRUbidnx
Sy9HoHIaEHpPTzIuiZYlZ3MD66l+KmaH0khJfL3N12NIFbpcOO/CnmdpFNP1hRRu
LAl+i0jSPDiegiatcxigOGADx/P4pytN6NDHTsIIGyjUSpqBIvmqQUTHXd6Tps+0
xWezqD1hiArNm2Rf4SzQcmRGLzSXFFOje5Lf9a/N2ppxMoSUHW4HFgTsgp7InkG4
gKWamRbUM2P8lerE8+bjU4Xl3kMMBUtPBVDvzQBJEz6SBqTpu1wsm6JwOzMF/byv
xlXFGmzwG6w1Uojw/LlXbLiCGSkTdc1ft1oMsmpv0CMa9dxCADeemaH96KrUjRHp
R5NOZ3/4zX6ohkFlCZ+CvN4K01RZ/PuG6q5bzhIFW1dVm+dCP/CetVapggALyMMc
NTSQfwCqYmH1l0OMxlF6jIqu39iu16Ch7QXxmdSCfuu52/kav30MOQvjzUO+YSU7
zN2SQCq9N1SRI6f+W2qpr30hnqAyEJrWcog5Ay5w7NNHiC3Q/x9oCL4sIZLl8VWO
GRanYOzzxNdPn3FvgYbJSkVFktlk8uiSVO+1iHCPco6qZ2bCRsgaomUfdb5/S0Ku
xG9fzgbXZgw+NSevoPcfxIO1jQszBRmJLZOwE8PB2QOvttKZkIQMn168KQ1SN5Ox
wMjJttd5cD5n8IjwGVEvhsQhic2/Tw9zpjbmlF59XngjYl96AHWmDIhSXyBKq+nT
dGxZ2Z00MD6xtVtoEfr4gbqTTV3pppHRnKCzrJf7SCGZuu97PcfsfdI6EGIj0kDo
KFiclwkYEUTqEaAJbYyN3U2aKrWsPFly6vJzIKnhIhoMtZjzK3WZrEvC+aUSCI4X
cUccBUBbBIAGB5qxGtK2lRg9hEubheO2hMewjOxbCUmh2IvbIXMq8JsvtrSZFIPO
MMyPbze7J9OZeNzdTQDV9/lgGXetDizU8BWclaFec9TUcLgI6dYNWRp0c91DlrcR
eM+0F5XsA1c83UIuCpyQHOWl7traewdINTErDjBqQHtX1i5nlLZMGbni06CScumx
6BbKQZIFxD6WSWrOqeuofhHE2leXKZ/QzTNsxXOywYNMExNiNom6EWKfCXgXHB/O
taqooDpECNJ+qhaCtuZ+mWEQ68NIUz7X3NMJrdbpQym09CdWXiQF+p7uyS73oCgq
Hvg0FzcZJ1NO1cMpMHrP+P3oOzO91ZfKARNn4YEBSMQ7zVpE3M0q6y0WDVKFv5BX
GwUyg0c33UYmxHgyhyCjOEyspbBLJOIn/QyYzSuWnL1Snhiw6cH3zQGrz2WXpFMj
e4COxyFdVKvVVfXrcIC45NwyaUCNRBvbrhmbxHks0milE+oMKEXeQYKJ0vtIWacS
8vYdqUIKh6FmPj/7m+Yb2Hl6kMjH6cUqOohPuGn+x1LIVHMJPFQhnrDOXwwRiyua
5ZMQ0Iru4Y9nYfWmrj99GipZ/CEWlx8YuAE6eK4cKOAqQgK1OBw6nSIl+FhpCLb5
K+2/jdmjPTr3XE2z/spnoAQuEA4QKhNpmjS7Jq7YYL9+wY0h2GnB53czIlqhBblJ
bGm5Bq2L/PFE07oYd0kPbbOG2NcVe0yaj9xJ5cF50NtioeIVfYbfwfUMVeEXt6bf
dAjITIFLmVYD/BmCLGSJO2MuWFcLfOV5ZZCydNuU+kQ9huj010LxZGrGtyRbW7pV
r1E4pNDSIZFh6L+fDdz658Pj2aC8wG0kmnjoyILKFdb/uyxCzEmsjz06hAv2POEy
l7hUmJQxCTMx2RVx14cpzlPb7q82okbaFnlhm2YGLdFyElE9tgHV05Ue0Iwz+0qs
c6WNN6o09EZLEK/05s61hv7UqobuR3D5QE+etUwLoP/RYSdfHzXzMvC1TjohaQEq
2t1VWlrzGaUE31vvip06m55jFTpj5zRgwRVaJLt6lnAi0vJluj03UroiX7hZw1WY
Yu2VXTzgQ9vnJhx20/1PjOKem4mCWv1ilMxQDW8QLRRYesQngxAO9hB8OQYgTFmU
BDjCm2TsO4FyxTI1Dme+Qnbg24iLExJQqbtIud720Rex89HC2yVrx0Y9vYzBYVTC
vz4kzkRWpV+8aN6lqqK0gcHf6rdxyNN1jqwfyKmLyNmcteG4tLtcyiNUZ83kZQXv
dnKdhyP4FwaKWcSokFo7nbV+OSxeohdNW70rxWTNB3LNBmb+LDQ13tXUf6myHHB7
kYQKX+eE7UCjPsP1Z1qbi8T6rCcQ/Rm92iloW5BPR4XmwgewPPxlLeCYZD18wjBs
N1ko645jyHRnbTFEylucoxprYl9O9AhbMEsKKeOhBfrDZZBBRV6MnOcXtV6T3vTv
YIO2oOJXeN2QbMXCRhMtml+J4VlOfRRCe03wvKwqhGnczFc2n5W5+6DOj5MV6GB/
D9caQI1BluiO27M5oqjXB53OQno8kbteZub9S+bjBAD7dGrJ2mCyJdfrulPP0rzM
VUeILQx4sGMRpL2CBp1JXsbJzhc1NtmRKt+lDcrZGYQRzlYpspiHjPbrIqrCXhrz
E3Tmuv7vj3EXZ7acDdSV+h5QSOL/Vui0HZ5hXrp+zzSTUPDU5WECp+2iNCBs8Pas
5IdXWM5glQJaBfXgWIkzZ7yo4aDPVaXaeyygliP1PLrFHtA+ePpVGYUeBPEFgkyo
vUvlUEQadh6RNgX997zHUbeVwo7Zz9o6dAPpmNv9hhDWBLClfU2D0WDPS81h4Q2C
ZN3hVTE1bI5CUJFbrJrauwzCz3pYLbaEzSiPrBrCZ7PBcAJSPvSuxXmuaVgSJx9D
ZA3QErYJ2EsiKoERmWWke1NRgn2TlkfbpVdn2qMqpU28n7vdD2hvqiBhLqPjgy2u
yN0vluEyPx7Lb56U4/4gVgXzIrDmXEoBfBsgmdT9Gpd6gblIE+K6SAvcrodO6Hhf
u3+q508+OIc7HtEnCM9fqKaFEbPzwhRpENduT1oWWATDB5PxTtV+MBseavwN0t61
yfXi6v9b4vzh6VZl4Skhwf+keQikEBDkkZigJFBbFk2LD6dAQ6+J7L9Yz8aEQF9h
ehF7sJaD49gJP/xDDgLd17em4KzAyNkmfn1KOLFKi+DPQVbulLKdqE7jx7NJCWlz
dzkc5CjgH1OTUfaqmvt0h0cWX4anwSPH3m7CBDr+5tTdfJ7rMm1qwUAiGMPdZEfL
CVmPhcMeTS+NIaX5GXpbJI2YKLICN43eoM7W4oQTkRFLO9qwctAg8Xw0TkLVYHIl
e6oj7x7PcOIxIe5KailXK3C0TXwdw3751B+JHLkrY04VSe7L9sjOt6IMGI2YwzS+
DkhjSkuHOjeOe5Ey5zB6oRpK77sRWUYx+KGGTmxYRP3EccfZQrc11jFZkBVRjMZm
AgzYOa/NSZeB1lgxVC/bYGGCDalWtyBbsIndhtS6QsALBWHqG05uyGOaSlm3k1Gh
iCjgPXxjKIOWdrFO/J0+jXeS55aejQGFBTQHKYuoJKdkE9ezB19KdAoO5+eiIIeX
Viqf+ikBRTfvMHgkeYCZyQaWCv4+5ILUlaHDXfQzRbsxcrg78T+dycvWCxhKmYyJ
fd7XcqJNI9dyW2wSnqsVBz2v555ZpdykgqVTwLlVSlyi6KZTzsR++9wGkkxevs0u
I6aCFtzt0tVEMVAsIciPQNVxZ8rtyAhCuKpKJbTgikP9ng4p9Np6hiYPHGyUVjbs
q7ZcSqyb3IbOmlYUeok9mAlQsrURLeZdmlL0vk9ucM3YFmFMoHrpmFqZM1L38mmE
/W/6fHrDl0SOPEHkgop5DJuiQF+q0EPWP4/xDxiRBPCQH0s631oz5c2mY4bG4AXz
dE2yuXRmhfFttkcHA6RYCkO0RyfcQBStj4sC3Ch1qQx/6wGtgwk+9y7BIqkx3UYK
suCNdX83LFkvbexnMAH8oUOhUSX/DnwN0IQSKMyIZXI7+08JTsQ4bO6bTiRnPYzD
LN0dYo480oiNdNIgfDY12sVt9tVig69EO6ACv0Fh5eCy2swkyNMlw2+GlOz/FCKH
AdZqv2wry0RvSLoeLocwXpftRM9M0YeKlOiteiIDyBIoMyGrAt6FfT9p/8v6r68G
eaFsR9LKIEFafaBO/tUjn79kwrUda0OmvH6tkOWZTDAGS8dW3R5FBG8el76CDGun
btGMzaJFPhMZgitXUqFf5Cj/w9a8Yy/Ojoz/mG1X2afY8x7nQRpEC2v/mmPeOnlM
4s0Z9tJcmbtW7fTkiJYddXzOvWEa8V2udvwrBj2IX86TDpF/B6DTGYPycFC0VLto
CtFGCOG4HiCc2lUGId+zBbzY//aLF2J7ZHuY+L6SCgH/sDIeBJxELpozhmIuFQsU
vtEtIF+PVjrBXUJhx4YixFzN4Ni1kf3J0JKb+sVrHZkYvYel40db7vr88QdEJQ0q
Gsv+26AdPRbXtVPOglWO69/HxXW56obQzr3v9lNAA9Zbu7mTAfO0UiQGbmtoauBH
eCscvsMS8pzVC8XIpBffJOxL8V+EkCgmA+HHWA6lsG0G+e1utWwdGzrFqQqDRGlu
mmGbxz/2NkPhIfxWjC4P5g4534yN4XlMyUSeAcYLFNM+HlWZIXGLippiSg2D12G3
OZxWgAusCIxLjLg1nAFYJlE/taFOl/erG1zDANYxQrDvU6CWQESV56u9JXu3B0wn
RfRgEhs3EbpAxjfm+9ikdj9k7Un77OOPYjOdNIAWb0mxjIY3kR3EOJe3WQmARU2n
zEm72Q/Fwv/yrKWpzmouMV6qGfg4vOrLEGZNReJp4xFBNPudL+WFBI4W9BRwMEJr
YHkqwpez0LADNgqp3kt2rAgK060UulD2N6z/UhR4KDxcEAFb6k8GytJ0TPeray/x
NTszrURd8U+GasikNQ+QDANrPBC3isY5rxJ76wzenspfW7FdPSfI5sxCmPz1o11w
9XoISsHIO+/Xf6z4Hr++W6Rv3sE8oWzfVekpZbFesqspuV7oIEtHtZOTWa/OP+EU
WHu/kWrOlBga+sB5pUyW4ExBMr2LE8zrw/ENaAEiiFW12gOmB+rmZCnpXA1wJpxs
w9RS0NtLF9LTpiVITOhBv/vFPBLg/jWTW4q6xB2FrMMtHgQXjrrqGCVaF7+IQxK8
DLSBheTWIGSyHaJIlHIZd9IqL+j0uMfR8e5u3ty9goYWABX0kNPnTj4lWW0d3RMx
JuCMchpUc3aDLBTBYSs0ZJ0x9zFU8z9MEcX4oy0WqhIMBeQMIe46WqLrqU8jmoz9
D98hmxh92A+DX4i39ShbQXdz5ZaUDHpycP3Y1FuAkAGfbRT2oj4LekFLqFXZSSjn
6PMnbmfo4Jx4fQDxhiJooHaX2gzXPDmwGQhECeCRI6knYXEW5sao8QN9fNC8P616
v0F40kR3ZONBbytv975zwsKMV4AuspvRbPiKgKIn4eSJnrUWENOcXDjSiDpMRe9B
H7oiw2zO4o8pkHL5Y3bUudt3dRsSrBzj4rPdqaO4hyC8wT92pRQb34I84FyolgiY
ZyZRp/quIdPSL+AJ+87nNYQOEVbujqnCtt0Fqij2HmAokOZvpwVCkkZb/r5muhs/
tEYNEp0g5r+qieO5Hgx+fiO83Q1RrOeV/umWBRPtlrSMDAc1dgLS3+mqAOSUed9x
STu0w4lY2MNTZAdO2Auf74QSXQtgHVVyswj8SM/xGIY922UW/KxgXFX/nCJM/FE2
v4jHeTBY8fqeO/sIGfGVfFiLA88t7nrzH87FStb4u/mfptN2S51PGwsa3d87e31S
zgQeBR0aYUHD0vKuyQ7ex0CTmp1jWBST+SewoTb2WZuHcEGJWMfq8tZ1RLA9y268
93u/bYvd5rkDItaRpruuNVnkmMmeWDbOnp74Ram6E/yKuvxP6ZQ1l2x/BP8Xl2tm
LA2UHTw7LhNtXNQfK1ctnHZFbpQsXYvTeos2usbtubXeZmLUKwHrmKIJFGE2iLQ6
kjmm32rhd4rLKRKKNWT3Tw==
`protect END_PROTECTED
