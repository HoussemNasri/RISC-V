`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4K4ir6G64FLbgJOKzVCJkscp2DzGvpgj88zwtRKliNmDn8OYM2zptF/LQD1SAkr
gVztz14Ezc1SKbGwB0ch9SbMKVWZWLJ+OupXhdp6r/Mds5NQiBE3krE3bTVBbCMc
lHdLkkap+KHTaWRR2YGmLSqV81O7tOlh0xBXsAESsZv1TuHNVa/pG6PEDVeEOBSu
`protect END_PROTECTED
