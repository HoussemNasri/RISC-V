`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6piFKuew87FB6E18KaENWOGqb+PtnoNPZC9RDIczF3/2LQPPluTctPaCq0xiLhDs
gOULbXRD1yW4egNU/3Kw40yczs9Gy2luix+I5MDJx1iVGywvhPYq60PxFFisYLex
CoQKC5se9out5wrpBfwNpq7DsLVn5pat3ijfWl1UCe2rZ0Y1Hi3tiN8fCocpkU3B
Gs4tH2US7Cv7DplA+YQKhhzkHsPtt2i8PBino5WsmZNJt4VkFoW8c8a8RzPt5qW8
sddrdw3qM5h92JcCSHdVAlsq+AnQEaEOdUfiktOYT8rpoBT4C9EDASu+xulqy1/Z
q3gsJBhysc7gpmguiJ+dQgIwRNJ27WGLZJJ591zne26iZ2/Nr4Oe+0Bifg9Qcbbz
sFrXCncqQDwbTv/4hibXRQZwWf/Tv7etBbv5JjjUqPU=
`protect END_PROTECTED
