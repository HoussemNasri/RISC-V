`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETJByMzXqK5m/MpmPlN4PzC9fRT4tEMvZvm9VIuY/0Lqjj8ITig4O5+6d/SZHj63
chvUkLLCRPH3hTKDSrl7DQXOiOhUGF7G7brtOO76j2qVASBzFwVgwdzQ1KQ+GKz8
GW6v/RhzSgpR4JHLSAvmU/ooeWE8mw8m4ofHBSKjioSlryymw7q2qsucNczdu+Kz
Hs9ZfMygxvaP8/IgTrQrFZBifG0TYHh8xROguNA+icafNzS2TqgaoQuNtXqxav0j
b5Y4iMdgg903BZZkcHEINWbHXH8js3IBaBZfy2XVjnuHggZwvx0R0R8o8Yb4otAz
mVK/4q7lSCAFtDODkB04lapZHXg/90FiO12kivDz7wLhA4NVbe15gT4q3vd5U7UO
DIQyShYm5K8V/qV7CNx0DDSemJfBqG8aMLMmHvdsf+ZKRYqaGJ6BQxvKQng1ut1I
mbqIucZXCdoQ3rrhg5bVsNqPFDucajffvUtGJLS5CbFx7Xi3P2DXL7OYzSBwuWBS
kRxoS2dsp1Y8QoRzQ6GwGT9LDd23HKnHHvzDtXi9hGxFXHgF+0R0qkpEHMetsW/n
WzS2alJJfKl+C7uJx3qfcXPsrn6PKH8Zjw0whsRQaVOrtH9srouSDSRcpCmqHB1b
QKb7fMsIfGWUg2MSAn2YmP/MhR0gvi4CNPtbR/UE8nMZ1vMYc3blSgRQhSaVgXVm
nvSrjqn2dtKbWW4Hbs6goe8d7N0mnTQniZGbzMi6QUhNS5Wm8XPHs+GFiEgIcIq6
3a/S11rcY4WbUDtDzdK539o3id/VanTzGlaRpjx7Pqhs9hBpc61d9pnhp7wPTnkO
iwK7xbMfkjL6jzXouQYKaD0Ctf0w3sNf/6sYpTA208aREYapQnRWD38/i3Vt0qXp
Q3bGA0KnY9Vwc0u88nb36pBm7eWi9q//q1HQod5t/H1VAAfSKVvPUeQDXg9271W/
f4S8pE1xb7yqDiF3F50GsRmAN5O2JblXDT5wlBDLqA40gKle6Q3o2HtACmDmMVDV
lh3XWpwlq/BFSMtnoh1oOcvbEhd1D08bGMiRcvKpQ8MjuaxMB080aATLw558q9cQ
MhQ5+Q6515k7GKFUu8hfafuYE/EbmXIiebLc02Bn2oanyPP3AQEgaoYzRCccUeJI
wHVa5r2F+ZU6khyVa10SoCtXX/pvjm3S+aUa+AzAxruG429eDuA19iZKbBzedn00
A0YHTJ+gLhr482SzAy+jwMx9X0Dy3+8eab2plIoFxVjfO7V0goimmazC1oMtRlte
`protect END_PROTECTED
