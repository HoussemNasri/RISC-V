`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXah3Umfl1A/9rWyVmfW+jNTqsnvny3WHeA23s5GgBMIzftUex6gVX7PNHahEZIM
ro+vk2DoUWikFHkhrkxxHHZXIgsPIqKCGrvyS68+UM2/SqWahA5DR7r7mVoSxGmr
nafnMAwzjq/giHpnZBXEE4c/w/j/VnUstX94oG9j7KdrbwgHX5FcsiODNgEpRNXP
rYLdCZRfBcJJWSBbZXjx/irenHoNJhIaG8NT9AZEZTic0evkAyBKDMtpjt+D3yLK
LVm5OZrFVqxiEqiv2Zc7C/iYfGaHaVEKO80kcOGGbk/2z0qpvU6t+73Bqu6m9YUQ
jQp0WwANBIbnr1PJmNNjb44aP1ThH0Nr1IxI7n3fw+6PU45KYzT4swaBpNc8aylE
JsKvDyn9ZtnRF4WaHT1zsqfGATp3MQVEVrc6E3LkIMwKt3E+lsWbU96QlkOfdFYx
8VynMTBDKDOT6I0chWWIrEAN9Gi9eT/4VH6R3eCFFAETmWpgqJqX6B7BbrudhTXN
1FBMZFNJJGR7fp6WplVj2ZlCHPADAAyn1uEDy3B8oK5Q2bGVaaZYENoMRqaW0sT9
onTdThnw83E+XkVhc7ROft5XOsKLrje6tHamZjGYQbHnZ4H0VZRGMRHMBvcFYY8l
++DbBCokk0MHm3RWB9VVwVskKCL/qkin8ZMFdYbCZlemUBN2CBkmEhtmSKx1nzG7
DI8qbeHFZUm2KNiZza7BayzGqzz/TUs1cJqOhsIv75oyblRNMlw1JHpfMMZBGcSg
y2Kmg4s4FrxYf0zbMOzTdTNUQFg5KnmYoHYg4nZUNXboCHgRDkBk9lG4q00F/5XV
XXAxNpbXltoLGP9Cmdbwzgu8SmhrapagAPpTAZgH1lzGkXocLiACIOLfECAj2MWM
ZnkbLw23U3OhsBhgtV8rxcdr+YHxxcV2I/09srJq3ilasEOY03EjQJMmqyk8g2lH
FLemWrTKgQ31+rde/VnUQSbpmJBm1W4blmVkMzuzC+o9q7NQbrzvthnZfevmAA68
3xU06Jlz1frP0AjO4wByhKuQC/r6+zdm8Ij35bBLPNGRwEfVCwNZNWBIc97lvAub
Y+n3iVla8MigNXPS+gvauWow299zTQKx/VlrrZIulga7tMyQL7a98TybfxpwYhjx
kprKO6dMS4HaDHAMcTAHDsa5Tj93XIPaBdrFiJtifOoOMAPdeMHdDu38toNrloXu
Rc6eOI+U6ghUCArRRWC9pHpZTU9NEa8Mf2hKoYYA+tSEguZPeoMbKZK8+cG4aUmP
w2U3cp+ImREIX5VbihPs0Hn45g9s9hnX/U9vD3XjPiH25uGTThwS8jKyLW9MPKu0
cCxJdrPwpS6I7ym5lWdKxo+ICKNU6xJjzDZ1AtKosQbMWfFc70K2HIAUNYirx0uT
XoL2agLuUzYDYrxn0twSgQX+oMLU0ka/10OkXsGX1aTfVVvLQWGfLJ0AnpoAp7US
o6Q35OevfKFA74voV3NmYrr0eFnyLU4ejnKuE51CAVa+Nb9h0Ii3nrwQWrw+2y4y
6jE8ltPIapPLpRP+xiUOwxi2NWAdPZFD86MR4YR94VE=
`protect END_PROTECTED
