`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYf2WEmB8GBQSA+8ZOzwSWCUCbQUcqTMQN3m1uYs6OzBq2UVGJ7kqfGiqHMc7H9d
P5IkaLwwglgvQTxJnAUQkdReBQYzTUlYXZrBgvXniZC75wlQp2iOAF5H6FGx9OPp
EaXMB2nNuObBQPjbzaJ78SWBgzZVeET3kV80lJVRIwl+caaGmbCLsV1Ql7T2+g0o
YdnQkRqwr60iU20D1V6gn9+PNak6y56f4qZsNlTC9sWnWTDLVXWngknQ8I7Luew7
4/Hdq3QsYU6qRccXAwRBw+ahiZc5UGj1FdrJFSjXY4ZukxZFh3yQhC/PVu0x8ws3
EViRe540x+e6mlJsSrueXdTjbGCutkqib/w7RNeUyYgMcvfav0Y96v6AOs7ATrJD
wG+hvJxLsu9VMv3Yt1hDT43zCYRbKmL8IQXs3ZVzu3LssF08Pp/vVbtUwL2sfcDu
jC04ZwgGoXTPlTgRivecF1LsCN7+7Umpn+ZrzRiMIagfNwMRN5HBI5YcYAXzLFDn
7lY+3N4azEjqLg6hDVdZrryslnjpeXoiFx8SYyX87ATJVH34yuvYleQ2mk1jjlro
oLA36mscNgz8Iy32qnU6GrwYIgJzj6gOMY4sT6vik2NsGfT3u07jc0zb6XiHTScB
wvybO6B7skiky5ErZlF13IV8eAa21kfcAy/RfLrBwBJNVpT05yKpRzr27RGGtyRm
QQA4pKaUvDN0+w7fD4W7Rn/EoW593UjJmhpxysmiaVSSOVieWbnTqCU2XQ023VFt
r3B3h2Y5Sg0oo6jc04OBan45G6DjYiPgB8+PJiv1vduAPkS0+y1rlkL0uHSa3F38
siNv56Q5gP64f/E2pWR6EMVBgJYCGaW4HesqKtVtwtRfGLc86zDX7V2cGOKdnKuM
fBm4UQ2mqnuZEOrjLG0gtMmmG30eZJD1Tl0im8EVvCWSuHJbcPg8nfduP1zaPLsC
16QbicXoEUX8TBkUNIRQUbtIDJ+JC5uSQ/ToxCkeCFgncT2Q86KEwkgraRVpEbUK
boYRatQmpeeORE/cdkPyE8lADZAyBLadK/QKkV/BgwbsGnMO75IEyfa9OhkxnMrV
viLIvq+fsvSA91VPK73qzzeJOujKiT48xhsx4E9GtUowEACwUe7CyoTRDS5znA4N
BBBAxc5/CKREYjTi+/9XP8XDmzYatBG6ylnULcNEY+GeRsZobMFhXn3Gl+QYTlHV
rYFo4lLn6LlY5bE0tI66EBNzac6KGLd28sZHtU78u4XjvELx0Rklhc+sNFxc3OEN
f/3G7T5nW+NphzWDe7BY5i7XD7/WI9PfY4l6ZraYsBLgtZ5skexV2zxQMRji429X
qg1RhdlrjlX2GdDdKdvXIiuUXgyJ9LFrkHL28VHTuUG2eH3a76nmR/by/HhMEJpq
M0nV1gSFGw3fa+ao92qzZgYDr0SJx3TegSUeVryZAh1VpHfxQF1jC7vCGbDpx0w+
`protect END_PROTECTED
