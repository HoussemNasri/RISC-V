`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ErYfou1qD5KSgFC6PD5D6OAj0eP77r4N9fHM1/LcJHtmPAxxtTXc2Gywahi1ogyo
0OxryEOEF0jlExyL89wi33DWa+lZ/CvdwboDmDFmdjDyZtcIszcPqrd2U4v1iPTy
+NjiFkfvZmGdWCE7K4fz+/SAWEiSkZAfFzfS9ol4eS5WPu1WVVnN+PAi50BLG6DX
X1MPJxqjcOSretpLZaYFqwMYPx9ckg3pA/RZ7MyXtquQLTB3Umg2cfS5vwLwspyB
WbtAJszZc75YdwhSeg3MyLy+hzxw73PfTaVzv9z8T7Mp8Us5XD64m0oOwcrB4++B
IpeCpHu0+LSTXqkVse+vyY7QtIsGCjBb+RylUFcrAYGTVIozJoP/3RQbsATxsJyq
sop0IlMT+bX043xFlz24ROIme8Vecp7VGOdJbqmOp3NbXmcq+QrDgr7zVRgKZ1op
vdo7ZCjDeIanxc2Xy+G0A20y6XrHQbEUfZ5j0aJH490lYCFGZYbW/xsscn3tOHtZ
anFls0wX2S8dCzwEqU3WrcnTzKAgtxbT1J6jx6u9Sqo+ySz4eTgQN6rkgQ735DyO
cuFTARNqVENPSBYOGBVMIjKnr9BClgOohRCBWWSOToTDKdFzgHariVGMtAKWNEpm
DxBwBixq7w0eBN7MJGb1zFnLar+jaf7LQLeS5c7qd0eDtbpuqTK6XlRWGHicVjiS
8hCiLKbq2lscFg3ZAMR/ZP8qYTtB7j0u4Z2wHH1Iqhv9FvxH6a/ntKg0p5BY22VU
CkH7Sb8atR4Ac/ehCnWKT8yoFY3jKkbtuea2nqG+OpHUwhiULhaI3bhz8KmNKtpp
BBnuuH4UQJ/MazTWwkH/SwiVAQLIK47TEkoABbgexb5ARYcED/KXmNd8Z/p7L112
cUH12AJ/H201DMVp7mvq0S8bIreSALDZTsuVwh/NHkSBCp1tpZK63RxkZ2JCkGwg
1fIideQhMhzYjryvbEi6OUbdBMYgbaVga5UgKMVhb/az0WvypUSYc4zJBSna9ybd
nOmcTuA9FtvRaSDBH7PwgBZQD38P/+F4z8bhkqbWqENhkQee2IVqFogJ/C7jkD0n
`protect END_PROTECTED
