`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5T+k9Df8QhnzgAHzgaaqxzU+Tpvvf+jHXP5Wv69kQ/Vshb0wUzu2NnnSO9vl1Ohs
R/qAvcsOPfBjFexFVvr7nuLn+QeuS18KpcmqMtKSbPlXymQWjrcy+04M4dzjq+Pd
Q40Ls93jN9jCHtXsW8Cg5zLP95lou3cuh6xgv1k+TErEovZnr0qlnL875nUpWNre
pK/G38FdjKeAF20RoM/3NFRI8VCasDkEmioJPR2uVvAK/wKYP3B0J0MDhOQA2s2V
EIk9fF3OOh5tIX0LwapmRgao2fnG/UxlvzaNpPThAxHRssuL8uH2XPYx7b7f8k2u
dWJuA271TOS4v79PCnv+NmLiwc6iJVHa8qZqd13NM1TCEZ2Tekqjs6GNaK3ROMZA
A/b2pNIB+ivJWOPJRBX/ecmNCvmXXYa/4IuSxZROuQ2OsiEEqWWljKYAS5xn/0Bu
5voZUEsF4H/mhprOmpljL+tSWDNsWx0GX7L1/pwbTXbRv/WjFRH4hqCInc0H50VF
sEzubBAgQFwbRXy+AkFRPxtl47lvUf9ApGaCcq4IywiEowCKdJ0w1hXkrvvzeqzd
UHsEfV2BugFasB9GeL/divpbJXEPIKpm3fAlXZmmZwZ6X3oc9AWz1+JYm53hvBVH
n/M7bdXfUFZTkNg2e4UsRPyom3Hr08gn2vce6HBSlXLkRMZ5CqPbpc35c+QW/Xuo
yyB9Rd3tH2UGavEJAC0ZPzNMKeDn9YjddmVeoBBmGsiIYGV6JSnavxYGfq3x/O85
POq21wRC4vmVdLEaPtoZEJIad4xIly5PovxVI5xY7s0eoZBCN+AAj7kzmm/RZX8P
VcouNayFesJzbmaiNxnkbkEiZui1PTJmDfjprWS4l598gHnwnijTfMm6HIhWkgIs
OJYm/SIcjJG+v36O5Z5OCNadJishUKjFqKI5qze6k6VN3f/nQBr4EsllKBVgrask
61AHR2nmtJk0aRFEzxkxjaGGPlNoDbz/5ieittaZfn0p/5C8d/XnQdePPYT+NYgn
Js5q1zVOkpk29c4Y7uO5cPH3V1jRQ2CS+jnSXdzn0PX4mSqZy+DiOOaQVvTmS1oS
SZUI8uyUbZQYJNW/nqFkeunDq/aasJyCvhad/9okFMpUc3jZvbtFJLThv7o+dFkA
zaWdnG6HcgkMgoqVMNC6iTI8hbPmLRSfJLY01rzbYIUbOPiTfLW4NlJ4uwIKsqTI
/5NGiF7O+tRfHjPJUdERCbTnZrb+peo8H+G90prC1LPxtD7OadzpPKEkKiYBGBW2
`protect END_PROTECTED
