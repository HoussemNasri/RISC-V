`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Ht4oV/50HI0DbuJty1DiTf/dxdXRlaOVrSyM5LD/gSxDhU2654ekfmdEwQEKcxU
p6rio0y7QniYtCyQ6Vmlh8oBN/GU4DOJHF+vV8AK8Sy9f8xty9wzQfF5C8VHT/hb
DAAMF+wtifPxH6k5XKrcYpKjIi+TxFL6SzPKJk6hoinX9hwZQRpjA52E7R+kY534
ceytVdythMF5gagpEA9RTmHI+qbUM1UKQjY4Wwk70njucct61e+/73KaBnlm2rkz
A+G2swUqqnfSBKBI9zYR1duZbUr/9zm5dWqnZzNOgth2dS5bAhjQ7F6oWNBUJrvD
0m15IkF4WvutxeUsj+jCvN+rqqHOxTVdZ4bVWD6JFrSTdOOExgjHtZWwYJjjdtj/
d0/gbyWUObOzinwLJwad4m325NuIW0gf6EwmKYo2bE3MihvPrVLtxqWBXH5CsXnG
3s2VC38alykWypCTN5ab2HxBXo73CaPrxk+i1bZxu5tMTXnIebyvgXntYST7Hu8Y
lXjuJznhmE36Hj6GNo4d6USH7eTWGgSoV6eHgZu3BJ7IjT0qLJrXk/6Nfzhu5AyT
lc+6YnbRB/Kjl1J0jJjeVJ8YXtZZNqVX1LydL3KLxEjgmnh0LNm3a7nx5YuAUkLo
gIQF1dLEabWDg7x8E4VqljJinYkWkfFMX0DnD0+VyB1rkaxdi0k8LRHh21jdBx1T
+O8zenRScFvGFE4Ribj3IPkfcs7pto6Bpeo23tyNnVIpFXqJC4Va+M5V6mhgEJzw
bpAiB2cWn8byVF8JREb7+Mt+W+v+KIu1xzD51lspirssIbVgEmv8X71R0UEzFQkB
XXqyndWmqAj3nybxp7WL7z+hl3Mm+pgmst5qPDDjDx/0OPATZuYobpx2/JGDKke/
G5UckgX1V9UKxPbe4yjmVDwaRehrmEC1LMYrj8Jgs5ZxFOqr6FwjqxXkwgwYaM3H
ARjcHDoKjd7r1P44zAvBf+ODQ2fAdivz/iHGpxbVhcVOtOLlUxAORfL2mKg75Zjw
J7XtSUMplJFg2psaxq7qKpyFmAmRWd4gsuF5qaoyQsoWmObgogjfkK3yHbDalZ3z
8+GFHBGqh4tFbk0vQQOKZotP4pxlilxdHcqted/O7kzt7LsS8GQSKaSMtG5XbESH
0sVvyuvAlKUTDSDIRqX4sMJMdA9UGVSb3vcWtVtYqqs2DBRWCQhp2pAgihWkLiN7
VcE771mK7DUS74n+6kQ/X4oiilX2kKBHP6hm5TsBioOR1MC6u3+bQ2gN6brohya7
SYzmmwRkqvWkx0T9jJWrnryLwjUHIAhSL32NwD1z+8wj/Dn+QRglfvP5wO/9vqP/
6H8j92fI9LBUKG6XmhCgnIuLf01P1j81fOeUkeuS9lD+wQssZo41fC1PbL3h0qVN
FKrzDxwXX8Z0tOelEGn4RQ3PB0JURO319EzKHm3IFr17o9oH1kvnl9AxEoa55owg
8Ig1z3nf44UynVzqVSqhitEp9XEDBnCmWrQ4gIv/KXMx8Ax5hOjkBMr1+1tM92WQ
hTBEwyMtv4P7dEIlPxLbk+KlCRzp1ihPUSPkANVGX0IFqmkijcZWS0M29o4U9mTO
cJbrca/F5ILgiTU/Fl8rcosRV6bqibj6UDqEz00C9mx4rrlm8/1NNo6xQpJ3yn+u
QU4vaNpuGUJal/a9iiYhGV7qM3nD1ARLxFlxkSfiXc0ld3Dk7xvbpDka6P1MZSUV
IlHw25wJeg9YR0ii/4nSE6aosKx+EmrSYzYIbZvw2C73li0PE3vBV57BaKdce1gW
L4PD53LQOdTzo/t8WEB1+dvSmSWVvbXbVt7zwCI4v/iiMaDr5i5QBQB9Yqtdh6iV
PDjBd/NclJbh7z6JIKh/TlSLcn6Dr/8jloO7QgrqR4L+sFLNsJgDNg7FDP39IIrJ
8OWa89P0q9dna1gQHC17+NV630UhyxybdFr/MBVYo6ham3mcSszBKi/X6RW52v6u
TE6AQ7AhUwAP9W4IDPj/SCnPF5wFkuK4sJgPbPMZm4XJ+pFqB1Pm6xSOhS9DHx43
FzBTPvVVIJSMdOMf8UI0Q6P+yaV8GH93VwgFG7+FQiTfxXDQVBfwaHY9kKUlGdGb
aqfZU2kyhBWhQEe7I9XiC0YqlqF5Js7hfiW5yv6wYKIFPgF0vIOQkvlXxTqEigmy
Bvxo/JVws2T/V24JchIxUqylWtnd9CZ3KcdiEKBjB41/ndVv7CCyiR+jnCtVUjA1
tOv3K5AVXKDb/X5WB+eepZ2aKLSVGy7bbYOVueWTqVAQO6Qtsy/EserMmEfaaZoP
yF7eMDcyiEreZEhcNApNVF6pnzdQo17qlZpkSqJ9grA9+5ktyRFXNS9SWDob0ICg
MIYMNw3YS22byYSjkHuaXI6j5qEVLFi86QAjNKeefk/E0VYEaydZ9B95BZghoY13
o72qdsnt02eqBbsD6rB2NLYlLP3r4hC8va63nWkSS8egQ9CPWfXGrBTL96shXRZC
70gURKCGNTW/KLdBR168+5SH31fQ5axIS7m8aIYYs5vw2luFLhgHk66zdCE+Dlaj
Au6DhKt5+DWR3hR7eZ33pxW6OFYM16LDEhbUfTJGPu91ZI/vJSayENVw66mFdeAI
EIzfCbV4SwZ/onhjMfUd8GKwnCrZww8Ln96nvRl9A3NdURb0paB68sZ4Sh0ighYD
gi0JKDrIZNl+mv1RdWJoBoHyhKrGDUg2TuZMQVCIMxSi5P+6//WAPisKh6bNR/sv
PJKnbJJrlyO1U6dXdr7mXlzMjM+FWZfq6aIb3LPprhiFf2qWje9UC18qQtDf3BuE
UdLvN2af8JQ3a8H5uu1TjI06AEXWFe+7WJXbmWUeFF0z0ViL3im0yZVivk37pfrY
P4XaAtQoWpBZ/9H22vEhq3oFjSuCTAcid8xU9FJ3y9SJ+DilEOU5tWmgRwXsKrlU
2rHgxerWsHBZvRiviu//0xa8EGVdDdsh6gHwNi/R2YoWNql/COiolYPrTLr8Y3ay
U5hSgUS2Tu6Iae8iHqhxW+heCi74bgpOXVeZJGGcMzRFS7sSIcMZyHWNOG4wOr8L
eeRwxwqi+Qzhub2ql6fjkp5JcUdqrflspHnHwAWURue5S8oOVZm575pYh1hkaLXA
1VUJ/jlVB/AK79wTtUCQ64TeLRq0pnpU79gyOD3vE4/YyG2e+JdFR35FdmAKa0mm
IYewIn8pCdEo+VM2fdFApJ6Cwy4vdUn3bz+BJSeuk5jscUncKXI8NskwWL0fx2Hf
xuzW1UtDf8fW8Gd9qbQFN8reoamn6lTOu8ldFMVIbRd8t+Og7yVXhIZXjEUdARXg
c41Q/Ar6onaLIytmv7AKGdeHHnVebsG6OZJJnLvKUEO1VHqitsoEOX3UyfUD+7fd
Uj4qaO3dXVNjag331FqcSH43OpUHJ38fOWcOTg8i0gy009JmBz+m5Avur+Asdkal
cTCd+A1HcmED3zucfry0UcbLQ/xQKgvKEXk0Xc55bv1b5DWSjrs3ekcs70Qd5UG7
WTKbOl0tRJ8r42s8ceqrDesIPd46jADi+9vaxhpOmOk9OR+xMdKGf/5wBec6jEPs
wSW8Sht+xEniINQiGi0+T3fzoCQuBVLsojD6oAHkgDt4Q+opcFvXmatXaO7uh58w
9qw+1/qGTG6hH/yfuU7hJ8sYiCez10toC7voxFCtA8LU3gz8cUgEbRMDGrMVPqkX
aXrDrU+es8hHV8ZMfBFq6aRxZxRHFjGhkis/8cE2fho82wajGq8PW58bxMMMvVcM
CGjPNdAjtCBmeBkQvHtKrB8jWYp0Fz8p/E41Fz6i639uDgYOuYHgBezdmsJKEDWE
mL0lDpbvPphvs2RXMIUJSYMvf0oDqBrllgwhdrRuzv69Ux8j/LOF3QO3/lcmInh9
nNB4xN9xLt7cjdPQwArxTdhr8tfG0osYgMJawpzrVKZhLFK5Ztgq7dKjK9oRR51C
1hO1Y2FGyV1ZNucg1XLPsY2h7WEnDojCORrbkEBvp1Nttqx///IZ7p2uV2jY4wAd
cIWPNTMTMHvpyJ3jDDdL/grr54g8xlkY8mBGxuicu9eB5ps8yu0Kp4Tv2slnO4EE
67rMNp11ylCM7x8hRUabuGpGl03koVARNtRcVolr1JEQZ5CrryDGuEYLsropCBSP
xdh3XU5AeVyfX7FhLkzo66HoGdpvUdkKAiCW51Jp1bkTwKTEmtHnEQznVMVU7fC9
rDsxsXPVR4t1Wp/dXovpGOdU/KEMFER982Lop3NLGp+OUitEP2R1ulT/jVgNDqZI
a4PsUeyJkz//BzijaKFm4XYFPeJqOJBdnLQrgwCF7J+OPYOY9wLW31CE/G5qyfKM
YCh6LZUixQJ4F5CdXOgLzPPPJk7IZ4Ts3E8klqJ7bEn6hQXJpOqxD7iyGjqlebBs
1G9PFctEh4XYw1n3uptceZkWzdhevIxFodgCI070GKG8RMjJJAByYuCwCyMVReIg
mgrOV2W4wFVvjckM/5pTUDH226qjsyqH5viawVMtp1cK6BaCHPADEmx8fWD5bY0t
uGnvuSLIU6auGkDc3Z91DJNl1Wbs29J3HiIOrE/7nbHhEW19OCNOZ50FuKt9Z02G
JLL9uqXuZGd6hUktgcJcKcwDvSI4RQH8FLxvGRW5A7PrYi503i2VjjPSBiCAL/8q
xeQb0XuTeZ5it4iWPAoH+0hxD3KF7uStYYcohELJkVb0DG91OSX8XF39w2kIaMev
jYUaoWEL1HsL5DwYQjWM2vaV2FJejpqcmCkKTv+q48+wyjytq5ObZw5k5gIqbLNM
NwQGCWL0GENt38lsRZw3diVbKgyDPuWGXnl6sdrF16q9pjRK6NE/1VcyB877tOZH
FLYyNWvrTLd9NUlNSuJKXO1kpNAsNe0tXQg9CDzbkv6V46xMw7zwFPvHWX5GB4qn
0BWPSmWkAjuWKpOqsFBIEF/lx28DaXEkgRVscV0tABJIKbWvgNXXbD6gF5iMjQMK
d5Uqb0f3w1rltCZTVUTcyACbk/ypU8qCF5Es9i1jaVsLahsKb2sgDzahIv+Pfjzk
Tb5UVAJllKTD34gZsvzTPj5aC+AjcvXK63JToiVHqHYB4t5miXmKElxcndOBmBfM
1jSmuQXnq+zZKnEbTtih4Xi5dy0Hb+iw+IdMkPihOrpeNB8cECtK50k8FTQQiIHv
tXTQlv1150MeRw4PKV+i1BsHSpd8FCHflu0wqAtV9lCTJ9NgLiJxFbJcbeRTqppk
OIYQsgCJ5c/uFaYSvivF4AmkoQmQ29jHdV7pru+b9OTCa7C4BeBx5DjpxX+kz49+
a1jFlJGBvvSceA3vMo3tSCiqQZOmotq4vdgYiqyT6TT5AbxgGfCMDNrMypRT02mt
qB7X3xJD2oAtXHgW1jV+INPnTqiAavNLa2U0MRiFDUXJoL0wBojqgYtwIhXzu/n2
+sKuA2Tc3ZXTHoyaqL1+943TAe4AGjkXQgSBl+xSZtfw4dnHzKT5EOxBuWI06JrH
/kLPKzetomOUcQFKs20+8dKev2m6Bg3PrpONLSAVnQ4oEzbVNr4aFm08WIBllzJl
3X7HxpKGabjSvMZrordioDZTDiR9b4DjltRXXoNk8VPeqH55zUxmSiS9eXxn8QJj
1axqA+xTNfvk08bfQ5asnsPhp2T6+x8BKuY/P5QsxqXCsxzdpu8fm94No5eia8B8
BU2HPeSw5VPQIpJxYZdxMu5GuxBB7kkKf7hm/BL58FZcaj2vgQcL3hWF7KTolrWq
1lUV3qzkApl+FwnPfqr2J6ObjcIDSE4DiGv6E6Gl+MQgmfgxh3w9SGTseJ/efwhc
7ZzplbSPW+nFVp0XmlIkcgmLcZHA9Ko/0Ulyx7OnaVu8jfDb9apig4aJ93cR9jNQ
3Fa/Yv/QyQ3tbJyi6zRHz+uhIUh868qSTv4ZjEK/NrP/b7w6qpvDTflOEexQ9k51
74tjST0AazB7T5umJNHFKwUw2j8RsoC8HS+PUcChGHV8G+J5ijjihPahkgClQ0Ru
xKKM/si7fQ9gBkbUy1DNJQca+dBu3uTF7gnfRP/nzQdzUKAc7Wb40gPOh1VA9Nt5
Cm4DuMrgBqNGbqRTOlfAmJj0WjSjvXaVwlHko9PpyFIrA0PHQGOVMl2DHPnpp4Sn
UEI3ML97XfPHbJ1Q4KpcmlNNBH/g4wvBTjnF3wHyE2g2WiL/0L4OiHm2z6Ey2x67
SsFo1TqPSf9X8BSVMthE2CibKO3RlgptVCd9UYXME+3ZacwparaZ7COY0MaXF5h4
hLkmlY1Aua1qGOFGtdGDlbgDDnsLEEIZNJeIa2WWYjxBuKvyBExmZWyzCrM0ycMx
HqKey886eWfY5CEg9vJNrfotgfQM/Og+8YNU8MdSIAN/+28ykFIDHkrdh96XyN1z
IMSpawvoAJdcxXCb3TN8dGCEPWmk2whgQHmYVX0x+hzXEowVxDFvXN6SiSUTB4Wf
ZbE7r6x4ieQPR/Va9BGL3mjuNdq42nU+sI1TdnwuRRSCS0Ky0EEs/KhfjWRwbFMu
ZvEgBogxPpqQQcA065vgPtacvT0AcRZb9WX1NqEw0UmECk7EFKGe2hmQzo4DNGdA
rYnaZD3afEg7Mk1g7mB5KZK2bsMO0L11vjuelSqFDG6sMZtMxz39XrWCnOE93b2E
bz9iebenc2tsYwStXPYiBt2yG+c0WwL5P9qfrvj/cM2l0oTYZ9bpfbrbHDN5FgWr
UoFsfgZdTfyfUTjXDJjBmE3u0LvmUCf3MXsFAxnyYLon5W9hNht7YdBWxL7+m8Zp
eeOjCZ1g6yLUo4sEKQ/1+PSt5gFgKo5BIJRdniSjaj5yKLZjA4VwcId4hnYQPBwo
K1epwc6Jzo3esJ+/TSX66mRlwZ6YATiEyVkQtZAps1J8tx9gNkj9t9zfagLRZ/C0
PTW4fa+YK8RJwdxyv17qe6d4b4pxGKIzoGKmD0IELKBEgW8DLU23aI/l5w0MdcVm
HZTg0SssuelvjuIHusIcB9nORbr+lXw34/GN2YNiwlPdmUCXLz3lLy+5a+OLNZi9
Z4/FmDLnMgDH0wMe+TjotIsT8gW4dq+l7vG58ro05CLud6b/KKdh3AIWk0V5Q9Xo
asVGJRqLTRP/I4OdyAll4UNwsVJKpyUbsTlnb90oKk1c/tg5YOkG/Ya00yuBrRGE
ZmijOG1/10RpCVU5+bihlIyW623mMR9IkvHrgUDiaQdujW/QpNCpazX5/JQtEl6c
Cr3tGERU5tUDFMEh7oXSVWpdFSweCaW/sx0aL04XzIvynzTgDfQL3SVhwYY6hvY0
PqMYhuPxGgsNHVKdlyKprpfsKNmO9y5uFKhr66lnRhvq/JdE53JgwxFfNbWCP4Pn
9bRHkFNzp+Hu38B4Aw0WHPeVLWwDm4KjezSNcFkfeVIzcd1sFGLOMuRDGGIY1G0X
ReWEaD023wIMrAMuoNY07+Ypl63e6XbMdrUmIiOIzV+I4d/rttkLFGdd3l9N0g8/
rebt3SGni8JeJ7gYZXegQHu4HmuzvX7DU1Bo2GZ9zZkVmcu3IUSshl+uL/UUYn//
H0XTF1jrv6aT9mUfgyKjCZsbezVLtDSh3zpF3K2E5rKmJcOAxojPajLJbLfskgnG
xEw7KGz1+7k08k7FWjeDlqIAkfhezpCEYC9G1dCXwWEKjXMtZEtGzDBphfcsqGHd
tgaMz+G2aUDe5SEqq6Sitwm/ulbpNDM0wFI4cC3ueU9iEah37OvMXlTsoVI3k1FE
QBxYq+HKcF9UnhR/D0IYYm3LEjo4TWrfFqSYxFnHDxexYWqep0ZqHl0fOaxoEtjd
r9EKfcIZJmhep6I9BayFzPxD/hlNWl1I1JBKu2iyTOkknfKYKLYRY2rr2BmP49kz
swHRwmn/DQH+vvJ+4nRpRnV8OKpGUZi3dcp9EXxUvSGpW88jjd08/SAgnf1DyQrA
+Vg45nWX+/IfpLbfeYWeK1jeO349eqcZvePP7+CPs5pATT0NE7fnQcILKMvQY6ZZ
Y7jb1o2pMSKqPmLPqIaBh2Ij5mP1zGproDYhex0X6oQxXeaV8Ncmf5Go+fvS0rbc
oy/lTWlYMsFuZgGbyINVvU+yIIR7q07RSjBw1NySJEa29I2VdS0UZ7Zgr2xuWONI
wg+CL1MABXYI3zZOV1ZnM3YN6CaMg54jBRsTUoti7TnnffAvjt4OQau809g4YRGE
ytw+Os/+8VL1+G7RQHpzTotr6gMFEXUciIfuRvFv42SCrSyO2rTvZsSaak3F3D59
ZGNPW/Cr8+s34BAfGM/k+KLAlr8dVSvVsUcexrSCEil5g1HFz3V1mpR8NBFGABob
j+JkZ+UmMYWSt8XoNpH0CpzVlOC1+s8plo10ahwv/4iOpor1ehohXmxYtOTcaOzF
16rGwWgGnjdiTJ9KrfwHKeGrkJGBCaXxPP5crXULktmsM72//GN7iWGOBNQoiGac
w/8Tii6hdEoRnrqBcxbtSpJY9UmmU2Q2PbzCsFFWU5LfHP38cIFHuNCt6Fn6HZgQ
GCMDT8LsfvS6pzaKpxtReKylWuTc9Ss4WbSnyMOrLDagJe4ms9hwQzmK0MTxHSX1
mJaYg10s6gmYQVSv82rbKLcM+BQfbedBeMFtoMxhBCTjX3CeOd2XsvmntEqrPG0/
rpGksaSSqPX14zrbkEY5+UP9TsrVdcjxd5iOJm/xf4++xo1zBeTTpoafQgNoxGje
Jc2tXVb/unUMcPAS1x1WSXg+QqfZjQiDOIijUoQzCecnV00nXsnhbpLz9RplnO3R
ftVwgADaZcKuRO2o+vuBKVAsm7tRrv5L+SjmMWcFskuKRe4Uwea/x5bUnXRH7IK1
9cR9eKwmi6r1gsjw67+1sjLwwmh9PXdFQc4fpx5rSdZGoCh+wgtCGBOF+83PLvp+
wvKa4Eop74YAlaAz0xJ21Y8Q1ExN4+kZT8aP+Y3C7muEkFQ4iz953UVx+tVi2uYo
nmRTETraTAEXvwA2yvHph5Gb7vFyswaGmu9WiMvN9vAFxezEgUAcqDxEz7cZg/oR
DrseBwjXnACVoguC1CIrpwnsPnQe6y8yObp1r451m3q059lKqXfOiWhrHhF6FVab
aZUOKVmUAhXAPPtdXI52CguC3MIiSgOXUcHTPHulaNlEwLkJBMepjTXBuQ6Wsu6y
wzOYiSuX2HxiknmwLG8k+gT8ijqlitHpTKGyZanN8idNw/bwmVNdFgVCqI0Aueb+
hlh3qr2R5BbWH2xoX2CDrCasEkkqFZhnCp0rIKQjGs2fy4hWlfi1qCUO3JICWOQm
aMNjQRGxEP9Xw6wD1rELrVJA/cxOlr5ylHhe3qaJ8Kg7qoq2oLPqDZ+r+9HJFEeS
yH5dhODcnHsTOCW001b7H7HhYM0ruHG6iETc2ZAqEosHVjlvWFvfS9tCvY92bZK+
uaoOhOWeZq9R+c/RT4GJ7EzaNB7zmKdkP2JYNhJvat0U0uFtlIJl6BT/phUcdzK8
zuYZTtVuBe7YFsO0MU9Ksb9ANE/5k7GGWvBWc5wn1kDqkiX6/CW4O+CawhmNFx/f
5YoenQZEv++v3egYR6Bzl98Txk/lMkBBUPT+vW/iIUPGX+OLYRL0wSwjiGlIH/xm
X8jhyxC3Nfb08AO+TvYPon+GKBM9wPruqylZKu5gPzoB13HBfLD7EHSBcOaTkJre
B66HG75co+WRANjRqtEqUo2U2nJ8dkgxvrwIJvvwhpM9CVWMBSD/WVFt50X0eZ3F
s4VEwraLF3T3oiwms4J1HT68maPS6VfwVMYSJnTCbngabY2ZfRSdXDSGiOzHH5hS
Mlr2JMFCUIGFAKCul3zdRkGWT7C191bx+DhDmyJL5T1B9yEScNCIQGjIS8brLOfs
y5IlgBoiwjf0FsrSleAyxCGWRajlbBPXNj36R3qkQbbpXforDxV9RuDKBo91Hd3F
iE/1sVp+MPrD+SWmW/SnzzIGnccJ3PFc9ONwY0k3k/MEWS5imoNRZVO2RC1zLW1D
Jr4g5PLxj2GTbZBDytUYFqAwvgnN+lyBFz2AAo1zgQGKIQMFpQQ00Cm2Nwn/XOGN
zT4bCIjghlvFO/O/buZpFja+N0LI70ypgRQEDelOi+nZAIcdN2kviU6JijLQbPSu
0f573HvAtKJsDJC+EnOsY+1vKXPfKbvy6xkuGuseD8/ET3q2PayIHI6aXPiw9Yo/
EcSmcMVF4IGQElSD2Afjh+QUf0H4S9f103PD1RuO/X3F0hjkBHnW1oQn6WoHkzaf
yNHECcQy0SG4KVpxRRZ+xvHWBlOeiSYVvsHvjjmOUxHmfv/wZh8aqhnrcbLzcVVN
zoifh8LmjChX6uRozwiFyF3cXwcayJ7VdAg9nWzkpTTg0bwPS5Ooutb0J7ZY+Qld
kki4nXUS8OSqbodW1Yi/l+p9sbti1L2czyXKtYnRAsDTTQPB26spozUxGSVxm5r3
Z1/Ik3fepodpvkD+lbXUZSHBazIs/+aE5foDcmPUJRoyVkopd0s5i7ClP+lTYfaR
VFUQhSTJbR4/oo+waax5MWraU/yWbgYlWvK4gXOAJMiW1sACYqpj3TmOqGHh2BJK
OCO2GZdhrCq+oPQcZW+eBNJuFcgoFGFr7BbVVqzd1LkehvBDB2JG3R9qO5dgOONN
DdpmB1DPt/R3Dze2YLYuDHEjB53ImQVs6A0l7+TtqogG+83+Y+UGcXpYXjZapJ4a
nMYaQDtLugRIfL03SEGpB77T2xUgZ3PPYKdsOnNztxbvnjv3kNpSgm78keKp0XrT
krzelFyWA19kwRZjRFJpSt+3DFEEBAjQ8QRWuzSSXjs+b5YMhSwSLqPDiwelw3EN
lRdu6WKfHuC6jw/3qqDGh1z0mhZJY+CYOsqicljBwyCT8JdrSnJ/BqpEGDLG+3X7
6D60kmCDk502myFJvQpAXWqhg3ehM01TjcXpj75xxr8ODgAXnrVf8b/kcpCAmY7H
ElvnT8S5xqf/rmc7adtYJRba7CFVul64y+ZXu8WEPswFiVR0Si6hYdIvJWWHWUnj
MOUe1rR5WiCzba/AVYJBPjd1JFAVfW1gUZCPQyitS39yp87jDbmWSWD15MNVxd1F
byX/CfC2V8jIeYvyRW7OIFUh2VwNPqb/0kJ+NxwpTI7S9Ob1bmvfj8az7x5nVAqK
094kjfuTv5nCX+bzKDxBP3mvJ1W4MsVAA3nAuP5TSsYEJn39kTfAkf39eEiSfRSA
N2ScelpLYVztBFaxmQU6J+2+gM6fjQw23xV16aXW9Oya/IC/uKNNQREwrx/6GBy2
4YEBGSR9Nmz019HAl5G5nxkP2QSyvt0m1KD10W+p7QcnLbu+3HM3BVvDhul/jPLR
AELIN7GH59sUQBlAllRGN1z/U4YlY1LoG545b5EJ1TocnbKEbOKVP+LqlhABaK0z
SF31qNxUpyArjnQqLZ8mvWbrSVcQTVhU9fycBaT9+rsRtaLqBYrMygvC1/O5yHt8
GpNDJszi3M2ufAb/tPj4pbSQ2bJ1KHLF2jsLhqChnZOHtYIR5GFKGb7MQhd4fSIb
j6dRKVzmdhQd9A2FF3Eq3kdzagP6AVAR5nC9Zs7R2BmokI0zngwV8iu84gvztGEi
H+ixLGShA4OLABvIgMm7GGXFrLPrHnDk8TV+RWqcihbtJi86kqB48TtfVLug5bvl
TEX5tHigrjUZgTEHvSq1SGvnr+Gj8TPsCaZ/ytjlXsrS6v30G76wKYYF/XOJYQg0
1jJao9zGujgTNLK+O58uDed++iT5Df11DKMJ4t4IzX7eAZD1MaQetsufIpm3kHMR
HjdiTeiKyafZNcokmXohdDwR7fasLfCyUX6ffLQdFW8jBlrz91wv5eF5wigAKSfh
tmE84cV4B+msdzvrqx9OMfMD/tiY9xeXHwqiD9zNsvFTDJ4BHogA5PAx3mCdNUne
Bz5o4fmhXe9sc89LsP7bKJTI6nTpW7r3zI4cgtTdAprtFaZIhqZv/fVby21YZMi1
zBDtu6ru9Y9SvwITTmKwS6g5fJJKhlQQjd+z06Q4SwL0JYuos0bL7oj3KC79orfA
ipBOjbnTJwPs+mZ7Wc48zLHkxk7/Nadzq8za8OgUuuglRF2f6B0xgoJmqpO67AV1
vIbsACHvYrb0PKOugIFCPUHKeUsqeV0TqU5YtnmvdXT1O2BTWBOeTPXibcvwVE6v
HMaORGDCPjvSaP9ewaXIsA8f9saYf9GIJ6R6jQJWWpCRKqHN4QyPi/Qu1mJJnuXz
DsGgjrjzWVyFMakB31+6MYv/A5aokCscVbJZjNEwFMeLfzAp6YpT7EDZH8L+UQvH
SY8Wv1VO2cL7Fbr1yAgIGBra5XT6pHgAGzc93IAMxvZlDdOBXp7j5MojmXDincdE
uU/rqOB7gQLHRo99iWH2c5a62waDM+cS/XnsbzaMwVr4qpA+eMqPc1ijJTb/oy0o
cTA/GI23WhEV25lk9uQjQjxCNQo595eZAY4UtsCN7KJTYFZ8YQFN0T8DDA1b5JM+
SJst0/vjeo7JS1jJDDBEuLVy7BCl1WZXn+DmuhtdESPtIQNishn8rYqu6PVtw9o2
/O5gI5T84VFS/TcsE4+0MV4Q4O5Z3f4no5G0/SjH27Vtwo6u+krExnKUzLGmI7LH
MZwtRxI+1o7fXugX02YrvFVAYZpr2G0o4nCsZo+7hDmg6L3sDJIe8SrQGgaL2Fhy
C6A4B9fjAFHXu54fKA26Vx6zDS5Z8QjOUW/MFh+p4qVYaaqKZqLAL6hWfyoZB1kl
UaTi6MKrJSStpU/TumZmUrj/E5yuafUwjc/pBSrB1cQ8c1KasyH77jle24TCmRzC
h3R1ONmSXITd5SfuWef7rOfeFjaxwrrjNGu8VIACuk5AjJ6UAYePpwxZ45vv1ec4
P7dr57TaHMirkdGDzx0vEvu256Vv3IYbqk7DmOnrRmhSTg8vEbipsGNye4eAz9hU
/8LU9EpqSTqSKc0OfiBgemcWAKWTymd/KszSCTtSkpP32JiR0a6U/ui9EB7tPz97
cthHjKDxPEA3PMyFCMVqRny4j0z3JSR/Tdq58Bb50o80DY/MYbWawu1qihafmcAN
wrhnRyPDrARSTsnQxEa1RKTm94P/mM2tqfvVrdZxY5DuzSyFZgZMfL0e1DEFKZlS
xFDqcPzpLjtEkd3oM8MvRrrINm1l4deMLYhPj51QK17CQjbCzPXW3a5qBqwMF+0X
jeQ0RHeHx1LqyR9PueUFPme2CaLKItDMO1CUrw3Uif+GwcDOZnvbAkTTQSy700lA
bOfLunk2nDo+EshHHIkVJqRDm/8cve379diQZ1CBRzUHZSY7B/xyLCgvfshCehOm
cAEbSESw6qmsBKE1wFasAhvvwaHk4RrLU4YO6pUHjp0XEyZpmF3I/Lt7VCSqFHOY
EX7U7SUSCPB41YqEDBGGcf2pHM/jl3yymGQKVQD1DuOSxPeYgUHkPP0lJbzexA/p
2nAf0pZWL0pVixmdVAaSLlSURZgHABJxhZrra0jpGaV/7rLnEeIs/UUQkYGQ1U84
69U2ogBmSc+/NADQutb9glaC1trq+Gi9jdigZ+rnTA+kDr0bdmkfq33dEkFSnOMT
1YfgLbW7DG4U+xZY1Da0U0dExM4rxApqLFgbl5yXVtEQUdjrGxkkZQonjJiyuGxL
1AcGoxemJe2WZtrkNm9R+z1EkKwrc2YDQWB3wCnGYhnNoQwqLNVa80onCNadGw9T
f72hqDgXrtI6Xkidge5o5+YzGpk5A5ODDN/Jx4jxB708GaCUvJym1qN0L7bH8Sod
DkwMrNl9mciuL7GwKSIOe6znJJkWowovizdIijp3GnGd91TfEiioT+6ZJ0DVZVZN
wrxz7hDzrucMvmQi5sniTJ9EUQJ7EAWU+UgCod1h4xarKf1CDLfvEiTRshT/Qtwq
8kc0VPxI19pc+jMwsZJR571iRn3mFy/bvqJG9c02keDic0imj2erTFgcSAB9Pqa7
tg8SFnOc561hLN9WLqBXLEvg4IF7I3JdbtMImInSkiBs31/sfGhXbgUnojEzQnAq
NDJuZWm+apV1abEuequgv4/zjkREBaUury9y05VBPg8zuMDUPl//yYH3IW043/D2
Z9NwKEXrTEbzXhW4za8+z6/ubI0kt6blDPPa27MuqEdOv8864nGQzwureGYitNJv
Nf/381nCt1V/59v5kZeqLae/dregoeNA3Jo8olN+SS4bC0hBzdLN2tx+1HGhdeFb
mGCI0e0/zGinhs5AWVatzuOACyo+/jbw4IvunctNaRkCnoBrjV5kKcPa1q7kez6A
kWq6BUh0LYfBOpUeHjskvR7XvzCCPWkcqGoDbPZMRWu8CVCOdLlBxGzgzQnKticy
g0DLrLY8a8A3bjjkK3Q27PMekTjEivJPE+7qHOhcIsU34C0sWWRjL6mnaDX0hvAk
XMgkIsJx/h4PxuNtJ4byjqkFkAKVWvOSksqBPCbl9LjzJOwzt1K76P70bADfgL8v
JQpejjmp9hQyInLwh5TIbK4JuFY+i2RA8RaJLNCtvKtsGG+JYVtvhWgJLsdJNSlU
8Hm7mrWBKxcylqRKN+f0XIeDQs1NR1Tvwke8r8/b0vnK2dB+00e4uqanDLroZSQQ
Ea5cgfAkkAKYH2ZoA8gesRuVsqMG5tbkr5JsSlXTldnWLiJHy6qxwYHHtqACxpWi
5Jc1Y0RUOuRsAGpnfgugk/DhUo/zcMvLmQHqLDm8MctyviCiSKF2n9Hq5FFJ8MG2
teS3paJMbwfOUuvEoXyr9VENd3QailKDIC4Lqpojy6MHrFJ7wMoPo+dEs64LT2ux
YfJLXWItIus8d4Cdx6ZcsKP85BPf1b9u2TZuk81VfzxCmD21U8vGlE4pkSfiDth7
5qE3pc7Wv/9qNOZK6UfNixD/Ith/6j5g9DDs0CbyYY08FTmcTXX6kuEZoTBoOWX/
/jylijr1sc2rC9jolIy6ccwlvDPdw1/wrhioyRwxxEPqImbHmh2QVYlRoSSypzbt
Q4NOU/HeNtQXDMBOawNIiMKqbSXTMk4bk/I51GK7o6ezPWEx6ekiwJpFnA+BrF7p
aUvA4cfcSIsQRrTZzQuqA2/1cJD+3Lkz98/RLg9hjUvo2t2bpjcy6HsFa5CP14tg
WvdXuiYoGYxxJiBLNS6RU0sphmj740MTjmF6yq0Tt49BTZfdrMTzEKjLHwjKPjnd
xRprYwXczw7sP7ILyfaXrOlr9c9qt/n3dixTKaVMv0Xj+94C0flQmrqv1qN2aBCH
qvY9V8yIgDWIxtFKLK/0Lz9TQipNGIMiEiBhGBZo0UjZqJkWtbu2hUAKP+PT/AQB
wqwZn1eMIIBdx6oUE/Y1tF4EB2d2DdcNeaEzwDOlFEabRa4mEiyfZCn6QRaCxw2H
XIb5dnzkNDWHFjMMqmT6xl0t8BihMt3bLcuRGIivJO3bJYyw850HqNBEdY7h+gW7
T8YJ71LbabhcSjIWi87AmmrIk87vmIqgSgJW8WFGOYte+v6kwi50/lm/hHZjFy4R
X1KAlx5d3XkhD6y1FyYRiy1H5jqyR//tsmOR39saqZJoWBDGDcbV6YppxZca/Z3J
LCcYVe9QxIgQAy6izd1mKX+zTXF9vc7TdbIEqznqSTOUMWcSfunBCIsRGevkbUXa
oE6FHxIMusNY41Y1z/NEbWM56mHV8EjAMab1iJ5FhJJllokgyw0ZTSeTJblJxNsG
xmv3V5hfOZi2V93R1XxFo0DzquHMMJxyIAyNuLXITXtz+VJKT1N0esyUo72AHm/g
QLD/fNAK1SFHPO3owDVpWACoYeTjTkY9CYKdxUymbKhGJygLKZM5wc7FSdGA66Li
VDrN77Qd8HNgaS9KuTVJ5HngYDcD7xkehInKLYHMYlQ0mUhsUUL+si1TaoqTc5xG
Hs91DsQVGMAH2XaxhviwPxb94W4K1L/grR9WtQZJxU6jW/zSWr8g2gtYiCVHqO/G
l/PQpU4t1eTsfeuGFvdm302VhnhAPi72WzHQvBtly2aZcSxkJtF3OCfxPyTUyoq3
uhFDURSicBBIlnrPnuUsFoxoaFSh0lu/pv4CVhvv3pSHI8K7t0jtr+e8yFwJ+R77
mJA7w6RsnQVg68rTwhk4/j6B9Q4P2qXbO15CeNdV1E9k2YPWWDXpVLXYXyw2+Jxv
Tn+Wr18l8lqY/DlJBGE4XXFBG5lYk6uGGOBhsZDTf/gketmkOJzCXUKYhGZbR39o
E/3/YepFGwFoNf4ME+JhpmFXk9/UaHPe0rKqw8cSDO8O2z88ruIGsVs4onEYhz9/
iPPuwPtARJbjTGEUIYFJtJI3WUkUeMov3vCXqk7ez+W1jBNzoREHBohE/dc5JLFr
rim6vSOhbbtsaTLszHq5w0ZnddOY2RVjQWbMGGIDDcg6jl8j4ViJxvkc+8SZwiXy
8hfSwwwjSmHOojBwnJGFfe/phRI8s4qinBjTtiOmyBawav6yElqaIo7RtGNtpQYS
A6SZVnrZOyH+X4hkYTr63AC7kexDz2LdxacOIFRGQ5xpQZIYceuZwg0TKKB2Iehp
bvqcQtW8XwzsGCSCMgS78axbr6eZGffKwSIvvbDhTwtsajmfvo985MlB1uoxYIaE
9L/aJDKBi4iq4oDPF4F6aD0vDbakuBs2HkXr+gHNbL96DH1+zU1ZU/PUeWxAu31X
bmTndFr99tUJQqtLnVI6iMADbcHJUfu6BjHeJKDmBOtRrCyBddyGjnTnJNpM4dgT
3WC+Cyh6XTECxw2Ys7r7SWfnUXbK6j1zoBcEmCdjyWa8bEK09ONl3kIogyaQP1m5
WD9id29kpDas+PZokrJKJT4XuIBZY2+cyFwV7jTtiuMjAqJGEQA56goPDf3RxPPE
USi0DhRqvGVMfk7usR41DERTieMdfRD4YunkKJOou/pKoEm3Th2TKB8vIX+EPACH
EAw4kABn3iVslpReLZRmMiqByiD5GjuWcwvqvBM0rciQgqsBfpm3V6Duah8TZKOf
CjTefcay1XQb9OZ2McpbzetAFk77g1E/PJOoc2dZF/vno1iKjqSRQdfmDpheWvpW
XPqkfp7sU+KO3C5y+KtKJutUeckxCQFQh64zIxD6rYSxr4xXnXTa0vidOontXsj7
/uUi5Z+Ix18TZx0K1t9t+XWImcHOKlOwVKcBbzHetporJxThe8JygSNAGvsYFA8a
AQxmuJUy/4gWtEOgqeNt8lLUpJ5Y1t3ugPdNw2czUJX5whtD65BoALNHu2V7px4X
eZSkROxdtuyHGnX6e/J6UWmCVhZJ31CVhxl4goq4YqEKIfrJGrDbgVhhIoKCgY15
S3Fl5BalICeV983hkO/+/x2hxEsuiwh3Pr8u13Vjo/6rAUwSVaTj20Hgi7WGgHbH
SRWzn6opsjlTlLLci/2nlIiPxAL7DoVTRhsTQbhMWtTKumfkx1FXCr/IaUShwU9g
ghh/HPx3eNXXJKUNf3ZOj62XPNlOdWUwcZ2ZvJpjQDhPdLKcjp01DgyfHgz+SiYG
pNvvFU7T5p4iixDi1keirpIbt1OG5r3wEjQmPFz2B6VL+m+AaeTOvRndufkcaQgv
fLubyTC1NHU0vm32uGTwfagUMCEHWigeCF2gM4UZQPY/SUAF8dlMZyZk9TWAeyRQ
LSYAzTfIP9zaRvcoX329umnrpSa8NlQg4/d/CtrXU06r4l1R5jLNtzD6iDUMINF2
2UCAOui0jrIDL+ktfLRe7dVw1fFemgu/0phjrkhlp35J9RQiCPIkwlRgGygvUQ4G
76S2zFcw1+CjIXOdfpSqLaR2XhGi2UbmuUsp+y0Qciff6bD8Yl3klLyXTONLvDKQ
siW74VM41D66PS8M39SmFHevqz32Zf6p3OWFAjnXqH885ybg225+Ewx047XEUa9P
UcKwl24rBFP73L0CrTa425t2Poc3YodqrRFlKhPuPemmZD3N3dl+kmbJ8HbIEWCT
0mPi2kEeE8sNTeG5tzlJe/VNbih04sYDLIFcuLaZlajUn7oKpTf2pPOtsdaphVcL
5o2TvFGdenz2Z+R/X36dNhkxItFpOQVeyb2D8z4JoCoMQrfRq5PKqUdyV3xXD4x0
03Z3Y1X8Zr662bLHegxncL+VnBpq9gNjegVgVYMoiU5kSSQAVC3LqJXHxFMNmb5G
myFf+aLUlirbTWQTbEq1Q70Ow/Uf9BlgKnI1DpaWepZbH2zhOvsevpkuWzJaDs+E
NtU9BzKUWWnJu3tGRMFNRV2DDB6CrqkIBxcNkqisHAJdJGsFrYJ8w/0o3ZbkGfcB
uVwiWSG3LYFSvKiK02ETofY+QHtVhfeKgecpkhrPY8pvSoOclBbvemgueBD5HSUN
OUAeE3RWoO7+O5BMUWQiEv8mzqYd1Hx0ebeY9VgB4yfHu1PBU6M5GwoCuBTR7s1m
Wn7L+4HbGg/JEAf5ULb1nVzBbu46dp2UDxlPA4rq4LBAkmyaZeW2yo78dxhn+UBC
/PJaVtLAfw7nOMRPYE/FLYP0g1WsNnb+/n9n6VQnBfIM4Krhm7Aek7ZEUP2v4dat
wkSkVK/1jQ2L7aMp+ANieNsyrd+FfSrVSJ21S99fjXF9KK0OT/17G4QsKbuFFQnE
IVYSCaerUA0/HbrZBOi9zxG7EJVknG5vn1vTrdFMkbFJJaSf/ZK33V3aaJXUThYc
8zrrCATL6suowpj1VQVoxYnWx/gRM9mdM4d2YXzfzIEcTdgOG4O1/WBO6W+SzUBv
SPSIkBFx19g81OsAnfDuOo+DFIM2iTxPBtyKnNqrCFA1CMKj4NUf7M2NncqUB0YL
Ufw7+4cKNWTvhjuPVUwZ3UPNfJiRLbp2KtZZseJ5Hc8RYydHeeDPLSFfwWvBm+v1
zERAnBQ/OEIk+UQSwWDTusoAD+ErbMpv05j7fWO8oSL5qFg/Qxk2LLV0NS4KW4s7
Cwv7Tbw2Q80O9mASxFoxSi3GDKXnwMHY6kpuMFoF8Oe63GQsOJyWOBW++ldHo+kf
S73gvu1CqbowbZ68ADRQllS9Tt0DN+e9mu8l1OGdBy2eNvhmLp+vA9opDp07sPtO
wvPzDHyVuTUp7J9ruLt+6KmxgVcFz+PxXTFCIUMOlhvO9SIeGYY5b0AgNt4d0pC8
pGRb0i5cDVMs+5DjDf2xQy6/fWJYZHReM8fHD7yYJKqSof1FEPje+Gb0qXgVvuWR
O7HEjUuj+shHl52Zm9suYN12mRRvZmQlTzmZzO6wQbpjedT/BbKFVR5ZzDkQMbQn
qwpfP9QZgmgT7JhJWqis+ioc0WcgtsnskHo3FVBkF+OYjv04b5p6SeUvszgR893h
xVizBJpzu2zmAUWyYrOATTiVvqyzXTvwOXEeRIRPEFyxkqsHzHSn4XAfRo+mGDfe
bXyIDzDvIIVRF/Xm2daVt2i6iO3U+WAoiMN/6W4h5+ZQlxJUbr3UBfzI2H57YHgs
BwrCUs3LaR67fMIsv//UKuLvxg+9+y8wKYu115aNqm6j439PCvPY35NvclmlQSUf
mTMX7E/PeUxVh8UYJcT7wG7QBedp2kFZ6PkOYD2Gqvf36/Qi3ybAFs9LgwFq9vRU
b99hRUm5x/LZ1Jc0knF4iF9yJ6XJKivMTcUsFvMiVCRrAsjJqmYDBvpeHqMiw+iS
rZRDdHIsO8TfLCRMgC/SpUTXv3vFJEy5XFq2Fad0blHTBTJce7Y/SIvT8dE3NM6r
yhv9PqXzPqmOSbtBNyJfeWlpxYXFo4bkq/aK9BbjKic4FxaVJv8GFWEJLMjidMY9
bk4jWjM5vO7alGdqazdAd9dNgTUamSF4eoXqsycomn1pkSHQHLqPCgjn44eYJi+d
MxcEIK2EEg6BXWZUkV3+INY/mZcM8snfyB9UbfL5iDnoAyTl5xci/jqE2XxLkP/m
oM3zhHIdGt8YHdiEAxp38CrlgiDsLsuHMFlWXuuQ+Cse+LzBkGC1sEWChIBto5MX
j19rbyo7AZup9/lfA1j8mD/0H1e8meEwohI9nVz6HzJc2yiiYO3tiYO/ZKNmrypd
Tss2CGBV4D1/eWbgquEsTaffzce8oh+tx3Vb9qXZDwbNX+GAcJYlSEkkbwNFekEY
Zk8oj7e7T8ykBcYJO3n+8f2Nv/dqZeGTS6od8bEuiyv6ljtCllyUWOlKu6BTfHyW
Znb9Ix/vddnrKKfnDThbbyIWqmzywBrDE04xW+pyLyoZ0JsNSYG+6RxRWU9xuoQE
JcrPDj3u2uTDKs3929zlHsnGFN10bPLmX4Dm4Qx4Kiq4s/VzudzX0zs6mVxKy7d8
BvRmAONKfGHGrT6GZAh3WjrEYlNTuNM7KLiUPD+UF0xV6VoSmW2/lkXNsoWEPCFn
qonvvR12h9pSyl5XYmG/3jJrHEIJdd3HcCeZj/FrhC2yqleyoSlm3EsuJ23KmONA
IsWcIKrYqFhO9uNT5wS2AXTDNPy61gizo965oa1qAzzYSDfs9aMIU0Mmp/R8LD0q
dfhjuaZ31C5PP4cKVbIEVZhkRd33bHdp44HsZD/8RCBycov/xLzjPUNhnGoYNkkp
ATdfyxhRv8OTjckRo9sx9skNjpcGcT/0nzAT+JYb87uBuqc7OiL92ia/09fUF7WC
0N6yVHwbYX4Cn93es/J+BPmkzWm6kxHbkf/6MSG2w7cFRyRf84nzHVNgmeV1leLU
hdqMpTqZd7ZqS8UbhKb8GDKf/IZXRYfzkxQMltBrY8h6UFgrJ2tGwyK3RR8/L3kM
Dn8ONJVaZhL7L+9GIfxVKROh+WCz5LBJh/Fe8b+t6lYKCwfoDKyM3SCvlKDg+tCt
VytKvvarh3LBppvRvJnNAiZUN6ySIU7TqLjcrAtb/K2LlKfXBm3HPa49W7HzNHj7
Oo68V1fL8zCTO5jf74MxG3AfGySlF6/dL+ZyqNo705lNPTw2ORS50jaFlJhOKOH/
2M8p4F6g3sRly8W3oCMFcKHFEtizP2CULK2SsbdF5nEUy48AFLoJfGFwZrnwR0/I
HyJRXP6Wf9gIeZ2e3OvjlVtK7jGB1Hb1PIIujlZID8eeA7LNYS6UTzRc1ae4CjEI
BEduyb+C4KaaH8GuhmYQpdXNcmcXq/7j5lQX+P4fiJ2f+a1XKMEQKp7ktDOaUrTt
kG4KM/iXjp0PBOdUdH/Ea8ECSbrAhxzwow1g8DbQf+jL7N7qa2y/3c/10eR9WqhN
bm3+7Gjz5sPfboHFdbt2et8/2JKmBmS8P4DKLvYLE2SYBX15+DLtGzGcreEziH35
oIHldX5ryAUQuZt8JQwkRxx2FPmNiIPwqdTAp/Sv8dLa9aKBj5bkJV5Qf5FGrMbq
RGQ6Hsznb1jnWahY+kFeq9VZwG0auXmaXlcloTCyT696JaJ3IXxMj+o2kEsH03nm
osiu1VyTKpTPZZWlM+kFGB5Kkbxqanp04UPpfgbhLIFYQXD0ju5Iov9LjcN+2cMg
f7ORhYu9jPek0A+n/tmqrprZYt3LdgEEdriC5gPo0pipRl76L6cGkBkVAWpvgKo8
eYXYGLYuputgWDUMUlpVg+avEN3AODrfKggM9LJ7Uvp0MO3d3n1KoUHwxVTdjeFi
DAwpKRDJHa5POJ9W4DRCuXESGCs1dHZSqCS0nEGcDqDYpL1pyPagcyTZ+Q+VAELY
G2f6gsu29eXoTXRDFhicgFmx+Y3C7Q4RurzQgO2BBVS2qJqVGMUA+pMogotvjARd
8MpfbOyU6YY2maQmSWawfpjp7g3NoWiejE6B7QIGGoozzX9zQkiR5lpfDL/EmmiN
W5D3Uv3grpOaCUUEuQFZP9NcwJrOGzN2zP1Tud9s9fYjDf2KFzRYiPyyeUOHjDOs
BrIUmy6Nd1hx3DaevX9d33fhvmOh9th28yf9eDvpO8+rBtd5KReHPtUNVdN+q3ET
Rwr3GP1irDk5e8/ds2mQm1JfzBGwajZC1ZDSh32p2dmXGk8TC00ZN+dGiFXW6/a7
ulbsBzCyqWoMkldzbVfeAIDTjvAe5DAnXqQhwLgsei8eiqX+kEmwVNcdm05gLZf5
Q96yQyBX1J2JHipyjw2fKHamZnW6AbI0BRQG5US6j33DW6nZ8dWJCYrPbBPxk74R
EqkVigot9xAJC8fq/eJphnn93QHSzcrymsd6LfXZn6KoCgaHrBS0QM2T+2ugJ+Ix
2NSAJg/n4IK42VDByAnwqvhRRhr2UrENruYJ1sm3oX1LRu9hCXKwKkFTZcNZ7tA+
8Dfiz567Srx4IlUFZu3fBdWK0kivUkReQbVuZQXSSDKmP8DZsHZ9MTpFbD6rYNBz
W6p9XsLGBQ9lzO2ohGWql8jZsFHEWZe5bxO+Jz+gnLtf4wBTvX4b5VSNse7wVUn3
/hj3NX60+olhgfoaBoFLLCpxb9RGGtExELR+gKLv5Dfl2oNIHUuDOsJNZQ8HzhvB
SfTygkAsaaFozxIUoYNEETWpQZdX4vgN+NFWeBn6uvi+SuVxpxkKT1sJifqp59q9
L7tEocavxRimEjB7rQzlwkwUWkHuC9PJIvU3XC7pGJDqTcsutb/DlSjPDDfYFkuC
czAdMWXveuYYI9Y4Mk7be3ehB1dccN++dmqmoT5a9mDuWCHbqwIhMhbyByip9cdA
Q7bh1UrmccRWdRnvS3YqMVibCJwhtzF9Pyl1r6BVbadzeh6JB1dqTcRgzK5RV47i
jztWq6h7KUgJdwzSq63VAoZFN4ENQQ0bwRrVfG2eZbAdbZkgLeRlqGR4yV52AKRs
Q6W+KwlutDzpWrGewO5RpYJG4JakTKWljP92+72WlyFd02nnOvsnbCIdDmSpeVVj
+hWTfBFlrZX8DnW50Llc+FVWCQ3j1cUr7Us5e8xnHjVzywskisdgajSPxYPgwOVV
DScQgEKotxsO6QDZfrCNRHGHf5W3fLO2Su8y/72bSSkROiJkVslt/J3OESp7MUwj
XESv9XkkUUr6F2YZ/1MMRz6S6jgkM9iHQVBkhW+gY/vUXBNsl/MX9SQNJBphZGU8
24tkqVbi7++uFttvrajA8RXrS99/XqR5+kQqTelqpiLIGFWeOZBvpPSOTnqFvzbs
C5dvm90dFIVRybP1hRdJ76XmZF6e2REh3R1XR2PO1izRRsnobZjXmD8MmULihdzY
5y6vYNaJ4tOnyIFwbUox7jFzOwEu8tzFFFNLNvAFbSJ/T0kmXmWp5YFXQTI6ziBR
yMXtcrHfZDB0t3yAhXn8byLWk5mOjGE6NHfjPSx/YCgn0G0dJBOv17/E7G835JlZ
Eq5EkpYV/ZT+lGzi0ipo2RwoZFZG4d7iypMN3Bd0HdQQV74/B5Rvpite4eO9+fXA
fkUhClvDmmyltQ4PBEpl2eM8PPvD6dHxagCfG56BxpMgSD/2nFSPyn5RaRbPtBSg
hS7W9xIyojQOebo1csZdoeLR+WrShRs4Y9ovJUKS2Yg3Li3PFnfjY41XGqEev3Yk
LBnxsmSRJgXOPmNPklOLXDN9P2/+aFHMTm92KZeHlBC+5Kw//etu31KFYawi1IDP
LSzAnijYHO/SJbsCkTmXGZstYON9I37qvQ4kDpVrJs8oL+BIsMzLUYzVjJ/L4lG1
NJt6WwuUrZK1RjBUeKlAHFLxRsWuzB3DFZ/b3M8+CdAc5fSYHZpBhd6g3pvVyRtg
ZBJ3+Uq80CJOByI9RixstNyR8gdh1IqRMHmsD4+54BrQ0I+qCS8yWpMI6a1Fxhy7
x8vDhE/bZ1tbByZ5lhXXqaaxD2vzlKbUKtyq48akwJfV3FLEWxb2RBKsaEnevBiN
byjO/eGBva8OmAfWmt+NmRwaflXlJuZlmhRk7J5pcV0Sp50MiG0UfchIli945dCW
tKZl7UELfFjtyvevhRrLgTC0xVQ+9SEjrHldT2sWCMFd5/2GUzWHJXHbf9czjaNU
qlsqKiJ0lAmBXX0bJVna9j1b0EyR/0kLezVU6qCEFXTQqkjjRvrD1Fn6lqLYjmlI
jo8vPvG3beZjWlmWpdpnbOKogKwhLdhUNi+AKmZWSjTcOuEthX6VzFGa41akupss
1kbYXDy842qNXfYDSXNQJZIJVSKVKBRgjH9QSEVDlQuqu0cxN8jXwcOnpnJea7Ut
zHqzd0nITpH48yzZ6HmvbGJ6tVERD5JjpXOhs6KQqva5RwiqkVfinwZH0mHaDfDs
BerT3OP89A/1nNncXR08vqKOXSrF3sfR2PlcXf6b4mwvtY6aGk/WsQQEam22D3Eb
fSKMqpocYwqdu4eTYkcuxjA1T/8aNaKdCP8PH3lGwsfED0nkljgui2HuE4HBZhoC
nz4AouEjhJNlNbEB38kIXJEIEHhULOr0mtrpZGBK5Nose5qBgV+bEX/rgmhfte7K
KDoaaZpQtxY/2aEw4XspTo2UvyZNlNvr2N89s4ymJOHwijkdVh8FY8SfjOc7SlBj
yl3ppU1s36NkrEC7iY5NBomKvOitPRjJhi09zMaW9Nck/s8gXWJA/2j9DbhzyhQ+
+fDufLLUxgdDTCsCoRR08xT4iq0ccWq/LnoB44aE6lhybrKc9ptNBDTHtqET1+kJ
WVDpiocNBq5zi43FouixjMJQW6boA9MXazbPEhyzoWPbsmPQB0xUEGvzXbasQLeL
BGmGljXmkPwZJ/fX9JL8eTNF0cY2Oo4gKEwnIu5QhtnjdL26IPXE1Zm4VkvJGyFQ
iiyryx6bqaQsmU910yH7IWdHQ2fLA5OdOv3pORR41O1hR4At3y4/q/2nHt/HTsXp
GVvq/7T58CwDewGiXMTT23KZdupwYJ1DN2ERcbIoh9OBcziVgdPWqBVmwdNpGOGy
T9JZsEK55j7iJ+O9JQ4PqfOR+4s+d3WJYG+SbhGIHLb+v7pVbQs+x3/XUwq1le0F
y4+1deAz4oV97Rb+LLUQsMhlLft9zvi52zOrzsP4/ojdpEN5a35TTxhOUAMLo2Nx
vY9ua7LTpJryII8L8yAjBu4twJx32/GqV/e7CTppS41tfSveDD4RDVdUFcM1psHS
DPV4m7JSU7VDXupw0DFse82rI4uN0984FMOxrjI7mupW6wObgf3WQAA87p48ZXgC
KiS8Vaw9KbwQIq0PAK2/EUKYgzcoJyPjDX6wo3vpuXZMU29ns3MCFXmLFO+K69Ea
GuqjA3yJ62TCdfSnYXYIakhxuipcKfp9sDl/GbYfLNjSghHS7D65qbom+1m7FFjp
OR55bFJNXXUG5swRgZNiHTB6sMpUPOUPWAjYUNgHbwjlf9YBZ4Bi2t/hK1ZDN6ee
yLFOnnuiPFt2Mj9IWoHv0NyTwYLMu3jBB+D8I5bZZaHokYBwu5Nzm0Oo+hxhd+Kj
3jEs9AcmI4ILEzcOpMIrN9BiKepJ93Qia69BC0jhCJT+f0nYm9goRjuD2jm0wfg4
qTUgIKB8rCVAiGqNY+0PVqzrcwo557csH8s/EAqFBJTV+l7+AGCTrvZsYIBv2LnL
s0Ljz3kAmcmLRhe8FbEy8TFg+GYCoaD2idW3atJVoNkT/X5Ej2WpDAAcuKpgaW9U
2h+PhQuuty1VxPh8mENgy7mbk2eykQppdnARkq7CcGZt9pJrl0XDjovwB+LKZUKd
TU5op/f5xWEnjo1axePvuZKjfZSNwr1YtPTRCG+IvVWbYHACSn1K57L5UkBoPBbi
U0qv+qdum7ly9Plhebjhc3BMcNxOYlXCIGot0rb+IomN66GvNkfLBc7GfcVK+Afh
wR2o9WJpi06gRF4kzKNPkt8i4iH0CjVfRLP2WFkNtZTwKsTOkB+/gj2MSvvN/cL3
SdPtGhSwNPtSYW6YEu+ReMeBlm3AYzpBlbbD++LYW49sXNK8EXVSzBdOa4bZ3ZEK
Lh7opnM+Kgx9AgtPX4v573B4EzRWig/t+DcAEZisl9gg+eV1KV9PTVf/aBTCdXCH
hRMKEn57+pqereOuwWfqOSM+xTEEedJY8ew/xwuTv/YHJ1O4TbSGcVpHHTxogCX4
0gbP8kbVLHa6pYdI7hUxn89219HRN1AZPp7kD6Kj1bFhM6srMQx+HX04yqDpgTjb
U2D8HoJ48Ans2e/nCAy/cKc+1FVdG08bu3beC4r1Jkccz/cIecwrputEJWMxUkeM
3SQajzMDzMci8iDirFoRl2btnrJdjBjxDI/cW8qcsgRH+sGsP72k/hDI2B6d/YHx
zCV7Oc6zoAXmytYOYep5QEcl7jWYpj6+4EhbaIzVxbfqSRcmfihfl44srOF6jVxo
7GsjAguzslWvApg71Q56lpNoQ5dVAvvyptdfA3mUdBv6PAw9qVyDHTLU4jgnak0t
kafkf8LxKBM3twgzbrZUeb0JohAIUUNLTgA8RkPYju47+v5BhA/yeU2gZn1TbUqG
wA7YaDF2kd2tM2dPSVL7RVZZz5H8N6lJ/+PeQkpMDaoUNjo1BFtwm4A2JTq3VjV5
rfWOcl0EN/OKjC3j3zVXtIWsg4MvpOqT8ZMxA9/RXPno6NdThPPVNynDprHXA1U5
YA6kf31KdmKc8ZDtyiQ/g4IH6RbXSrWnTnPp9EmzwGNA7KJWFGd+CJmQo1XZtdxt
JxG5iTQGnfZuGoGNleemrOPM+taA3KoYfesT6i2dm1AVXQkkImYHiMRCHrP/UqTF
hYYQguC9LVQTrHScG9Mj3jhDy4px5dwmg8qjnNOUDB8/nGipEWzgpXqF1BaNg6Gd
bigs7ZsUk6vjLpFuY9vnZw1kC1D0NlgaYEHE/d6GcLyRRCzOtGQsq2p1uYPsLuOd
QSLxz2nzO8d4VbqMZ36jFLDHBH6TwyYQbo+/olqpRuxbcwRxvgsTfGGvueECPtQS
2QWu+BLyf1O+Tfu1T5K+n9TQmFnbatOLrA6x+O1nXQmg4BowvQvQO5BbXO5f8LNW
0DSV0EaJq7gFYQx60er8Psc2YkOKAS1e8CSM2c7fYIbR1jElGl293J+j/tW4UcsU
6gQ25YzxIPirFWPGng3Tz9/eNi2xHOxB1CULkFLiszn794tjnRlObkS3hvJB7XLP
blwox+6zV/0TGB+1NUiDSa0bVH7ayCT0P3l6VwjVoWQgle9uFRcbpM70g7qR6fGh
iMRy3hun/OORjqw0UEMXxE9t0lULz8Z1TGXJ8axbkM4L+yvt9rnbwsZrJ8UZxbpt
yuo7ztEujJzsFFhD0fAfJxwMmrYvZvPKxHDrZF4pBA//MX+QofpJZUrMSzL5gFtU
R1R55zG0OorWLbN5gGMo0idvfeFTOadaA2Oa7sU1JDntim4GSRBQke0oaGJCEWi9
kugeglzmTmXAWWgt/RcfgJ7IveruYl6vFIL4oltjyhOcqPzCIeAkEJN3SJOtDax8
A//HUp0w8bOel+qOkPalVciHvvL6T8Du8AaSiRKaA+LBemJ/5iFEt64PuHbnt8sD
Y3/RYXsoQShRmnzp5HreyfLv3sAz1OBLdAMMs+0WJv+0L3eKKukqaB+Yp/V9qMTM
Tj6RPCB0HOpsudVki+i1ShFct3QrTyuCZ/TMKjKI2SqZmCYS2qegnFav7FSyFNHd
yhvH/3kFBBByG8a+vLIILNTLi87UbtodkJOWX1FHB7XdN7cth0eLuhVGrJkEMg10
M9yy9iKIeIfYk2gAgR/fLAOTvNNXjW8rVQ0jE5uEPgD0mWl3NjhsgxXC9dqBiTtM
Z9qnR7/gG+vOIVL/8zV0DsPaHefrxO2sk+E7+ZuyX0ukM6FxA7InqDO+Bow8QH9e
S58veZItrrpIAmQOIuo9lq4QeRTYRemwcb3xhKmRYqg5Om+IurJ2cxvdDO58d6HJ
IHCYbo0W2gpXx9ca/S3UsDvi5Hw9BWyCNg7AlbaYJ7Nd0QLJJmI5nr6wzVt/4vWD
EpisMBdEn3BFeIHwycJw9t5sPiTNdrP1wN8RR6IJZuuY01DfVn6JFaEcuEAotdG3
sERFMwsqISNgH6QtupV8sk2tcGndCEoZi5wWmjWO+Qn7AzyU9nHeSrI//PpY6E4j
jbIHnakVt8LTn8wjX202c64QrxRogKxUpGthVKZU9T9aoJ9gAgWv6tKPbUKdq6Nm
zfQZ12D+Wf3ZoQeAj+gpRcV4I3APEsv0PYNmVevvjnjvEJd9ijQjEo9EH07nPmeP
v6rboykP6/IDB3ZXual3/mwDld/XM4fGtlt8x9fbCBsBTiXlwIDLjHw86WaSEIp8
X9zIVBlD4Q0q0qAFSI3e4bnrZdtEiYJ8ozvjTT/HbP1ecG/qkM3+yZHj4orZpO/9
ThUM9YIF3qbVw+X71BSFtnc6gGdfF4hvrDajLnBs2UycClRPkEi16vstDRfjiWye
8T10sNrGBoXCUsVOw9LQie+D+csTlq5HHymYJDnakSMpBz5lkYw6SLxqWinxWMkO
qxFkbPZjbR19ffrQ6qVQvOeBZ9pywQXKeirtNCiwtdzgAHvKKXuORT9jbX0HJVKX
eHXVtDj450UlVcysefQdSlB0KcqH5/upoXcH1MRUgg1zUt+/i8Mqsw07z51wh6xn
vo8wGPMREBYXgGLYbXfQguD0R/CvKCvSjGEoaonWsGDdB19TWvtZdc65GjXbnl53
vW2GhJcfwP7dYjfdhlMKKsC2jPUJQCFYNNEb9x90tCzi1Xe3B4Iv2Z5h6b88DCZj
6IqfnxBSm9F2rqFlxR+SAYfUqE5C3riuUv5LOns6GGKZkZEdGb2l7RIs9CHRj12x
BWQ/fQHaP1gLJ2DB5QU/aGH59u35NQbrwNqi/8kG4HmFWpjMvRHt4Ec2awoFL2bk
N1V0+/WFvWdt7RtxguuxWHaEsqLjk4vqETiBUS2P8MPUehi876HlVjNj/3+3Jc7E
2qBGrSImTl7TVnahmGsOfpqfwmZHA9j3TORacpTf6eSPeVCXUXcZEWDZAM0lJxVe
gqAcY9ltzZahCR76GDVIcSbQqhq5WrrLYD8RXD8amvE5KvjLOFVKVcR58tddVZjM
87xA88Aq6K/34c18mgqvqqLnLZygNmvuCu/g/5udAyr2PrnDKL0GbM1XfghnJ43S
bka2SaplFVH8aiD1iyP3Cok0gv8eFZgv9gD22+3C+1gg1HxsLsgToLOI/zEO+HuW
RQ8op3/r6znO220GQi8fdjgcfZsSpOraw7NhD/qlPlWvVBufab4cWz4nuhm7GMeR
aSzr+AXE8yriFufcnFKWvwEilE8dcN1lSSxCSqU29w27yynBCs7p8vOcbRTAiS91
PUVrWDKeo/Ks7WQten422PnaRUpMDvF+/mFUkeYC0xnuv4vExB08AmOs1hPqrg92
b3VadX7GQ49AgecRT6tD0l7u5bgTmjCjjzD28xpA3NR6vmNUMpuPhjKRADANev07
2uOQ0NIH5zAlCP+GVA3Mm7mv9ki7K+um+n6zXXwWdFR3K2qy+dex1lY2sxK3UGDc
/m5z1TBgIftb2L3aO5iNXgWQ5Kr1ugSyis/I6xHijh/hN31DK7Zx/YTGWCLANbr0
y/hsBdQH5ix0BFK5yb/tUie5ZdNmSrI+mV9Wi6sAjNgoxhw34WWufRZU+vQJ+3jG
UoDhq2mVr7Rj1GSyoiLkWMsF8FrzcfDwi6ijbN/1cy/FmobHR2XLKb2yfaOTUXHD
KnzCOJUOeu7Y3lbYl/JJdd29/VTGIYlJnQlfJPdyqj0zcmZ6tQnfiWMONl4tH9eB
o8EIdr6GcF2BTTWSr0Su1ebgbx+nhmSdK2aP6kk5l8usJYBDOJte2mPvd3JcsNET
XXkar/HlP8aoWDsg2Zyn9CENu5gCTmH5H1QPwsj8L2q58x7ntK925rfZaMdCSs/h
PYynfwpfhWs5QF7WkIE8dMeNlE8rG2eT1+VesKVm2UoGcRR5WWuF7JPrQPvoR7Tb
fruXP4vVvUPL7d0AaXbY39dJjOhphkaqeeUx5YwvnCZXXipyKg7e5KlrQoauA/Ya
NWpV/UmxVvkKV86bEYfSGu5uM0P0GKRwye6L45Y4AYTy1RpKfZaDWnT+cuyqKayi
2YhdT4oxlPCWJIzH/ZDIzZclFiDhXW4ZdiO5ngAOTbJKALdWSJ1LWn70IkaslCyf
G3cn7hPVqAxOZ2Nw5mOotHZnHvWulxb1R4MkAR3pZ+JZgbon1NWcJK/38uGn7WWy
yoQw4RzOP6lqtit0kT9Tla17NcMJmekAF8VB6Iaj2z0F7ipkDsK9423dMkSmMVEm
80Ql5oKYe8maKPsUaBAPIjvxgVHlc6bkvhqTzl0f0tGA0A5ouBOiCdf1wUNxdSzl
CK0OydSldXANrbJS5xlkXf1Vrm9ZxOqdDLK/Lx/lhBhtMYk9/bU3ByJtq2rJ+JEg
zssELxgkrP2cgJfqxsGOR27fQNx9FOveSFZPowk6aiahU0ZvBRILBDGSJ6RcWsP+
MY81eSe3GGmJCSeg0C4vUkj0ws82GMJ/NgvrtGQEUMhGD4r7RRaN2wv2Yt8lzO+4
qJekMOdMAnDzi7LUUHczA6C11sJJxKCB00QUPs4WObM3NYC39KxPvRDNkjH903p6
BBUkBjDK5c9wBJLP+1N/wZXBOORcfRoLy+fwqWgpc7a0kup6XnJYIZydvXzXE+lH
XXRRa6rKE9iPnqcroB/kKCj/rJXL5A3pwN5GGOxMeLKx5cWkzAI0dvTea5NILIQ0
VPR7op9wZi3nf4A3N5GPSY8CfFLf4bZ/7ZHohLtSa1XVeq5ptqsVtlPsswP+Ts0H
8jRRopepEVHS4fqcvcbbffGTbpOTeEII6Lno7L5xeiCAFp5yNWhJsQbHGad35JhA
9CHU4hRWrqR+5eimcfeaexI26gkfVLqqoXtxNIcoHLKfM6b8q8Jb1jbw0HYgEfIa
Qa3bt0h38lVPF/ReoEw9g3M2oyB9G6zhhhwH8M/19P83hEt+S+gazXlAQ/ls4eyx
AsUvFKJbskLfBGJETRGQf4mIgWBUTrFp1u/WpnasQubwNTSIRye3CyCg0rZZYcZ2
P3Gkhlhc/VRxVTOpc5iXh2wcLK9hBz5UbCmkMSscMXGgkWHc6nRnTLFeOaOfZgrT
F22LiaUOsOyXs2nr6beRtvXhsVs8/9G/Z/O8mGZAIJhqN1ZDTJtvLizswfg2Fu8c
FAek13wmocCBOCNZbpvACc09dfxMarOP7LKWnMLJ7wU9hnhmCjbFi5KqysaPmZtY
qGCxSEhWAfdAh6wBVKUd/xjSGa/s9BR5NBnFz7fbm6zioJJs4NG4eaMyJR3+oTx9
E4ocSaiQm1wS+XgPLFj3o65LylDct5Ku3mQGDZqo3wuWh1+byKlzWvzKsh9uTVfV
2yBd9I85hWT0IAtKRnB+BMggNf4Orp/4nc15lb9ejuxeG3aU/NDhPoNkDLsUz1Q7
U/yHlOrLJ65sbC4h9wg2AA7U/PV3eWIECHqjgLkc2V5x+wiIh9K1Q8UyESiU+Auk
sZOuO3p+zM/1iTyGMTIPmA4Oevg3Bj8iYuHwJjD77ePmkv5Y3O/PjJawg3XUAYKf
ETXMowWKk3cW0PQGrRbj5EIlNCcQAX6QSRIQt1YzSULG4IpjouOOmSHuLIj0QJIN
hnDGzEb6veNBPGOVXh7TSvrRk/2Wnf26rmL01xFEJm8QC2qXIY6+MBNOZ/ftq5tc
KLuI2LXQwUv8c9pTMNIGncmXJ9BIR9lpifqa1/nAFcqzkqvXWMaIsWg/af0I/iA6
++YIMHghJANWd3PP7nL3KUZ9F8COb/N3uaDEudpuDIoW+kyF1XxisXJTICJLcg04
PysPii5sDz1gzXa15z9t18SNvqe2vYfHNHxPVHSYSYWjUepJBVpgF3FVYUPhl/Qu
NRhQNUIE44K1x02rXcYhyKDbjjg6r2dK2QR3GLJKEO4zq1UdjdOVRjvzqGjMNkEC
OZJoVtmkt82PYyXSaoyiJribybt/dCGX4dF4H+uL+hRUkLUXkoppWXdY/B9XWUsQ
k+DcBtYcCJU+fK5jrGPjiXoF2PEmcOUOkXydke/8RsUedqVGwdSz/F1VuezsbcXE
K/0+GPE06SskKePPj5vt38gS6YyDjW0ebAPDxf5DJbaw5Z9OXgwipsO2VP/wBbWJ
HXoDAlhk1gyVb/EC/28e/wmL2Y7k9xuPD7DYmNiI6omNTpBuMvMMHsvK1CuCjDvI
fZ7FiRzIl126MrgCKzNKy26rz2m6FYgYmDBdhkacCpLSgfsnxoUGPAEM7r6lCO6m
h6mgk3pXl1nxrjQAaUsA4KSIEvsI/Pdw3RHW1dnrOXiXyS2o8vR7QmXvGA2DhMzX
tJJY9bqLYxus2HGUU8yB/i9JDN5CvX+7Pg7zx5/96+gm0q00P/6Lv/f5kMRURERy
Mdpice3/M36EBM7+waZqHgPt5E+dH8ObDzbMNbBxrbJVnKQXUnCuQIm198YoPOdU
F1647CEProrbEo7kqPJXhBpEnsTYVbWHUrlp5q6vdIr9psuTdMg2tzswdBkhWHiA
oZQupElHEMIARhEXRuyqqelWr8JPMKqJJKP/AU1ixtdNj0n0qSSCP4b/Qz2itY9+
7dKFDthmnnIpFWqu708oq1AJp5xGqQUxL6AvXJ3l+1y+Z+3AnZQYSceein5BO3tK
XXi6U5uGodjzPGUMCla9y0A9CNnqsMHG/odzCTN9doRDSqdybNfhY9Yc1D5mUMkE
hbw1q7lvYY3hZEY3vZjTZb/foFvocZpm03dqyQnCqXpLcaMLUza8LW64+gCaabj7
BmJKiCOK6bLDgUk3dKYedtDWDDFPcctcXAsqjwPez4aTXqxD3rEJA6tA9EzwIcFy
yPsH1/Sux/FM1WaBbRoBHKopUDCPOASkzQD8pXBczjN67rqm227GFEKkal31C254
R8+kRkD2j/vKujp6aMpS5qCTWHdFP6feTTIAXx4Dvn0gd0Komn5UMiThemELqw1W
d9xiOSkyKYTCWpriUf+ZZJy/ybhanJ+HRVxLSu0plGPjoi9DcSKytnuQ6LOirpxr
L7WL8CKNnZuNX+q+df8uNC66sAhzkeiYtIJCTSTmcBut9PgtdUd6tA50VJLQm3nN
RRFh3RVud5mi7AcA0HsBpT4t3EnrYIkdspdGGAQUPqpZEZk+bVb5TOnkvdDUIzV7
VP9uzNPOGwvyrV70seXv5JnbRHQon97UiumgFV3cli/Zgcp+zmDf8wDS0vdR2hj1
PWhnXvCR8KqapYMLAsWqjFiFI9pJtm67xqJ2SbA9zfjrRhGutLGoGKQJGwGFMGEb
DpaLF4HCSFwx7LSP+5pJD6DCaOOrw/0Zn+cNzPDlDfyRb2m635Y3A2bWitFDUbG/
MwhoiMLRcoqFbT0DfvpIufC4o3zzgAJrw88nSXMR3FCv60ahnU+/ZUwfXsljats4
UO1uXnBdRysbIi3gt7W0F0VOcpvS9tc21dJNEv80N/05sNu7/YY1Sy5Ek7dOUXy/
0Q3JguhJgyT0Nc2a8coUxA8uUtaVcHTaFJw/DTsD0hMMwQCso/vyfAXW+XyTKSmR
un+qXLGS1mkdvy4PFMzUTQ7DKEykdD9BGJRyGi/jQQXdn+a1mAU7NTaE1nCeM4Av
M/6WybQp4PHOviR5Wk9aDQVCpEEkvMyxO4faoOhN3gWfRicSZGmCKLJC9ZvisMvy
evSe7cPGuJjyUJ5cccZScncuYLLHqqXcAmOrVyK1qRo/uIaGcYZXNPdmC0l73csW
W4ge++6mU1GJK/J5lZhPn2y243nWZXisR4+6dUNZFcg55iN5yug0gpcNItOrIswT
0MtnS+zLnSSO7LP8i/Onbx1IyPj300tp3434upRzM1UMUWfJ6L7a9XCRzroFBhpK
PrQf0CGNIujnHZwC1DqThiPxQxyKHaxRIgCf4AEmopZlDeWg0/QntwVdrDoU8HN6
WnLpNa8O+35W7Y6YR7DCEfAssJ9w12W2791mUeE5LloK6t2tYTvg18/W3XVOL63W
hnkk3TxgDBNuSsQZw7PArIvsqfCg+/botBR7yrIsTKwg5jiIckbEqe8gsXSKZch8
Ihq7vx8ra1yCp8KNLmXK+Qxh4GqTRTQ8F++0nJl710yKFr68UkGsDIv7DS+WejYV
Kdhi5HdDYVD75u+tWc4BZOCB+E5tJejCkeMAFbfiyMO/39+v0DLKi7ne9sasdnfz
Dj6F17WzJFPx0bw4JPIOGwR4w4VZ+1GnpLHL06goE98FT599E2UPbhWgYQU+7ztD
diBawDNRbVkoP4VloBW1fMVUI7YGykZW+Qhxiryo5RFWPrjP81tn88yOuK6XFQk5
Vc7BYdzffs8xe4dYhlOlZkjwVKUcYKaWxCa1bXhgEGJNMmKQyxIs3RmqkUFssqVV
bA3zjf71UUiqVnXpUXT/fFVqPa/6kNbQbnXo2eVNzjHGcGdFea7CnqfRLyJjUIiJ
9DErVxbtjNKJqOoeUOdhXFDk06jy0Ibh+3WMZNB0eFwS9uQkjzVjh9UJGhVgqLgk
LgM3PLvWc2HRaFMFjABbwdr4KIO+7BGHWZC5sokM+sIViVUEB5rlL6il50X9vlPj
wvTDauc9YQbTX+nRg61ia4EHH5ifcq1U7Wm4aOi4Mx7LoacZO80eNjGNxtRK+yZs
NCilmLgX02ZEOtu2Ta1m2MI/v/Cn6la/2quDLF6x2pwUq4X1F5m0WSk/BzCFMhZq
ElI4MnuYB4T9J7WlRT5yvZOxaTGMGwiotWxkCUtmYFCzLqd9+KFtXUS1Qa8qwPg9
sQaOKRew91S11smRVtX89++fHTWkNvkrqGxKJLrzypc2lKOzxGq19mMEJFBtEnyl
uBCqciOcDJvh3QtSP7Fo6tpbyqrIehUUWNIvMAmHzmK+qa2z5mxRCC2Ukf8rrUz5
7rdQ/3dCPQArTxGK36qI3poHH3PRDwdhDPe0c+ukS6ukPprYwTBHhiEktEq2GE+a
h0WF5u6mfWI0GH7tIGLQq1/Y2VhTaR/f4W7Oz/HTHz7mSHuhhyWkMTT2rkjCsYWX
/Y+Ep3J7JnAyXNCRDTt/kHAr7fyIV93xGmL/WzmxoSAEPg3+t2lS1Q8UsuK7k6Iz
/PlDBT2iQ8cUI7fk3Xlfuo1a3BqCzuftQiez/9MgdhwY00q2sUsqfX/Aj5ncS5Fq
/21vyF5F97OA9coMZnNW0zkHGE9sWX89SkBB9OIJax/8gbwL8Vnls5WQUHaOQ0Kv
NlXJLjeT2CMTXWx4qvwWjpyVTjfVk+K3D2Xv7qydJ1ndGi5Jp2dQLTgJMtyGg+6G
592HUNEp9L8AFizXpNJFeMCPzn/cZGcP9pxZQLo9R/4vKqwVVbYIXvwjnZPaR4q+
e/GcvKoCQ8p9XIAy/bKqJqZv63fyTQPsVFBN5xyHp0gpVyD4vbdmOUldhiIsyfqP
ysdH5jJG9dAymJT8uihh/EdzpA3vKuwcDGPzfKJ9GxaGJfzkiWvGPkXda9QFirlN
CD33GyGGFW9Vy7bRUwgoTcsJyLSJbhaT0r/I40CRckF8p3LWzqCOY/HoTFyPHy9w
OJiCQyyl/NvfvQEKG15JT31Yc01/0iDvgS0QhDijZTp8z3niq/FG6TanocMi1Cl0
X/f+KeD5BhaLfL/hjNLiQ+QJBcuK8nLrMVR8ep9j3H59ae8hR/5mLl+mS2Ps/mUJ
s0Xc59FbM71a10qJ8SfNom1APX7uuxgLYuazDUzVTw/sXjODLFBFm76pcRoyEwGF
OMnAHTpr1eLrG89uzE6YLWluXR7K37JkV54j63tK3FtiLfewLLympMv5jD50sgx7
4LECCGFFac2+t7PxyKz1oXKC0QNXVxJBoW1FLOoq0hErFk8yVP+3/J1vPQW6IaX4
nV29OUgw+IW73++6TmBZ0HWsOsqEw+aF6fZR70nlqozyLAvTGB3FdB4piYh2T6yh
ru3c06XmVc3b01hdhXNSbIt1fYFDiJ/nZj+YYi+tbm7tbREP3QoOhGM0C6sBvTHv
51rYPuvmYV1q362OyaqSqP2MwCgM2pNUuGU4f56LuFatolAFivL73mGcR4CR8szE
MHzDWn/K1W7OpbF3ltVp3hmLnAh6u29Jk7Y/RsTvuR9wors+T1l0WLbWpms41FnE
GgvuRHJcLrjKPgFYNxdGvZyKZa3LO2axUrVJZIf/nJ02flHcGkYXs4K5F93rh5/n
u3fv+juA1f56RCQAc9brh3+02+S/guXsUlQjN/ZQYWBceF7ddTn9Gset3bHnHdBK
AQWvRQxzYdERMZIFWQ3MeWTTGiyc9LWq3FRuOEmDfhOjWJaJsni7joPIQWaQkGsA
k8DEv+0d5Nnu57aG1hM9ZEm3UkJC7eVOyQuUcZZE0z5T3TijmgIWGHcW+tuyDYE3
eep5qGsOIsaImrj3TmGEpSGplNskUKs+9zblopHo/QcxFzHLAPNg4wa5T9/mR4cx
Xu+Zn/5+ADtXbDvJ+Y4+9EstfxGXMvcPiIgVuNMS1v06eKllA++kdMqN90QZBk6H
ddhSLoQ5Kg5cL9pstIkw7ZoLnq548aNabq415ETakhL6E37n7AWXhlApRKnEG/2z
6mDcW5zK0slvQx2Y6+xfyOL7GzgeqYoa3pvfj4DIy/e5kVS7fpAFMbm5A2ew8zAL
ex3BXmBdQ3Op/cbPM1qCRIAqQF+XYKYDKLypzlwGwfwB9FUvrZdUIpUD4BC+LOM3
e33//J6LzZQG6UdzY1PbqjjXSronvnccxjrBRcd17ggRi0mcWZ4NOyHjWL0Zt3TJ
WdVTNJhoCXKfVxVF3Oa1xYVOoYpJ3zsUkUyGmaYdGXJ3g+dRKFssVRitXS258KqC
az5mI9TvzLMi5s+AiTJKXjf8c44Em7VfXmSyUixXe01xbmpw2xaHLd9IvxW2/UI4
Edlsz0riNtsLRlgCFJ9v4zXCguuOloo6jcxMQ/zs+VoOMKPZRf8Wj09lEvlGYRe+
UWlHIbqibs3jlsPO0k0DmjBhI5Etqfl63qFc0R3qNOLG4rispHGbX73CpdQukv07
r3t99Pi3ZQ/AX2whNLJb1rjpIn/K1XGliq+ZxfcefMfp9IHIwDyji3XLArHlDZ6h
FjztnfajXCtmaXgt3pJC42PVqyR2+h2dHXvz/57k1nplnhl1+uF//3ZkxfgbxgZF
E7pGSpyNJ9sud+5mhBh4pKUh63/X3GZqyniP6i0R2jioB8ucSUsqxPggJ1+VheOT
z+VmSVwVg/4BpJmoQYrsdYetcX5Yi4kvI1f2laKG/YS+w3WYtjt2WCOnpyEUrWJs
DWujJb6aKR+mroqX6ngDjd0vB3kxS/z0N5gh/jF4VW+tlWrNmepTbNPcT7iWK3+8
WNLybH0vKpSTHqii0RGa4XlnCCnXeZmrPvohvBV8rPTSzGRVeZFapaddcRH4oivh
YoU1Jqw8VgSp/ciM+qBo3itrBqhvJ8Dk9CzdL1Nze128tw08n+0E5L6CBz13+KLP
bwAr9lE6fhxtCgTRKZjONhmQgmjx4pUH6QtPLr0xlKtcA4RW4KVuNETJ0ScqBdXi
n/U4dml+9is2G4EAboSdcgU2Gnt3P+7Bi7RIF1KEruKtk2FKM75ONCQw9qMMbhlJ
IaGTyysKJfzSCWkmOhz+M5Obo8zVpoOfGOq619zw8TTzt+ng32kek4l9eMm+9BHs
5aAxN41QzjefYh0DJAXEQHKfQv8opJLKYkz4avYR+WAfZqPS91oot119UOkCTEJg
FT31gWEmIeL2WVCjgJtDTmQAQSEV6KoZ8sAdvt0f2xRNnJRu6jO7MQCqoOm5X1DO
DVQjgV9ccKIN9bD5Huv6zFjhYSrbAmisxEjgGgkE7bi5X1nui3zfPmivglLe2ED8
G9hgdSlWRWhh016qrp5n9OH9xQcqpONHLxZqL6xcA2RssPCWQoZyUn22H6xRJHfg
4Z4lu5a4+gUuTb3Qs2tZSPvv8NuV1QJn70PBAHr0pvS2MP+B7bRPJAAYXSaLHnyx
Q4BaFkDWwuDurMXJUdCU8FjYSynsgepYpuR0NOslW9Qy+ZWJ69dPTZPV8I58rJCn
QqAq28KOkqR+b7aIfNYsgPqQKTWVzMoetoES3bYm6Ub5a8dtZhHerE/u483aW+30
VjPCeyxD0liY3uUckzHfZj3mcfnY+5RhmBekX+0e0hzentGb+BajxhtM4vTzPp2G
v6NZrtts56hSfbx4Dm+ZY91kKOJ6CHzG6N4b/RFaj5Qvep/7aD5a9vxS5SxdXTT7
Z6VdZvxb0SD5ZTLT05FakAVE+P3QxXaUnfzIPh7d/rmJ4Y9fX90bYhJ9wzFBSs0h
CAPHWzRSW2NokzNf0ogigALV8flcFvlRd4isJoiwnX/Lbf9Agc1fwzh7ksUPXHzx
cgSVTQdWcjEFALNzp3Td36IDjzOUQl05IkWcXOzHZh+VyMzudDskN53llOE8GJDa
vvVopGIgFkTDVmgIKkufrrzcbrfUXHPALtF+b87L70PCX3gc6JKaFU9HODbJvyeX
AEiequqzapOZdLfxrq0epycORSMXLgkLyemP+fPyKrODg/q9KFOh76VaY/n1pBuZ
EVhUjXWqOZTyNZByVW6OORdD4vSAuiBzVEoyog2NKSlMPqArBQLxeUhaWphHGS4D
XCtSHIXfBU34Jh0qRwvdY1lCfAJN/v2sXvPw/dGJK1tKYZWtwB7fl954W/G2KPM/
f5E7KruPGK1bQpZvEjPQFNxLJo7Mb9uiGRhLzSfv8JPfyculH5YSpMU/K+97N9Fc
3Iza5KSSAC2WeU5O6okN2GLl4qHgJsEsaKrtYH5f1Gur7KShdWeXOIt5xQC1jR5l
Y6vZBuZJhEwXtGhvba9cS8/r8IjAorFPj29D/Ote1idF9ekNUwhdQBBoxakI7ma7
rhHszPM5ZMg7DXZAhBm2477S9/6/VSFBS5EcBRVPVr6rqCeSkXCKGTeuRa6EbR4Z
hXdDWs0+luZU2ux23bRplfkGjVV3vraEu+birlhRiFyzYKy6a6AS8UWP5Icr/k+x
OUZdo/sFME+XmOGuw/f73ndjT4Z5zL2iV4BpGQ/Z3RxGWLEjni46DzZWA0lIUH0P
7g0XLLnkcFWNTXZBHLNGKxoCSKvl78jglotVji0MV9pzL7qm31/JAzUVYdVuGVZM
01bbypM2+wM4+K3WPJwfxme+NuwSqJFwfKKOyQRi+iSnPJI1QfdFArJWF763VaSp
cdtj6cTumkQcC9WZQsS4zyHmuCfqFeaDXBOZxOZzLTMoFz57djkVYMwMquebc/Zz
eaGhew48UJAVsfY+haYIBPg5bfNeXBe8wjf43rHTwLFiZzXBfgeRM+5C5rLNr5ix
hAN6mw3Sq54M5mw3RYXSvUWR1k04DVvaXvvY4fcRSkOgG67qNQWbfWCbAMfpt37G
ZfAGWwvewsy000XwtbC8IyDSwFEpJ9n1fN3mOfNrL1kJ7Qi1vY/PKvbvDh+/vaG6
x1Eg5V3knSmUAvp2aTas7xJVKcOHWbUQtBC39kqQO3EfaP+cGOuJ9ediZqC+6ORb
/3j0UX4SgpCnMQa2WgDfwk8/RzFHdTYyLsd3cymZluh08E9ASmAvhZSjfFsoG9FZ
C06TuCCL5HCc1YKJwHg/7KQX0ODx/nDVrPsDQMIE6YXLwe+WNVLsWHVvMmiamYPx
Whhjtqo6L/9SKViz+VqcOckefXxr//rFfV7J5emjkT1seyQQ6Z7RNtQZf8eiB2c9
ElyiDOuUjLP/fJQIK6MnUw8NauMBhFeXvn8g1IFZNW6rr66Mx9E6mIXw939B4TYQ
QAKl83UMiSFNyUosl+/gyIPyD2pRCiodKR6Ns85Ymh9kIThF1tlCaGD49pmteJ3n
ohd3Wol48gBkNeuSXczQgjEqAtXhnvPFfSA5xJU8L62D9pT/A3I8SyUPFEVaYEFy
Chqm2QEwZUjuScQw+0gefmZR6nRJ5DdnOhZ+V+K49GAB10+Ap/HcOU1wD4iq3b/R
IglUr8V+whXmvxfypAsgoCX0e4A4vMZq2+IT01pix9owfjpTaXty++Zl15FbWWTp
m1glUcrXS7de9/015WM0UG/LJAChHaGrYJf8vKS2K33tw9DNvinlvkqIEsd+NdJf
0C/HIYtl/89b3AOieAX1imKWvcH77Ckm71PwJ1/Ywa7L6C05gDsQxe9u/RVD8K/o
BN1b2WMdgD5z5/n+qh1m/8QuCbJefxhdEflr9+etykeqFyjTje+l4rqnUNaHO3SY
e/dKXwVfpnDLAfA8gb1+V9x6jO3BrDmvFrQGi/Qpjc8ZfLjmCXjiFF7bE2eGjFRM
/2MHc6KwTMReel9t03P3wAcLrD/6O/8E/bsVK0uDv+o9IqRPxxhJUu952mKugi7e
QVEewu9WzutRQCNjLdtonDWnbe9z+XMkIYM8zjXBDgjjmEVSbUJqdio6jJxZx8CS
KwVZ+oyaQGwMdhFsZULguTNBQ1zoCFzttikiYTtUo9wgBn7LMVuA359cvHriUe3q
1mtlSW2VrO4lMh/O7XqZILRyxT0niLbZveT76rJ2hjRi6Bb7Kweuh3Sf8hgxnrBE
Nc/Aoey6JnM7cPVwaurx5Fss91HAX/ArFGdri2jeyzvUkGhDbVEW3DpEy8kkloXz
zJkQ0mmkRYKttoHRw6sPjL9l6JoEjnTMkCrI3PdPxE+HxYQ2Wh91gVYt92HQoORl
4SYCJTVSOzEDR+CpQxyuBN15JuSkSeUZ34pqhj00YHzXbh5r1NDeyBYaFkyASnkT
Z48Wt0G0eK/AQ+QPaUEbn70jtfAkvZf6yuPbyn24lRiQ4909QcfXEziLrIU2MqtH
0fGkekxnBROUp1lqUhINJm4nHIJ8prS4y72pOdLhQECw99dEWynGbeu6hzcepm4V
ecVI631nzkXC29zUSuIO9xcfyBVupm1cThyENFQjlHtwo1faTZA+ACKV4ejQVaCq
9qa7xl9BCfG5LAjXo1osrpUBRfrXHOdiZqLOaSKHOSwTZfmpGDKNkSpU35vhEFqV
w9y1W6HC/mdRxw9iBzs/oW2Lf86g1p2aHqaOW8JXp3g4jQRXnESYUBhhkNJb/pD1
a90iNVMLGdHY17kYCijI2qfUYnCpptZNDN9vq5KIMtpP+C0zZTzPS2MBi5JXLYx9
/bgPrjAs9OYkcYaNBGbzy0iuFjMWlJiWO55uO7G27YXieH2byGKlJj5JQWadkzyQ
9SAlNXwBOiQ3FGbe3l60JYgAGpU8Q79UqBHA+Y04ELyDJb9L6/7eoDw64NsYSglQ
c9QAA5qs6cBpuZzb7EEL4Ku8p4KldTz2DoD64s/W5exO6hXzwCvcGI7T4TExfdsO
7INnoe5ts9gl10REsdIDkJe5ioL7rdRgXlPnstVqg/N+StVVevZDDrZSPbHEYRJP
RlCzFTIlj5D8gGwG2jK5toYafWnotR5G4au7M3REFTKUb1xYOOoMzyw0ZvegiCxU
o2qyI3whs5Bk9v1hC3vSeDyOYShzeQXsfIELKeZF8ufmC7xMDL08JvLtPTaRfIxd
hlLwAkurmwN5ANNjOHgelm/P8acZaDg8LZQ3ZOMBtGENv/FquC3aP8CmD9Tdt2Bl
NybMueML05zIpGw73eZ1vuJdrl0R5yn749TODasbMyBsYc+nD0KA2rh7tIiQpvsT
Ia6Co6epTTg8vbel9whx521Wpt3plp4AVfZTY+KZoGqEI6FXmxrfNaH9gL0iQU+T
Y/47Le9efAJcDfF/+mPNepfTCO+f2ZZh4Hci0t7OWmkw8uXffGvyh8vqqX4MVXdj
CzL+CIO2KG/6KGphzKM1732ugpbHRr8RHV6jl7bW1XXJ9PgaUVRSjbOqdiDUZdRe
YmeNgyQpYJgiG0fcEoscTmkTHySUIrqvt2TMj5r8dHpNdygjRPLT2dzDuH14QkAA
hmdKm5Fk5GlPMZtddakc/JgyRxvG8YZVzMkEgj51OkHuxPwlmxwVUqwskWWKDx3X
0HtsgKhYDJcrpJ0vBB/DUArTfUGNcnrr5Y+gBAHglQCPAWenztb8So3shVV2efYV
jHAKDX8ImKwaR0z7bg/E8rSyarYcCmVajsRVV/75Ghz2ylsTZPPI8593CwMv/MDq
F/yWABN+HdVQ3JBuO5ynbBG81h/UotPdx/UCRk8lOKtISN76b6LuPN5G3H2PkkUv
e0qBq79Y19eA5lpWK0v43kdvu0rzimZ+kvRmQn/RIfa9vCXFU8kZaTE08QubDvFd
ad1YHP31/Pk0bnVbHyy6bq55fwS2Ls7hlQL85jap6DYlwt6sUkuAOuS5tObm4VA2
uqyo1+fPDhvP0SOnQnGl2FlQ2qHGvCXdIP/4U6tNVix62H6U0XvwGLBn2tcTrYvy
Mmw7GhUuDab7vqtKBUMkdOkIt3yYsmOOnq603vyR1Gkg1Qgg3/0wuatqhWe676+H
hAWsCN4FuLux4SiLnvTaBTbRMJBS+0mcRpPHcPqnHYzvciUOGbODkNf74DiwyzTO
mAVEeb+NjqosI54KJeKk1axUJ3g6Wrdb3qjmsG+f6aNy9M8UP3G5x+qeDu9ZJ7fN
cgWqR23l/C9/AdrM0PX/hgih4GFt16SW8f3s6GPDip8e3BdmAIk8YDd0/9ujpvvI
aVrSbItjngojUD7K/Sfj5qDyakrf+iSSvpH9r/JmYim2DSd/iR1JlBx2x3Cuqzv6
XtX7ya1lnPxtcgqQe8owddzF20i+ys8J/wSG8leUfo+ze/WScgH0kadhmHtR7k08
Bn5PypOsq1eTuewoQCFhMe4Q+qgb5vrmPzRoFOr7J+AAlYOHthgNdgkExX3HJBCK
o/vX1453SQHIPLq6L6ZU8l92EH91vXz1SIan1DVXKzigAKGszMg0wQdmSTsePd/K
fWmQrIrejPFK5ZW1+Dn7SL0QyYhwC7OpxRPiUO4ChXhF1gRPBwxJx8w/hIcuWF1D
kpE98Sji7yoo15X3B7pmHvLcdYNaeu5yuyJuEjP0wSLKGzx18ImfNj/l8qiJt4sX
HnUTAw9Fe73KEwq0OiQ6unAI6KSaKUuNafbr9MCdycEqECTR4nUaEkwEiKeRAJ5c
NYejU8WyWeYkTVq2lHVO+BrjXPoUOpbzvuB3c26ONrAj4UdSJNPvsvI6A1StZwd3
TMZG/joXhLNJLe7FH3XDuEJ9KCvnaS0Rsr+nqPHgKLinMYgC/pkEqtSY5mXNYyr7
W5ETO/Hr1Z7p70sgF1XlmtXgqid5zbhzmHVpHgGeUPN9pD9BRou9K9lf7lla0Y1D
6FvozqB+mFavkDVYymBwdi2qRtlkSLcZobw9bVR7vx3QNmmzSRUWjlXFYg0YtDpV
vZipefPTy1kmT8hBWD4f4ZlIJxcyQSirZpaoqxeyDneZC87hTKac55P+7LVfqBZ6
b5eV4O4IEs7VMcCb89aUsCFRT5phBaiPUyDCgu9cDW+020PFY1NdBaK/xumj8MwD
u9zMW92ho1RU+yP7Uue0Ijv7pUOupqTxLBXyxwr6/CQ0f33SO+ssa3vpPPNyz1r8
pJhWL+ZBAu3TpQL8nbo1gXtOFXP7y72mWFSfw3DkbV4z/2LZ0r/lDveA8A6h+TmB
T1mLR3oZ5xRhRMNRihMoFKp5sAstVUiBRirECS6gnolY7TVkpBDkQgrjzF9hKdYl
AE0g9pXGZPP/PeIacYDAJnIf3EOnXtElIHXLdnJIxvhfj6lR/1hpwh5+u4f9uWcf
A1Df+/0XS/ps+9KxYV0D+0QZnAw5wTd+o9Nfet+QkPSQUcjEGb80901JIK2QNxgJ
NzRd+cq9lbesDU2uMQJWQehHAtl340XmvSCGqWZA78CAnBd+q3niRpz13/ktxlFA
eRuS7IIuaRETKJaL8DjArRcL6pa+FejkQOH++CjB7hqty4epLzZY4LgFnguURTCn
B8et42XnM5GtnqGbevDwWrjlxqm64F9ruK4z5DAgQ7oefDy2CPiDnB0XzIgzJNYL
Qusafx9XhQGqImh/staYC63A+kk5xEQpUxW2wabXZHl63SEy57rsfWSawGRKWk1h
2gsXoiPxCplZfEmCmQRjWho/T/xK4jm1jcoNJq6tVjRlEVDZ9/ZxOZZo5/119XA/
z3f0WTcRmKeb5dMOsJMcZAiD13hwZOdBh1kGqgQ8umhP177LEnU/VIVQveJbU0Re
0XEhHv91TjvtgA4X/I32buf/9oSaUqSKeRySPYK6UyzGL6zUxleZh4eckDfn8EAO
MxADllaTWLhUEOqYvYdW8V85CoA4x3oeNO2tXXv11iS61MfrR9x5NPNKxqIwN1hi
kCi9mpGwkWBw1Zw/GFuhzr+o4mttSnwgjB1BJiWbHC20mKJqXDmiQi5kNG3tVaKv
XMDAYpeqlXmiv8spC+tspmm5ID06hIyFyfgiWjaa1/LOPbrgr7u8khKid2RyxW06
D2fTWsQ88dwXlGtuiI91PcyG77zfWax2Nqk5YEhfcaQKsod3/t0gwNY2WYJWk7/R
rIhvdbqPBQlCaqPc3OGuQLBbEJLMBqngAxfrJpbpL+rHacmaVlVLhfG4jntUyXvT
Hj9rRvi2gznQc096qv5xktXHHykET6rGnfnv/fqGAfmBKv6GmgU8rtVjK3KVScQA
0KV1L6zh/f4dPGpxA//10BfRIvbHtCz6rFpzYRTJ+vUtzy91HPao9enHPUQeewoV
ZwuqXdqiWTffqJZG79gO3jYlMEkVWqwk0pD89m/IgzHJ62geRVo937f2H1LDCOQZ
SZBsf7BgkNLUvkP9FzFWru41TRzkvpZpQJdfPHtTDBoMc7zBHED9JPWLZX/apVZt
45O26ETbQB7VOj17D80rtM/+DGOc+2Lbo8pV7j0tTirIfi6KgJDa/SUy5BnzXxoy
IewM+H6JSU7IEbvfbPIDMLQKN4h9WHRPmnNcoQzEdQuMY8HgWFp18VWWd9Y+Spvf
UimbfD3WVzEluEJohwabYHUioWcKQhkCYgPiihe0rXxoAPDX16qZbFXju1ckh3fg
+YEJ5NdcWws2PiziC/QTTI5MVGUrX6qhsEqOCvvH+EC3o/TSaEG42tOw5sXjFJA7
jAeNT9nW8A9ag9xzJQJ0b1R33aTseh4zSfccOJs9D5hyhh2KSShE9RWuhh75E2l/
FnbsK3D0ZZxGavOlKHoJm7Bzl6ptU2MDJ3AN2TKe4NNZjogM656PbXz6Folm3hG0
fgYurXj68M4xg99VCUW5Ylh9U/jLRbJMLy7/1l/erz8cGC92Ac+QNXqYZGW+gIaS
//uP3Uew2G6yYjsvwOGcpiulQQgGZzK2Gomq8LD7IDSMF7oQ7XiPlDFYvbx4x8V/
V637OJcQyIm/fLKmbKW3MbQR8l4CvOS3QNj9MoK4p4AHbXgdiOcSpBTS509EgH6J
rN86KbfBltRiYsj9whxPyOFKSdA43KMC8y8QYFQ2KhtPMKaSmfO7rBg0Nov8DT4w
lKL1gHHuGA+Jhy5Cw+UN7LEG8tOj1t0OBWImbDevdEujNyPyMIEIuI9MaDbKYn3y
6D87uruoxJw77OKyo3Zxwcv26rj9c8AirCiZNe9DicUh9wbCYTJInKPyseOlGyAh
kS+Wj5IlyQ4I+j7qSbrlJCy7wEAUy7zVdkSMRlQEaZhz1d+Xr+W1HQZZfF1Ik43Y
bEP7/hTngVRut80Bh6mDrye57uKCO+/2ZJ9vMvaXSbxHwzlU1xkexvDWYPHp3ErF
ouVfuWg26xzbfizYNtSs37hLsyjQg2pGXc/j5N4qqQ4IhtbnoSSYrE3PBONdk2qL
ztTuEAlQ24IfEjs9+M+FStEB7ThsIEtd0EO0AUxmmgaAQEpdRAN09ZGMZB1kS9Ve
i2vXeoukP0cmXS2Gyutb+q3b2zmHA9MoRTyWOZbibdEP9xIPuqYV9QnNq0taG+vF
fppenWEXIEHqqpXci4aAU28iBqnLIOSl9VpqSM+AiZ29Yf/4PVj1dWPZDE4Jdtun
fyWh7fqSwE82kdd2yGd7YPx7zIEcNY2YrRov5Ji5f7WdiEENsv3Hxj7gjEpoENoN
BGPOAVsyTd7u7FlSkTjRGLjEFMteL8upZXlIv4crxpwp0z+YCTSva+W5F2kLzeLR
60Hsw7S6l1/Om/jRSJF3Qjr3zMEZPHyh32w70UMmE0mocOfDSVgJEC0Hd6a4/lfF
jSTdYSx7+vsiCQzqz/P6kLhQNJuRDYkeRFAeQ9a/bbU/T1eCztGrdI9wI01Vnkeq
279FARhUWj6VKkHUrI52A/hDFEdYPeC2XQedgQyrsEAH7FU/QQFee1a9VAvX7L+L
kXh9Gzdtn6lM8MHFRM56F17qg69nP79OgzfXxi1SpT3WXVEjBAd5b2BwyXGoQ8sG
Ix+Vl00/A2FRnTkmanpvM9cTT3FzfDxIBatukki4/vzjCROtUuUqZtAS6yq+e88s
ZtTKvYkU+r0TUaGGX0NP2JyyaiJ5aOJ6eeOw7sjuaWdI8oX9bc1b67Q+QABY/Glw
B+SHrAdWzw5idVdBi8WHXrXZ6FKDTWVmBnwR8tziG2mGR3S6ej59xfqW5SO2dbU5
O90m/zVgoE8BvpnZZHL+0QqbqlYMMnuTUSGj1tqbdOksC+phxJHfY0PxwEDlMmXI
e3dBh9gLPQogfIWya3w/sB6UezQFKwHBv/bwYscvl4j+3KmmLsQUsojFHLet8STn
FN7UD0e7aqWiRia1tRX9C1A6ZDd8/j94TqRN0vyPCO2/5QCP77tcYpx/kH6Y86vU
gt2+wlfUT7PL4o1gOd+Vw4qZGHzTkfKbRfulZSNwUYA2Cg2D+TVhGOSsc7XExDS7
fEmpEy/RWXIH7ThzoYML2G/YMATj6I3GOdD5trpO3uU5rISLGAnFU1INzpGD8Uxb
DBRtGrGGkc4q+6vT0lUP2Lr62jQ0AI87ZA6A4OYSH8n2hXYtQHwXYSDFCiQjqxGP
6Ygy447UOajmTbXnMX/KZTWV/MCI3MZAtdbEbxPisyUoA7UbMGo0x7AUn11biHeX
NYOytNQd0sfb9555zVeA2EdeiMGUXtgAZRTYJYhxoVw+NPoXmDm9wvS6R/WkoQkz
1hcDIg0Mo5D7YhBdmSmTqx2m1aqk149+uW/R/ilYOS8nUy04UkUz76+eQubvkLyY
Sm4R/KJ2dE/u4bZDjUBL42TVfKLNRM9OfArYCm7HBIqLzsuRCij40M4+vVsesGUP
XCtTyTbbxbi9GqWVtzr1huy2y5JzcFieZ1ngCtR9dLW25Qkn1MjEKsXHOT+WDUyV
PfGZPcIqhCh20rhxAYHGgiGPGPFZUVTAU9hIM0g8V+HZuQKKZbHxhgfVC0Mbd3QS
Bx4v2hX0zrTkUXoZ78yjIfj6ihJkdFnaLRSFxsCmQQOp/l6/vonKa33xtpDI31tE
1eJg/HKSkAnru/7mYkt0xI3sEbHe7MkUW1DeAek6XReCsbWfnZD9CnFrrblcxEdx
/lhwBR0yoQvz6sskSkmbAFwGU9w+NHOHwUZbUkZOfITBYOappsqa0HUfM/he4KBP
O6YvjL+NzgOoPM3HT/kG7lpXmJgVNCpgozujvS/RoNr+i1ztH8bj9hwhTYyafcdo
mM7ximyHnQ/IS3MBQDPGNc1Bs+cuCueCDEM6EXTxEM80/ZiIJvAHgCOyltldIV3+
NFFG8o45VcureID2kXSsjqjBRkzDAr6b07EW/vqe8wtwI8BO0FgUlB9ui0uKSMkT
8RmjGraSxz4XH8XmBeLdIGRVTYaSIOUVoigTImCRGrQv/wNS07htkG01Ei8dHPjF
g74t77MKsakonAyHdrQ60lEm3lWKVfrgtN8GUWVDNSWM6BVtLlnWJXKTqQZJ4sCB
B/H75/ZGhzeuhCULxOqacYMKtZIEfAx6oYUXuMQUavNFXpS9J3VvmmPAf3Il4s1n
lElQZy6EtNfUx2JXK5wSKlPUEMgxpwz19bPCsXYasn3uFZcW0gPExvdkBEawV5yi
GzBW1DJnUTBzTxcTDd5jpzqtx5DJxfzt9fyz2+jzQ2LxfHPx7diZu4VfmxvBG7Rk
hxLgUqB1E0nXH7ivZtDPx1vQK2DbuRbNZMnELPLi8jFV0bVOGWuxzoScq31apfe+
aJZG6DFyynBAFf4D18Mxglkr9oQQIQ0ozKas/lKRr94Y04g09tAOzYXU2V0e847C
KxchPMoIXJeAfRCAEMIXLZHniX0MfvIhOwXJyKbVcpT6vl/LBHbqjQo3U9enI3NJ
lML3ZilPnNvmumIvJ+Idv7HEzJYTdLinAOkCyUnaw+Q2nor1g7hJbbXyaNLOV1Ds
+lu76Fef8TZ9ZvHpbzLpC6qYKSsHM3JpdoJdEEMo2xz+DkCkkho7OwSj7WI4eWEB
mjpyXsj3ulux4BnV4ci7Kv4qp/A8bijBDe4VOGGSFBOB85eQg9qFXOQIwS7/DDlU
9J2vA8+eQYRueYunxyHWDlZsqlEo+W8a5wOVCKlLprhWgv/3pxNC9lti513Tts0a
xk+YBrz3NCc/CcAv/JV+vkVJ9Zt554XeJY+QnFg1WvGN2oHpqmc23FJu6Z8zI2xP
fB6Ueo4NOJKcAWEIiwjD1HIN2mWknVwl7bBwvklNoKZkIF+NQ+SVxXAqbdgaEWGo
l0dRTPYK8ZCwpEKB/Btb0aTEQbxhOiovlVD3LXF/m7THfWBCKsjQr/EbARVhpTTt
xrZ8yricUMMxauGYI0gBeWdQHvAbaWE/7BV5k7bJBc3iTAzoc0WZiO0bWQeCJ7Om
qPEEJg8H0zxw/a1qBJT7D8eSIp1oceJliV4kteO2IslhLzK/Ov+ymkrhz8Tq+fOJ
PB215YsGF8LkzSQ/3IyxMYVy39e3g/WZqaY/473FNP1NG+KJeBmHxob+6/TSorQg
dp4N23X+lWzotfsx9lkm0KxsTdAsp6BAU+Y1i3gbTqqIkTt91++X5UwjxOUq4eGg
rJCL5i5XjcnoSynH+NfyofqoeOSbv8KSQK3Ynd95XqrW3v9GIywHOgtrbPeZKyJc
SzixCfVJNytWovQAAW4LzfELRLEc+LFWcf8rUV/CWM+2+DdV4TpGvngAPCdjxvNX
zlPwIH6BaQ+nIzZr8UBa3AV4vsZp36diyaC7WEw+IL6qqM67NGfrCM84t8zyzsEv
OqL5o0CFl9hTJLDVOPzfg0zW2SeArFffFEH0bfejRRSMC6rWWtsGFFlwZJplS2Ie
Yx/kVYVMd/4SQxHynGz+mFQfhR51i7DYmeoWp2QYFAzuL/E1VGBLaDXItZYg6739
z83l9y4A9DjG634Ba85RTlyowGBrMWXGF3tT3y0PvIItBdOWbdl50ImswXLGnRhQ
vQDVPvOf9F1bf//KsrrXxdAkIMFKlvDDJYPGXc5NnmXA1lGx9q8/0bpsPATv2q51
fEo45HkvnKD11U6oLm0JEFGwXAEeOYZr6HpwZPZ58BOhotFkgOgK0tw0Wgto5Gjp
kkxe/hxZ4oL2lXqT7Pp8gY/5HRr00CX9KpLHzv0iqEduLyRRKusQO1cS0ESM+sA8
NgvFNWoSHbmlNO3BCYTp8Dka0ATdzs8WgP4y7eDCjngVsCCofJkFnkinWBBh+Tpc
t3gcyptdBng5nJacojZBALONfWTu6qDzR1qFEiCpQ1oIT62+qx/dWYsLlhVN2gkJ
aZ0MTop5g1VzUN3H0yC89I0q70WSr72ciXzas1HiHYsieJnLfS2TVfyiuagxbvL7
9E5tLsX4Hv2ye3eAT7gvwjmGUqhQNMGJICpUh437zrOIJ2IlUs843nv53akT8lSu
iarEdUKfB87vlz1LzATkCAwpMy730dER9URtb+GV+/Flt9F/ld3xHWS21jRWbRMG
FbWaa7rtN81787mInQd9jWQbm3j+GxepB29L24huXQp/tBNUBYAujLTm538vbFdG
5OKfI0O//wrSdAVwZ0whMMbH1MzLVtDv6r0SvFhZYCBmO+fJ5xwEcpZdzxZcfIjS
ufURLD87bYy//Cmrw3virxNp0b/108bksDupNZtClZBwnJH7cpVS7NPkSBfCAoFh
3z1v4M5NYss/ElNwHH599x+vG8cWcZHnw5HL2yVT4PMLgJu/mFhn7lNcPL0ipDAv
ky0vdh1S4Cs+OZbmztvGOXHN7wuwBPHpKqILuFnbMlpylSBhvAx8hJj71BZQAwpL
Ll9ziXjnvjAoglMt0IvxT8Rfv0kPYffVMZrQF7yP4my9N6sT6Om5Zh5fqD5Xb+jv
RYpMKdwYbbPwptOvE9hAimahfZFYTKYM2ozwEFTUQUiBbG+0Bkpv3hkOujv1bDIg
nE36WN4O3kfLqwnVZscQXEEqA60q71Tw0T/0D5wCqZqifzkXo6KLR/V/fqQ8EWad
K7UdC2prMpsgDunD4Oz1ICJTPENeIGtVJI1r7fsQvZwc5wFHUDs6OpuTGTTCM15P
cbb6fUPcKPdwhWj6o4M1I8GRE8RA/R1AYXiULoUeYd1ewGSbmgG5NWkcmxulCUL9
8HqS3cRNR77cCR1VAzROKLli1LCVp3beM8up9TpdUnU7OQ8u+oCAdZPynNtkNaAH
9JQn86dRIM4gnk3Z+9SIR6UPNi7hXAn4eUydEahKiUonYd21MuaQRo7NzHgNoRDm
6SoMYRGUUd8sJUU/q38S0zdaVE6SVsfpsJMvstoBMIuYloz5qSPLeyusccLtC8Tm
d4BOClyzoCbp3+DnEZm4rHmKQ++pxRaT3JNDeAvVqUjitZsEMXg2wwUg3ZOv3rcr
a6uH0ZoTUcFrZDviAQxDudrlToJVCN4C5SmyWuaBMLsuCi05w1KWWJivkQzYmw31
3RospN/LSa9Q232R5/FNtIDRd8aDW1n7cTRREnzXGGPp9hFMd8km8k6y605ErLNm
hwZ6qJ1lXQAFU4frbKn8z4WHfC0a39KxXwBtKmm1vqr7YT+YG4YQTJxvtIWcMTzH
ZSDNhCcOgiZseqVqaZ62h2aQhGQWHO2QNJ5e0+8QqXMuMpxFaGnS00V64LEU3KNU
g1tIuT5LWNk3KycNTPZ+xSh29zjG54Mj8VZykhTQo9dNPSN6ogMW50UlkcniOPNQ
yItbvvwcnSkBxRBzcDLW/v6TrwUWjp/Sg7ZMnM+FTDHmEiwUeqjvcFEjsr7S5C7i
msrWyh5lJc0iQxIsn260elGETfzZliNBbDM1+miqOIVzOKmrjdGhdyFmA2ebsFFf
mciTuH+KJxsk1N3ZOZfRxvcgbXh7xooAgajQbvLVll9o1i4pCBJ8SZNL3bY19Tgz
kn/NgW8w6wCEubmp+tUygZxF6I4qD6QhWxfyi03TDBETD2brFobw3oyXBfRLYDyn
8XoWyVBB11I8gYs5GyqAYT6/QN9j7sFb1EczBTL/wK73G6ccScItKpm2pnm1/XfB
5DMrzjCLMBjFnHSrrzzPz3MMh3A9suterW1LMbirnBoQmlePkaePtzFLqQc9m5Jd
ECgrrlwuTZMMd2QNhGrqcKRsVyJ6CTgdO1FFWWkc1UMabOjOWFNegArMTy5d5h+j
+zeqcllcwoOxB0Qhjv+Dhkqfd1QHr5cuoJ3a3TTjFS5Q3hyyQkdpYFl1ogDmkbyI
p5JFsf04Y01Cxx9SIdKjk89DnDIc8TWoXltYOEik4PTJ67nqNJv0vP4ZfbFGvN3e
wqECGRavsT4xRsCMwAvCDRotzdTeKG9gpDT219DaaL8ORvva22Dek8yheRPd5kJW
rGcAdjxVuF3hCttdNIJmo84VWZ+p4kFlFSchTW1twv/xmBo3bT/q1x9xXXQ7o2zg
15CTrqsYHGswZDNmObU2Icy4mU8OFuwnirRYoJZIOVtHkULGPMxOGmYdZRWUD/zf
9IyLs4YUqOyMIYIPToraawN3poDBwIUyS6uhbqaiiqlzH523Rd2cqnDh2L/TuIQB
uPyxIn6IxDoneieHK4BH4wln94eYjriGdyG4svCI0Ynd4l7Uh6SWSt3XI9KA2uGp
BRuR4Jz3X7krdZ26BfcoyNb79mUvTMrxnv0GxzPtVhOrqgiAmc3xasBU5ld0VFQY
U7s5K3jUDIRFTe4p46X7Ixj7D/tSGi9zLx6szsVdE8dy4TEtyfEG7oj2m1BrQ5xk
lQGqZil0/hUoqkMMzMf/XE7qc1rA307HXx6J8ncaNn/jQISwc4oW1QsNUFXoL0oZ
p+/3k++47bHgXsEzAH2d+yE6bwJblWYVy2UG/ayZ4YNW17ThYggr5IrIMmgOkxll
UNwSf5QlAjtdwkoK1o0T4lprMf9oi+GagLiXytKk6JZJkFv7f6T8qRxEafBsbIG8
COREC5dVieiESKnOo1geyndxDjKji01dbCb/kWNQm+zhiCqEyuYYxZi7uX4oayUs
f/OZr928oDWZnq4A8+iKkac6YRdEq64hnRZSUdU2Bwc2i33XD1/bI8W5JRIuXH6i
9EPv4Wk/jCfm88BzrIQNlZ+3Acnv6TmF9xtNH6zmqAQYB/xI5nNI+uh1Ds6jzYFG
DlwKgss+RM/7Zqkxd3tRfeKIZs6v1nk9kbpBrtNpZBaUwGLu0SMbyN/xWA/zUGUp
Lt0r22vIftl0koCnbOT5PXnW7wuQbcXLLsYt26Mc2suo9ANNzjubbos0JBlrMHKx
JYkrGDO8GkmKrVnZy2QKFzotIrgvFEDiteJ5huCgcAicQc41nPUfYvitroJ1/vMJ
nAAbW1dwScSyer10gke/LaWVx3ybheyJBnSzTc0OLYU+U4gOMxiiAdkLZUWtr5YX
i9/XF/mE+W59bRGuxpEbg9i9brfT7TV8378y4nRPFeu/EIncuavZ1lpTPj//HrmT
L8bT91KeKEYyVL3Sy7pYjj554AjX71/MUoDn1v6055pFf+ZvVJuvwv9bEHWV1n2b
dZKtalUN0sJRsj3fYYaNMucocjkoHfyJJnUmsgk3nfznLJ2n+x0F2RjyF6khbfRX
l3LOTWjHLk68Uv24knrkjcMSY+bbzGDPZpBzwCst1+4VgaZYfuVLKmqzvQBRyLxl
op5ydrh85zN4ZVZ0n1kpnAM5pkHy6GkSPcutXchT0GrUClRM0QmPPj+FhVSK6Axu
oasvIQVSHw7XcJuqB32RtCYBIdDb8P3HIHwrP6g+OjsoGuBnehdN7XIfjvYaZkSo
E5bPf7tNBkxXmIDK9IOsXOGXgnw4dt1ZNwx644v4+zWrved28e0wxidlaXWRuy4T
aQffg/NCph3ubUWqFFiVz0eE4x3oEIPNclxlNLSE0bPbO6D9su4lgJZ8PNotfb3Y
bXcGeuFuwuCJibSHy4lrRcWqE0K7+txb+g7IDx6P18Pdxt492GTVdD0jftrB3E8w
UrC+RG1bzNUJTJxyHSG3NdI6+myarOjSg3TqohJPi08AvOh4UgNj1IU2qWB4T6aS
tdQ1JFKTWTtz02DHWKKwrSZE3O08jLAUEu9Kjtr5hbww4eqFH49XEwegXV6+gKKx
B3CKevVPwApvudz715pzIe6W5sQWysaTGETSiVqkuKK3npSKQWOlGhdwjG2CJreZ
L3ZyZsByQCxf6E3aQgf27Ftc0Ibfal9V9KPYiRSwaT/ZEhO3hp3S8cq3YS8ZICyJ
6toVRezosmOG9KgoNMMf12aacNEYkJebpWaUmD5v2xR2raI7Rmb4MK/ETA28jQEq
wKvPsBsxNARiJKyDY8YdvjrGZqYGWF4d/WEUlf/8Bp5ly7VNGCceFR4Ig/AxQL6z
TIJkqzUeN33WVXECvNXpfs7khXy8txljBX/2ZreNlNnQTSf3015fKYkeIfTE9rf4
ZdycUHP6/4VcP1bW27UaNbdsPJo8hpnPHK31TmnnxuTuq31NxHKZORO+1HEbzJRb
ilEGHnFjTvUEplTg/Buqft56rTK9rpTihsgVlZ4W12+p0ic2qzEHfmeXmMoxkGII
OB3hBV5r1PXk3wpE/BnYtkhgb4xYamFGW+FbeiYMaRUZDP7cDeGMj/wcSlH8hfhq
hzRZ7yKsUHg1aaUHyWq3bkF02oSws5SaykakWmf2R/dGd2tFH2vkaJNDMIy1Ei6Z
E47egEK7in9gTNBdgptdoRgqVdsUvN+FwxaXRxA4ij2Sc8gxfvwx5EryzlaCtAkU
E4cijFQLFdn55o3GipbzKZTLzyEmBCEMU971v1KWuZvO6tFTZWgSSJQF3OoWv9Tr
Yzk1HrYRgHemE6Hd8aAxAc6SnfssMV04lmL8n3A0X9u8VTyTcDshpmOPvOdL0ucf
lkPoBmYGRcKdwo6UZOqR4gAMxCLs98Pk/2Ee6RBIgX5SvujmgCiRNZD8+xGLW02Z
Z2NbmPaLasZxLmBdnv+58H9gpMnIGO3qF6nr1YFQdVTQNqZ4INjgYn3L9P52HPfc
1SBC3tXaI4+ENp2OlRN1DtOrrijFwSxUafhX/n3+cedyS5VB4CE0v/ECxEjf+C+K
Igl2CdatN7jSs8lYOEf6b6zNDeBS7mMRMkBL94hw4qkJ9YDPqJd3B+itLMEDXfvS
mepcAR7tDw++tlO6dhmlERUwsOg+9NleHL1H7PHVFQFuB1htJ5elFaXQpuT0tvwO
wyjChH+RRyvCdjUPoVtgPJLUgoKy+i2Xl/2PdZrCcx0Fl6JVGMdJOXGJ+WR1UNEs
bPvTiSdZCPA/kcwTEhcRtq3gvy4WLbW5dOu6By03M4SDTacCFHqEnSpVLcj0ZB4o
/hg9fPPSnsj5iKHdl6yhb7QL3Ds0gBkewALqt/DRJNIFHxanwrBayDL6U+EtF1Wm
pQ7zCYxRqg2qia+uZ+eiQhprD4X7ekaA5HT+K288WwGrNjEtiTsdb3+tpuGf1pPj
l7aDF1flUYMJwOUgOy+OI9I8i72z9x+MAph1HnPjl3BkONkVCvFHK/8UpX92QNj7
g7e6p5FL88G+0kNerPrq/1wVq5013TiJmC90SqS/eAvC5s4r2KtXTgjg2lhqeCnD
Dvl+nbIMJNP308Smzg1QRkhpZETbcNqLv6B47wDm5H0pvhx1HMA6oswpv8Fg6y/L
7SHosHT2DgCUw9uyqRyj8oshn23RLARLj6WTtyCySci5u/0n8r9+GW1KWSvXFY3I
X1I0cgHAX9ogBcZ055/cSkXdOeKuElTCUMnrnHLAr04bYu6nGRyi1miiv9kXoGBf
e4FYXn9jidr4TR0SV7zNHyhNIssQ2wgAnfjeM67aH3Gmav7mYvuRv0gpjfBWcH5j
26QbzQbOl+jR7xl406KjsXM9OTzbC99QNfwhX0E6es6+nYiwrQOdjVOuJ92Eptgl
GOs4E8Wz+N2wkFy1+FqI547pGR9D2MYEJQ8Z0EdfWtZrACYijZao60ve61z/XAal
T/M4Ff57JYP3LvsHmcBTtdL+W26wMRkmvB5pjlE9aqtxDhjG45quQzW2QRdzz9cI
DwJjo8eNZqKItR3BCS4jxP4aKWk+UmdGvL09KvwnhEJKMGGqMWlhxm0uTT8wNUae
d8aGqV6z32MC5fA9IewvT6cFEvEkwl2BDle9a9szSAfd971NIcST0e+4ch1zTzuj
Xi4ueYSWaQIgBRWnXJ9ZNfKxWajFt8KSYjOPhQjLI6wVA5uFbY6K7KENUC+ak5Z9
qwVD1BcnuEmQj+YQw4nqHlJYutONNLDhbGe02sCoCpV6x0QvInfmbDpkCxejD+Ey
87tBjTQYSOjqviztnU2upubi9Fn+LlRXimNv5x+FFWZfZEpi3qoDxmMxA3N4rRyB
Xsj0SMDQqNPWr2mGl2QAdH1JdrRi8iRXLdX01h1VpM5O8678DGw0RRzVpTwMeZM5
y5r2Z2wqCviTeXhhnBSDna9gn0lUPzYf5W7wBBsTmEN1QfQbdr28lhiLzpOtcG4C
WUw6w+tEgS4mS75utPnRIw93f/erIVZ6lk5OAC2/oFa6Zy8RzVMSnFsWj114qktc
B9mji9LoctQmMlp/05Gh3cci6tJpT+BGGJr1whMHMg4yjDbWQZA6siPMzLXHZoYO
eShewJNaA7xOZL3Jy9tcizYSpOTZJ+1fer51sB6jpT/0YNUZukP0Ksa+Zm1ZKWaW
uXP93qkgdoqDQX47cxHVFCGeXHuzcTA0eKqaktRZ+z7jTfjqTgXqtBQLc8ePpAeL
8V9u2jNNm6w3HzTn8mFIZ1MM2YQQkVC0l6coSZCpncmCY4k4PVgs/yPHqyJ6lBJe
F4YHUuQ7EeJEZflmsdXAg7GGpWsqxNnqis9du4L4B2wXJhk0HPIcpVirh9ni8x4I
M2L04gD9YIbX7y7q+2/dn7NRawJaexMlxQFGr2aQ/Yr3iIQJsYZ9+rJk3mUPf/mS
HY7GbG/IvfMSD6a9SAJkbzfydKej18CLMCBWGJSbq0HbfMK6lgknHWQI2ZNIFVqm
Swiz/U6jcfkcczv7woXAZ/w2kAqcxn0dHThn3xIUIO/4dlp7u15me112rYjbYPM5
1HH66+DrRUMuhPnauL/OhHTmM3bw3gKxBVbhtUGeOlnOKbZSUPTbblDvrmx5a2gK
fMS58E03gOd/VdXNwYc7WHPyMo141Agovg+shb8iw2j88EGMvlaSnfzxRPPovlJy
s2MF8XDr5TgZkK7kPalxfzHbacTSJuPauGF0Ks51owhbM++h0A/xHG7CRLzR9Txh
Fx8VA1Dbr9t1KriltMWTNRBLPChKsd5WsvWrdEW9z4e6mjhT1NtzTjw0pjxWnc29
heFqICJIt+1obmONPfwyT2gXRHIXS04SwKbYk+f3KSB0puGS+ekYdYUckkx4gm9t
6EpDw6U98eXUi7523GjVVl8gCveFQ5m8t5uyt63T+oGqleclH1Hv/wibexaAa4Fr
6hl1lFGPooiiR5iTiHwBFYjaXKhXFb54W2dT5mrljKY9K9qP857qgTeCpAOEJAZM
mpSRMY8xO7qlstYm/zC4Rs2qyQYFaq5GTlFpicnDv+KO29QxPYrvXad3M3R8AT3P
7cCiNe5vnGYrTs/g2xlNqXSjZ/RKR3d+q09IAjI4j/8f4ZqIUlZ7GZtP267r973r
gs1gMzd3ZZ/rAyIquT1t0e8MG+NVyFF0BG+AMxfIYUk28wdq/v6hy4TZARm/z0lf
na9/FyUXRduNeOgBvhX19mhXX8pbfs3wUOntVR+9kiOZ1BcGJSgBw2vBbh+rf0/R
Tt1QfmNZkJjyDZz/O6M/SmJ0u1Bno1PDGrZQxpT7XpEPXJE8xKOFB1m+n+WtxTs1
0cnLl50O94NJ8Vb81Xeh9MFj5NRotEq8pvZjejTpcFqf/bNKdd33EChgIaJXH1zf
lrIGp4I/BxUPq3guuVRUGkoQZM3G5aPGgY0cU90jvC0rt8V6sm24g9B+uV34POSH
/nOacnwD0CEumJ7Ad/vGaHl6Dlyl9zqP1ISENrk8ka3vyBcN1GLVErEthHuoBOp3
TiOmwR7BpzvIVmf7BISezx0+5T5I7g4pa9/JCXXcL+FKs4SLFcE9zhGQejdfcNTH
AaqcepopGNRFmhQLnH/qymrYWycSIgui9C2EPDbqXnGrHpVClI1Ds3wPDQkbRk/C
ZI/Rpu3LmW2ZHQAn1xNKyOmMTG0YSPeZaex57X7yRMmECYNdq0L/dBijR6vcCWwj
uKtRK8mU7qppOzOW2of5dlbSXRjv/8QXj315/kaGhlwa9/x/wzHp0t2XBKYLJCDa
/Mux8ETXh29znNQzpIY/d/5ubzNbvZ9wuhxKAdpLME0+5k28lcPwFCoLwaLJSV3d
AakGiLzFT03Z7B2xV/dF8sIFlfxPboypbmIrcsdItS2estFR+eTAY/5uSdCKsOb1
NtB/G4/gjec4NFTmoZVbEuF1Xco+RoWYcZMGC4zzkDbAPJAOJbc/cFY9oH3mPsSV
pnSCZZ5PgegCg+4lqWVzCLCiyhfDa4O9yRSeVy4x+z+NOxi7Puwdill5V9uL2I32
BZgGbLS3MjJDUSfQV911KiovAohVMMbIYThFq4xUKV2oWsSnKrBXF58HdyBXmlbV
JVCgfaJXGSDVe5oGv4ZkJsahfC08rsLYgqZLDXjp2KRpcKJaHZmh1o9YX8gHV6NR
DLl9Q5u+HTl8rzhzzi/rfgaOr1nRIIZC3kV0cUv4JdjcZWC0JKS9DE0yuQfLcuFa
lVBzffLJG33W5iFKUIW1wgIcVD++kmDDqHIhGTPM4E7B762UMAslExbBgZH1lsVb
u7HUiQJ+2sYJ/QIvfnckagDzbmmZSObKOvynvDxks9FVe+IQHsH/w7ConoSHuukC
S4v8Y/Woup6aD/+ZbZB8Yvp4HVqRFb9HuDnBe63NPYfKdRK+sTPstHPRKMQM8eEU
tDHpBoYsJnFA0/pqALg+uozWgD0DfvjXW03zq6KC9N1accmURZeCKwsR7wh70DXc
pAxfeUPLMyBkSDHiF2FOF2O/FFA+rQI9AKBJCgfX7YpZz3gAmlWNO+njK8RDrvy4
46qGae3rgbFoX1JqU+zo+hjh1BXu/8OKaGOJdbJ6KlemMOVcYg5tYCZ2IdJ9udRO
K70JlAMVtiMtb+tNHMAdNyf3007gwC84yXKEpwEjLdwBHVmH6yCih81QU9GyvjgV
dczB3MQM23x3bu74e0fN8Se4mSVcpnF+Z+On8HDXJwK1E3Pe62oVqG1zgcTvgDMX
6bXoqsox1domMyhwptL4iiL/j3CF+wwyb++3fjVPfEvvuMuL34MxcS0TT1MOJ5HO
X2T1xkZPtannU50CGnIsnu4lws5ecGhc66j5B8g+3jPI2fIUh8s44IxrQQH+u6d9
1tCyFeiMIsMEz7n67UZSa9OAwYwRMbEAbNphr5LdcWkMVRW+b7/sgCeHISLE5mdT
Gsgz0MTq8uzhEQV/4cDZ23wFGTGhBnXrJQ9pjOouc3XmePVvlsr4JO4+Hs5KulFP
FjG7tWxyflQk0cVHTNMd02wsw/O+AJPCriGzWQ1Y0RRqHcolcqMaLTIyQQTdVNn9
1ZkkCz0GJfDI+e1Rsq8IIt+gD4hq6DJ6xN/TULkkoGV2AT8zVWi50MeDuLJ9WIZo
e9aGfv4rCdGzCWIjw2dJvNG2yg4VWwmCMeOaM+HTJ5EGh8BMBGx2+kmUstHlm2SF
hV5lpvFDzbBHbJih08LERXxKZ4zPgNZr1pF6PBi4+Nz9/Glq5LrGukDPdaIeDAL6
6u7jjn19PqZUHH6bUAbzXxrAgocaKpkfUv8eCKAC+8dGLcsraTdyk9M/qlCmGvqn
/E+vZRGs4mclDBa4bXijsZtN5dH3Nq95OLZDnRwKsbZnx2MqhGplaDgc9Z683NxD
DFMJanaAybBIOCv/9H7tgJybal+I0MTTEizs1wvY8D/m39fOkKU2oHfZcDYAYJsP
tUSpKnGBQZisGdIeBoqUTS0L11luJMTIojeuNuBZDySU20o5P6vv61NRsTsQf3uF
gnieUpuemrMTIG+XBHTaGIaGW6qJBA+idYpzz9AO9dSVR5Zu4m/+wEnpFb7a9aTF
GburjwpK/ICbfrkjPAHL0bsGKN+eU+fND41IlUSk7K6IgwUe9xeQQLt7RDb3lCvL
UMzezTnTUd3SEqpBzSytp4K49BPGMgqeeiZYt19iryE139NezEpN90YAel7eUhPV
FfGyq5/u7C55S2oF+soHB/iUXcKC/F/EkVzK78jBxS91GJjGI8EjKryRZ0nKtybB
erDwZN04Hw0gKN0wf+e3l7sXMJSJ5Y0P2Z0AwZi9oAwmeJ90s21UfS1/P3S58Kqn
F7eOZNhVWx8hMvazWX5fWI+CX+Z6Gw3ppEorWMV7iheV7WK9d+0yG/221gZ2LZO7
HkOhV/uXoBdFqH705YZpwPgF9VNiApKzbdXeR0p31sl8rluovTD9itrsQLkQt861
5ZZHNEt0tsDoTfI/5aAB0n+N0wdzcpOoXk58z+3yEDB7QVhitV5qvPGQpRAJuNQd
Due05F7wJme0rnN4xF78Eph6S9xRrzcqfOwUiJAls+vXaQwAdKFh9dAB9cLPMCun
WeEBzEWYmDOkcgcdzRYf4Oidoo43BphFGFsOFHMieRNJMly/xNVXiZ9NP6pIWnLR
RMSU+lDi/jG2JXdfwsIjavswy+aVK/NX63NGfbLeN2tm8XccO27Y9ehpewB2/QRh
Q2RJ/EmSDMZO/3WnwAXP+/ovV5yQ1WuYe1ljPiP8dTMaERJuyiG/xMZLm0ULww7I
d8UgZ3/li/aTXPuFpDOPQD5mSalpb3J1GZD70w7e4kEZ7Q7tV4BcPecX6MqskSVt
ApsWgM3HfXoOYIG0AmLCwV0hlIFOxKftgebCLRo675cbw7HpXt9zsNsZOItal8pr
97g+PlEXplI+3tUrzOs6q52gGNynQCrrIXoIRsmpTWsQ7TSOHfvOsPMTPj/geUzq
x0noDvSWJ4b7OAICu8GDtEiChB0vm108nmuPsf/mwFse63eQf4BNPdY/81ODJfYg
BKYH/hC85xaUEObDQGMSL7v4O/+dDl+wQHJ3YnnLoDhLAx4eSfqnosrCk5JteOkC
SNLRtsb6Fz03cwz4w3VEU2HzA+Jelfo2wpUPj0iGMZ8uNacfHLttzKIn70d3Wk3I
t5bWblrN5CM41XnLM9wiz2fWRTMFYRh5OQIxwU10c8MzOmQPm6UBst+gnrnZ9YG5
wKYHQaessykJjqFMt7cVKSuLpEqJiE0MGjl9X3Iq2oYtSNMzx38yeI0Nj2vC1DiI
al+MvTC/yMA7NZ1UIdd+ILFiiYIj5xgqj5S4k5ef8GX3OXtVYRySQXffYWBOa4ZD
pQ8eSwRW7H8kt16aAmybyya5Lzf/n4SlVdhszm1LYvSdmWZJLzldB1/qs7HC4zsK
wZbJqH3HiI29pjAlt6VdHzP5TVpyZH/7aRMKHkHn7aOSpkLDZaqdrzzqbsnO4Cup
6BA2iiWzK2T6AMhlo7P5rOMjd15bUjxloVqJOMxeQqwua6MFt35jYdxTubr3s47B
GKJOxR+/YM5Sij6r4IdBJgzwPxMFc7zu5c9M0+S6ajWii8joKHjmkvVMCG2Nmk/l
QH8A/fLsnN0JPP0sMMmuPbi3AUTw4Erb417XeknoCWfJMI9mLrjxO33UlsUK18pG
VpjWq8i2l4Ea9XapzPsI7WG5rtC+wywa8jJ8jKTMxDWZO/uE8Jc7uAlsXXTvrh3k
z8hAwVQKNKJBvJQ5d1nDs54YgtTie9ZyTGvmciBxT+PucjQUXSGvWAajtM7XqVyR
CTiavQdAj2mvZpXuRsTDot4/c38FklRIQPasDjRzUdsLvQHPm8umntAiovxtiVyA
IXBBengrJOZaSnm/5hnn9TYRu3owsYXNzonoIbEDRbyN1xyNZT+8x2tDk/TLKQtn
b2N9Qiv6RnnzvwwLgZKSElPbjNy/yBVcLSgJI2BjfivT+3DA18RMnWNReP5CzmP5
YyRP6cRwT6qN6fY4ZDB7l99jNG0H9MpMgB4syWesdQAqUG5srl/tfKnKVIw/WKX1
t6O+Sa6sybPVGIoxhAc5erYxDhK/tcCq/A6fl47vK0VOPf+vfaBjTnXCYwCHSsqg
QYReXuY5yuZ/saAceqyLIwGjHOsLqbqTCvMO31MbTHCP3MQ+MPiiW/XDRV1mDIr3
xu6+tQaKoGqkylhYUA3wb15EuvwiW1y/0ldl1UqYSTdxmbyIVd0HLcovQ1DQj511
YeNGTKfTrTCKV8P6cUjmdTyZlI61k+dG6zuN3ZfkzSumXoy8o2vpV46k9/9rphiS
RZAIFcOqL3Zf54/Gl+5uDIZ7eKFaskLtivbUPFG5F8gEENRx5/NM2AXaqUurYQ8O
EFeHMJWUmqqIp455ZVmPMT8kWjaSbrpQdxWwCTK+c4Ds+qyYAofifnIfOJK4i9F6
vTdrtzNCUJXxMtl4+9bGv7FOoXq0KyKnUNYY1Xpd3OTycHIHINJo71LL7PozrBuS
x1Ws9KqV+P85frRordr9csaR1gxFDUDTUnxKPoTsLIexku4mRYacQEqnHRM/nlig
iK6+RdxQjBivxtwB+jHdZj7ni0XmmWgbxoU47Tv/ttri9h4lUh/Cb69yXSF5JmHY
x6Hk2Yuq/ETSUBRO+wxnd57VLs6YMzvspXTyHmBZ0XkbkjAdBfu4F2oO37H3djwM
A+FSBH0ggxdzQKS9S2p7yJK07u1UJEYOdkc8WAyXp9ne2yALGLD2sdw2Mh1eLvuN
oc6p0ob8qtasjjfr8mXLvoZpgYLR3NN0ZSHEoWEfF9HwG4hNHsNKHHH4VPWmue7U
ADQsEEle+FNz3r4EKTV2aX4VflAiOGM309/+sICnyw33yyMRWQ/zIfWyVYqmjnka
WGWy2RBlqH9zlO+w1kAbhBHm6/c8OyQl0XjkSoGUYDJlCaV5pq4aE2A6irv3nihu
hMkEY1wk0YzmW050qdXl7rJZN45a5qee50N18dJxoZCCGnEOihwUmKZEi98uknqO
6oI9yPRNlMtwRSTv4N3UTI4hy0BCyuVBr17cRbGwYTY816/H3aI+zVLuB6ikxUYg
t+ew7uxWH5FP/qc1LSeLCyoLrUdS6TIVp+uH5I2sL4iuIgiTDtFhyHa8pg+vZnOu
TnBMYI+7zqkRDwL4Cn2sLZ4z6/+ft15Z/GGdQN/WjadqAKmCEdYBpf5nF0pUK7u1
xqPwBDRGSsnMsUkD9l9Ieo4/fuJi/HMj01m05VNui6d/P1kMqiKAfADmNeGBmlHG
Y/Io154MNH7AbBP0WALziEGfJvWLRdZsElwuo/LhuYoPHr+JfxauXXGIUeOVwNR4
QGenXph3NQceZis4NzKki6wi+vnLHvqlOq4yO24spj9ye4Ptw38VR09lRcFeFkBT
Ikbb9VfrbmzWsrLejOdpbP3qDyTcP7NwbGik6eYZcDOC17kznzHyrBbtwuyJATPX
tIUx+Uc/lki/2xGWH6Rc8p3lKojEOCc4RzcgYEOFfxXTRPn3mMkn/SWc/gbaW/u7
pAUx8h6lLoZzgVxxVj/g0EflZzNF9RPTtTUI4mI93S8QDd5EvYcjUKzdo3fa6Ujc
Q/uv4OVKr2/kDP5kXNX8nUAS1esGnnSXh3j16exS2YEYVnCQv8HqXyNNr2Jk9xjL
cNxeR1y5ZpQdtW0n9pdWo6mD9cBABmd67k3LW0QsBw+Vztj9y/9Ie1ee3iJteLRw
RW82PR+3/gcncFmNC4Sg8Jq1eFRIVOK6Jj2CbPBUZ4Yb3fyRok0ueutiNs9SpT0X
x4gyZIOZjhL1Z5MwF+NZJTk11dsq6MPMkTn12r+j0H6vam7bwn0dDXaH0yIKn1Qe
pMby1ybd8o+wPS+JDRLw35FvqYpjPKt4yk1X4PnmhymQ5mFdKBl5Aqe7wGr8bcen
ysBxkBhh3Orvy5Zuq48+ztAsplKYKf2qKyzu+S8XBCpve20zbxqtveR/xEOH7GL9
X59Zlgsz7T1qCJRiUSh1vXUhvu+JVW6k4ofBAtkt1OKENR6jLCNR56Rb60Ey5XOK
r/R77wZeLocZdwm/tjqnnNcEx61AX831XxXHCnbLbVNyMBfLr5ebABX8pTAoadTk
sJPrN2IZ6K7iIzCD7V6fo/DdlndCW6104076yDU3LHQCyRnB33+epstJCDtpN8RG
ubKIasq+h8kb9yjZOSme7ZxJkr8+tQBKKO8vWeB62DGWLdPOchdqaY/w12KQM4HE
7WCVIksEwpKPhvvNbZOpZdZWMO23gju3zhCxZFEtrEYwaktrx06G1AE8xKAO7pLv
2WRinz3VOyVZgv8vNgPZ+JysPdMenOydynNsUz+UR1V1hQBfoQg1Z2fT/H7B/5vY
34Sx0OEPJjQu01mP4Zqdo4JsrNtPyA7+C6zj8mBjRTimNuEFzO7hfw3r+mre8LtK
xHehY4ZuhxpRh64LV6LRnbzwEApkaaR8uLBg8MdLxJ7GE7dpxXFA9M1N1VHhjULJ
oBlcZ2+MiueVTHQ1WRUmo4a6F/I/KequxqsRvZztTkQw7PhKUCeo2eQEJPEAdwmt
5yZxG6wWtOVmYUgv6vkY4CsPTuMAsNMTUrHf/igKeGsfqEQ8TY42Gduk3mDNLtIC
Qcwniw1hMMu3FmKl8NUVIZPKIRIzbXj34IU4NR9VVIluCIjsBJVtXXVP6iBuC6/0
nTmiP2djCHxsGavNZKIucnstoUp4Fq7tGuJgOC3pvhK3r+DSOj+Fk8qyf85FQVqg
CIEfhJjBV8DBjcKmQgiL7JdfxAKGkzDS84L411eZdrbtfT1+ugLTrOZqq1vDq9QE
UG6VDyGz6VsQH4BPnv3Jl/xdt3PFLKzBjELghpRVhkTNuJ2Rx6kSos+KwV3sd8ta
8Bl4chT+2R3uvjqNQbK4oyTIiBAMapjmFZqNh7Hozw8gLiqN4XtwkS9plzueiv2h
/jHWHAv9Ta5vsPsEyJpSMasbWAWKRJDs+4B5Jj55pTwTOZ2u9ynjow9iVi8DQzep
dNhTzFNiX0ZvSLSjCCxwIs8E54jOsE6+op24pbga/50VaGfGBEUct9yGgWxxGR2e
Jb9T3TLOKbR6gwgHZGmjslsehL8cxKhou8YT+3gK997dboAz+e+kGJfsaqsr84jc
/dwnodlLkNIspDV7+gbcQyoujWlbSLNt9sC5y84jj9wbDpA6cT0io+YJxIhNnz0T
OPt4vND9Kfpq//CY15vRt3TjY+vEEoYPTTda6VrQofLf0jTqfRPUTTz5H19OCFZw
sYtPCH4049MOpEJ4o1BZcoqtt5SjNDgQEP03c3mVSQ+3+wXbg+jKuA5G2Pz+nmZM
xYZ4B3dbf/iRYYlLSlwQU4kqO4huoAhLd7MR8/dJYQ5RvAkDtDxxQ63sJjZAFz7y
+6qG45rnfvG41N8qLe+SBikn/WAL9PAv8ZmklEb18hKjknBrqzcE0aZJ3+MRhgKx
CSpxZJ5zMFJ0vCYx8WF3xXuJ9qfdMN3nZRUOnR4cOWYHc8K7OkWmyuLAewXnQWMw
w+dSuhgIeAK+YB8du4DjFeRTuDxTOACDigJzyx3Vncgo2+AEsULUoc1waG4lojGS
+P/8RvuZCHOkU3pJMbHnJ2HRIsyk5hnrqS4yMMjlRI4kN6mUnvo6iBfNlrzR5pVP
pDSxpGrtrEOBiQybQpVvittPW5CzZDn9v23LN5OvXzGlb7CCrmYMrCw+NrJSyi75
35CuIRUcfSdk037tlu6Fo8B9fKLwYmXBQtvnZf16femjV2CzTFJOhu206d80JSz6
RcjuHIxqhAY6dxcNc00dtJ8OuE+oEMlxlUiYHos9LlFhbTWwht2mxH37KZ3G5UsP
H3nWTLsQuYRTLDlgUIoE3n4C/QekmyAmO3esu7u+MfrIGRcPGuyWi3U4qhXvUG9D
mSxuD/+qX6t+MN/ENb60QdbT5xOIfieQ95aWLkQ4TruARtkQ6F6SpFNrgl/AeYel
nPg8+lxqbMq0neU0aFuUjaQRnzfwPpHKQSHJgwcT28xMMsW/yglmgy14vCBMemFC
o/SLZ7weRwlTXqZkEPUrh6uA9pcPPccRzqIxxyAtAvU0mJh2SGjwmbHrFLBxS8ft
kpYD5jOEMyIKdSsCmXw8egiKhRDmtb6PFGO0Ho2OanDyFmvxEph5Ad3sBlKK0p3Z
hpdCHoKDOltiXk9AJFgK3JceEjun2nTWQfAzx+eslQEAjhJkP3lOw8TFkM1mUmRF
YqNP3Rn1SDN7B7WTVqOg/nBxMjFFpsN01A7uCVtSZtvTt3QJ4mKgzuOHf0D+Mx14
m4m6u+ffBCqvak6X/GNiqcrbVs/Dmn/W5oxDg448/f5s0mvMIvKlNYmOxfZlPUnO
A33XAT5mNmtrC3bp5bipLMUwweevY3Q9lYJLVswv1+jDejtFUmLOT3RB4qI+GmZS
TS0Ffa+TR2cS4sQRP3DL0UfLRHmyDEEUXE1xG/vFQ+0KLjnpIVT0544hfxVkuEG6
D2MgiIM886olh2KXFwY9BUwxgPA9obr9glAzoigAN81ubfpfix8uh+MSc7ZfIQAt
LlyUPbJbUE2gtBdC2O0zYLSnlpMFDf/WT4zkuk4YhJ7WYQQ35P7fmQt0KpTaYj5c
lrmHmjOL2qdQ38VK22SzixIYrnb4cejKWOjjIhN471uruhi9qxpmTBO5Ky9880zt
CGe8xL0LcB0OJZtjf0wbafxzZWYyHxk+Vx/mX62Y0D4gwBvnpwtGK/PIuRW/1w3g
KMe036unDWAuE3ZlCTKgFs/DsKF/eEmrJq1vUC8i6cvxOLKTMbgJA/iHDl2/6q36
wvFdpkr7ZcY1rsUocekSvq8KSFgmkDNzGIxJdA4S7v9txDW06GhJiyhbCTfJ4dG3
VHYkfBZxA5dnVUQehmN7UbGdje1cE6kUEVqxboOfhDdPUa/ub1PjEfRFjMrn8ovi
nAou+8fNWIhikgSov8rWYjBJ2Ngn0epudOVlHTD3disSguSYa2+nNlATU/Z33hC7
oKGdPctO/Trt9ilY4ima9YLFoaPl+77rriMdVQl6kaxRmwHZOInL5lQphqxg9+LX
pWGH4V5yUhissspNCgnpivE2OrDYbLoTxfTFTd3+bwubSbAhGYMjlNVraPH+tZmC
4ClhYde5u0Ndw76AFSGbYhPoYgYNMPbEYV2OPwICt8vklpO2/BoJcUq7bDCDwvVz
+GEqjK2w9zpnvOZeNf+fhDsWRAI3rPheMZB7/84OqPZqioekQVIea9HJo7LtbYqu
LNebnLjqYXqz+uBs/2DCY3MJQiLFoOcm8Vtub50767IOOn9oFL3XxvaCBObNmOfY
QLTKOBygJ48LgklXlJ0PSv7NBqCw94xrE7GZtYZtisnZCIAY2G1pMKDRxkQqi0ZO
/TZx14PhaWtibvhIGYJrRMqWgSB801WzSZLdwQT2aKKhsCl6a69YJyvaYhUPY46/
3edgP6BmW+RPKsglRlAFu9u3TxoXITdAUx3WRMx+OHXkEpRKLNLjbV5A2g/uYVAn
0zhoxtWNPwJyVOyrnUgmcdruzNdZacT06JB1ElFgie5vtqyhPhgxGTngJCjfwWGS
kKddPJ++Vrp1zschEiKTZNxja9+IdiZp0LiXubEM7svHTjyKnIbXP2GtM9ED0Fce
/9YrRFFuwesxtBwUvI/FH0KYrrbJyb2115xRyhlp/cu2m+wyMUnSl6u0BdoT8AD0
6ATprSelOU2ox9ZKpexHeREtHykJ4E2kArwXpLHMUn/MGZ7G/+DGkb+a2265TjL8
D7FY6vPIoWJ6hu6SU099vC76cyjZLRNN7s1tPe6HP0CMM/Cu0FgL4Dxlu5YxFf/7
hqZdxAZT7w9lda4s+r4G3GnNjzY5sDYepfhNdbeHpXvNxnPlZMH/IQKM0V0n5xvq
HLdRgb9RASXVBwsT0BUVfb7BPe4+Mhz5BCfuumj1ITTlzk+OA7jVtGhbEyLMjv5I
AnB0fzMiNyfgMSJhAYi3+oCXJV0noQJzZbZAboaeJZX5LkLXAQc2Iutzc8MLpePC
oAJL4BvbZ0lC1+hzvfE1ju4T3aErg9MOe31SaVckT09sdR4sbWduK7uXFS+NE6XB
DTeVx9j6/vPJWd8aSBmIt2aR9iln9xIHtQRunSz1AjvnWOvpNGMY3GTzllxRmGTH
lmFW7YAuXlkYlf9wb3ikKQdloFpHwdEjEzXu/bj53oPDmWypxXAXydcb8ui63Q6G
hJtHGoYVODUhDOO5B5skAxtVRR1r8NC9moHyJjDaRWBzAIHuHDC89W0GKKbLCoZq
cXZYl7ENgoSr0Z2Ry3ytpFPkAjIBt8dILkL/2dJBun1gYHg32iB2Oy3Uj5IW5PR0
GAHY3ii6ckTNqfimo49fM7fUDHPpfJGL0dIi7ke36iRJTCofQuHL8vUUkjEL+5gC
uhiWcC+wi/gmXAOL0Jx4bwgIpnPCGCYUWmuOTiCOmGy218P7/83+HvLbPeieRgZO
/P/5jusXPeSbA2Au8TiHDHlykAnLuJ+dDn4CyFzhUG+x0T+gkoQbrLI5sCCDYXU9
snF/7/J5sbv6nhetbc3tNU50LAhqJl6z9/tcmpfL0TjlsvDEfYkDOEdLFPZzc2mL
X9oy7w7YIeZRcIj/LjrdFPr1Yv++jM4etKJg6sOu+AUcrsmhkYAjtmqBngZPcOUt
iOgkmA1lpJiMOMN8gFQ3zujadNM2s06cGuVYhBh2TCATY8JimD1m2sthY/1nY0JG
cE7Sz/mOKWIGgtO7NjZpPdq2jZdXuDZ3QKxO+ajtkSRGAEFezizhMKcqrVtZLsbC
h2fG7nw++r3l+QG0YUmXseXL3Swh4s3qPppaPUZ6Grkhh6T6/QpL2DXUDYr4/z3k
yg79I2AcFtlLrEwWy3759VYy4H/cZ7W6/4TlvLZNLR+iGN+MxXNacohbrbZtRBIu
Ttds1FqQ2XcJWhoRx3rihIpIAka9jHHhv6a2gWv2DHlSad+Y2ueMmUuUuU8gdyOc
RsTFhmGY1pWT8kFNL4THqiD1x2DakWFc6Tl3MSaqFeF7HY7DDp8E9IgtLSL5dElk
DArQ8bAQqF6thDYdfOusHWkUXflam++SohCGfFgWCpdLKKEglEYfB1+F3yjlBcPj
olT3XAregdH74ibyGtePbHjOi7S1YckDbF3MteG/lua40wpphdJLJ+xI9ddP/0qP
LylskBVbxS4BUzOXLHx2Qr/vKpTdUx5fiZ3CGrZbWVAkrS5Tp1i67zSXPgyy8kBm
fxunO8EE4+Sq6JoXwbBIIF6P1nLW3NxVBKd7/x21TfCQSuNf8ooUgABqP64w6U/a
V0STROTRf5UFa3qHg/X9tRRx8CHWQ1hXvzLt2sTQbajZh3q3ldsqiAVzc5Aw/Bog
6t9FUOwRPz9HuJMFmJhSbQ1kIjmt5YcEUv16lAGPcgu1s8ZXdhuXIrLNfHT1gZKs
kbnnVhaMcLVOtdQN+kGTQZZSEFwWuVC6JhHef2aXpGPVaJ8AeQmcxMCR4xIzQWYs
90Lw2bJO6ssoICuugZ7zashyYN5MyV3OdlOM7Kue1AJHdsGVIsNVELQBVohlypZm
cJ7yhT04s2jtqmTqx/5xixPl+LFTLyjkm7Q7udB2eH5NQpPEs1/mFZTGlAPN/mCK
+D9pXKyBn6ZLTmd0NESe/LcFfUadzGgUgWkfX0Hku9DydPcaJhB2fK7z6/P/G15l
uVe2v/3If33yHdI6KhhmJwwrMv4u+Vp49A5399pNXFHPzo71ThdZPQ3lcg6KAceM
1FtZ21iJIqrps1seWzJuLfqB2X79jq3ucB5T0TSyDStGzUAgITHCGoPCWYKv+W4H
4V2FjimxHmxFHbkJGwq49d6pGnUISmQgYo3Ik6lTZxF4QQ9Z/61DDaBP7pU9cOyx
WtGBFsSC3Ot+m9YItl5FokrX5ERT8d6m8A/4YjX3R7N5stJn6eaFkPNxhzk1tnu4
TbdSUgXAELrv/FXhFd2sAJk64bZZiAZfQq583SvZc1/3pVs1VXyEtEgwd0nRry8f
97ZUlUIABUa3P0tpGgI03HU7ptzksRcd8Lw6od9a00DMbskDzt1ULFJIcF5blpBp
DUZIt/w/w0bhu3YDZtLDZVxB+dFKCYuC3Pr0ywu5gvtEhDhAIGaqJEPf7ZGw9vGG
8trSdHRCgFkY7C19EoKMuLqDJUepmOAmz6Qd4GAg6E10N89pgaS8udoTG4J0/J/H
TLN0yBteSNVGrJFo1cJ4UiNkdgMfE7HXyQCnd7e0/JBBMa+IC8naQ0gDhF5uFP7u
1PjycRzKUfAJE1vBOSBpSkmXB4eXUIs9jHk9Lh/6/xwRyBKNzcOIKR1aWObi/PNC
dRapy7k0tAY8mvC+NnywT6NbUC+YGVJzuQGwV7AY4Op+Bnm9EFUft70WEno7pENX
Q6uNOywqcdhxHhG+0QQUfjiGBVsvLtzG6WPebU0Dydyd0Y4SmG0sbrKpSNEJqD5x
MD1aTAHIcvS4v0FrZuiIuU2pbc8DsrxFBvgroNfoazz2+0fvD8M5Ap1PamP5yw44
koLLIj8mr7UrnRRxQgG3X1fnUlTimKpivKmuKAprMRgIIwDIYeNtDuu8fgtETPBd
YrcqrMVEyKEi2wICa1zDXgtI+qhFsovGeXlh6YtZTT+rGqE3r5S4GbVb0m2lEx36
bWpKQt1s7w5JEtWXGa23xUXPwSksOUsggch5hqoVEhmrahk6med2OgPVU7jfB3Fq
cFdZW3MDs9pYTnYjWBqI1c2eg48M3m7E0CS9f22imZY1ZrBjLV1nsP1Bzj6FLXFO
Ue9Yk4raqdovg0KJQG5xIcba+XPOD8AdUBRbFntYfkSkhnuRfTzwcvXJ+Tz2Mqlu
fNfps+ETbCGcHXFg3E1ca7FFxzb5xEjqHqh13azFH/OAxFgyPBOOdhFPyiAyIZ+B
qWz+c74L53ssV+SXYqvqFD8BRoLpr5l0KfS9KMNnoe0LRxDKC8eIFhA39dgPi9KL
mEdXzoyjMVIDjF9r/XkjDxxzQ8SStyVkoNxKNsHyizW3MImqgJmo8HiKQoIgXlHX
LnaUmwxyCDhKq9IpJIX3dLsvECv/CpvqiKumvDXqbQzFtzHYsjhUr2YAWhohvs9S
GGouqoswlmLuyeOCuA5ecEcPZ2GqivMW6lB+vnxRFwo+nyvRSo6QHeX56OZRMuWL
4AnUviPVCoST6LYwrwsgHDUKipEB35y7wQ/9FuvgSz/Xn7SRVUI7/yMFoZzbjJjV
pnhJmGTxjPWbDwXCMaVIaePNA8+4oAtA5VjkoRlDnXeomOvi3+0YMtjAqSjaHxNP
3NNqRgVludIV7XhmmARRxe6JR99dD+1cI4tIJq1yRARjgRMDffhxXC3V+FEsalFt
0SzrHa8vglEEP1E13MiAtQzD+pk3f6dhiNKMmMfxZDyXYV5o33wbEndUYlBE9umg
wqwH2rUo5TYV7oKjQCJStjV3chFpEP6FPVx0T3G4SIegDfJYg6kvbm+zUL7V74Ai
RPdFbTVbsAjuOgrirORXmkZDqR3SJ7+9JUTDUY60sO6rr5OrtvWJ2iosTC7t7l92
jDm5kJ1vsz9eHkNxH5aSzXoydGZC8NpLCOhaaJAkyMMri68g72lrUMxwUdM+4yEN
jMCKz08/hSnlyfvG7tj9YB5PeYdj2UIdzLOE9sanEWe5KBF/Z+k9YX7skYwrtkNb
Zds9Glun+f2SobQ4urb9Yy+rpoIKwBKkkUxOCIKeuCkWZRFcOtRcKuLVC8bIHtSt
rVCnPIC8vMwZPnaA3kSWnASQniWT0UndWoq9R1J1yFbA+PzF6Ee/i+Gr1Q67CB36
W/W3r8fJoRJUALdeRoL5OIQPEGaW1tQDJsG6kWFUbr9D9BYl1dSB4dCa/frJY6CN
spND4nxlwn+sGYdgaqjHKF6DSx0QmWkylQB7f31REsLC+ry1EDY8AEbojYOiFipN
h9ke09h3BR5xemjcfKcxMTCikqRsOWC2TMZb8CEffCFPHbXMgqzOVHWIOAcn6cN7
DxcwcCTBWdMZp8AemBhkjgnHIn3m9qQVAIzlmRHD8MLTHxRj7bwn58VHQ0gIXZ19
TnWZB8tnA/J3c6kiwm0mLdXTmXvENHN09HO9HddVmslnBVojBop2iXFGXWZeyaWE
lVyAC5jfBm5ncC+q/80JVfjvpOZTSZoY0dE8RF5q6UQHaUibOP9/BKsmKKFv/814
e70lfmUbgOYw2VZGT4rxXFHcSbcMaMoLjRS7QNzsrV3A1AAiPa9fH5U2KKXm00c4
wMuEm5Vc2kBcLaFvJl0zV8ygrOHuFTM0OL4aExLJRnyymvTtyhVMo3BdiXWBpZy8
UOcAdwBBEgD+8blyTP6kH9D+iZ+OyLdFoRyD5dte+X0rrnKzFcRMLW5urd0YOKUh
tRQrMluluG/+n2anGyfpuFdEcWzOl4fBdel6WdAkROWfFvp34f3WL4YHFYBtnDzA
uPxZw9aY3HPrCaCbwLlO3WLbnbjC+FEMmgpxhBjB+MDxa8hZakSVhiMMqrRZR+zh
BvLmtA9TXfav0WS+byeu5pAfAdB/t6mDuSXtNKz/DlY7dtCTXMGXHE6wt+6gzIGl
mG36AcXDELuQv+pc0r9yLiGkOWChVRuInrlemOIGwXtFSHEZHxtNooIACYYlpXcn
7rpaKZ90i/E1iMJp8UadqoJmNC8sVLhJU+1EmABHM7zJExk6DYGsDfP5HCbT7sHR
LAnmpUeGiT0lGiPKFfD7UUJvL/cyPs+iQOatjISitxnnPZ8nhq3U/Aa+6C3hZiOc
URQWhgGEVqDkk+hFrHilk6f2lsNQ7y3PN2maCej5PooWqkMZdxTMOlguS0XGieZX
j6aO+OBz/9wHFhFoCuZedV/wF77N6SKkDFUsopYt+y03if1wc125/GkDOW4O81S1
i6Lf3L6q3riCTrKardE/cD7IP346v75JYn4jQ+UXExWTFF91dtfrjGI6K9eZ2Iqv
iWtQ/6RwiiWxbZUqSgSwt/V/PmBT9mXqWqyb6Ch3o9bb9Ljyq1WgqjuzCwqOw6OS
aP8T2yA5FxyrsHvxODna2L7H27Y+IMz/7EreByV/JfSvPDWots+SNVCK358T76qI
+6Kbwu3CyyHCYOam/U8ZaDx0DZieuge5UXPlpouQzU7mt7MSUZvfLPjxMwn7ZNHK
ZXnge3B8IaPlVfZmrz/OyeIazNZ0gNJVuGJV7SPSPOHSu15AdQi1kecCWcF4zBr0
BA4Q0WHOm2T3g1Vbr+iNbqbpsfVNeCeJnDRch1c9xFZqh2UrknCGhybqec5TbXCO
AT2iXBqmfL25SBSlgUkEUqhBJb7NTCvWNbdBjBY4MuzUL0VYKGaNAvd47U9JXIR6
sCHp8HHemV4pr8lC9yG8t4zkp7vcY0InCogGvksg0SLVUAq0UKqC8ColTE57tkOa
/IrWRbvheDC06Z1eJZnkKM6lh7UxsGCZBvIwoLFp41/KC7XMlst8zmrH7pPLsu0w
OTOrW/sUQO7x9nBAvQXtu8AXsKyrC28n0UtUDLnPxZPQd+tSsoaYN+bXWFrSmg0H
5RBFV1ZHQHJFJpfZ5ScClUIZyjkQntEBVmRylBHlTp2yz93FvZBiB8A0qqvUCUfA
ob51Fs9xmxrny8hf+MjvrkBOhzqUsmUqqpNksuus7KsCVKinqBqjKd6GNVlZaJ4D
9CgN88jTI2v14TA8fgPqkpo1/NNe87Ovny3ZdUKsozaRVuk+XpQKwGf2Qf4wEKGw
wM7csV8Sst0UaAKOjU60mCNvzDqYkCWllVxcQGCo+VgXhEIvGD9x28AeGwatVSO1
Cx2s+KQFPbxYR/Hk0CrjjXhBsEHAuDn+b7PrJhBKa2VMCmEwUzXV8t3X/wcq5X0i
WmyGBX4FcEffPvxQJg7jdUG1GKfSgIyQiPXnXElPe+rQr8M11lYODWB5AGnQspce
dXAaa/P/00QBzEfT5v3RHbfQzsl7//6AbPpYv2Jg1MF7WpxpmKGG0+qHP9kypeAV
zElDCN1yU66I3iYo6z+BLwFLU6LdDAFNz94JBKChowC569ryh6ZfWAxL8digVBqJ
dQ6jAaCE0Joyws3Rae7Va/RIlILVhMr3UcYi4/IyjelPFEF27pvOo2xtpo5M84Fq
CbFQApj8EC/P/NxFhyrvOPIjVu1q14QVJhY8y5iRp32bS8vWlm35A+5uXuaSHJTO
MfcpZJy0/wzXPiKsUqJMvLOvt/v49zd2X9rhccn9FTIx1xWkqQlWr5ZdoVVT6pBX
wnIXf2FMUVT6hngujFJucpcp6AsCXozYN8HOjyD5TB5E6jXIfzU3eXsXC0LM6MH1
wHenBdUod5QxE4G4kIkW6ymCLkEAYsH9p4FD5ACAVbwLuHkxCnWgWyZaH9TaeUOj
OcQhmvqDnkq92SYZATls+da4KotNz+y/5KiL5iPI9O9HZuQazh+Ul4Q6/uMR0G9M
2QGen3taRLERo+J5bPci+Lm+2Tjb7+Xh6b+Hd5smdjvxeojfRGCP9jJ/bAkBZU3t
6tz8b7+J8pvG8d/NoZBP0UqyugjkRi+HE5GLqjBSoXREwKUfBGEjE69fgDw+Wb2u
svNLFRqEzfKlAadadBCvpIS2J+20QCaWqrPWmhxNWDQ=
`protect END_PROTECTED
