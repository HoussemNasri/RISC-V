`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLG6G2tI58LkgGaYoFSWbdAHIvLKuzwgzt1+AH29odQ694vAcFweZ86bj6icKK7e
S2OkZqBsyYG+J1R8C5Z35O8jzEZ8aV8QCstinXKVQqsAp74bv0L/auP06FTHRMlo
2k19jP+em17RQ4FqnzFgEjLhQXtYRO1zfIJDpsficQU0yQ0wVrGwwlCzahY/JsQL
szkGgjJoc3H9YhUyz8OHV16unasUAK+8B6nmst0k2iNcXTzTXsEsqRmuQsivbmLf
35JFf8lnJvyS1aW81ZbL/MpArwwZXsnsyF6PThuLx4QlLyBlggaHVrvEiTB4Zv2m
Ah7gJIGGLM0A0Qs0c85ucEmu+Ttx8jYughKbryMnXRQ8Kad2R8GgAThEc6bMX8cH
c39wQTcwWvm8sJLBnjod65Zcpnu2xTMt78dzEEiHNLWk/okF1FfU2f5Y/e4aT7LJ
HGUZCiPf4zQDTpOUhpMQtFEtUU4Lxks45YeqME8KUt8NRAUPZhrA7xCA1npFqWFg
VUPqNyeBlA1Y7+TvLRMH6oxPfMeUYjtvFXM6Q2/DSnSoA+44BDq4FMO+yqsvqkwm
4Pu5oDovF25zpGOSNc8ZInfncMaDv+6EjTHuyGhVvU34+AZ7QV6xTICzAyqEjtDV
Cz2OkT6iFB1yz0l2820KJIAe3Y44X0/VpDGR/mGNKw5nfr9IGvEFmVuvPtHAQALs
qFCsNr4QCfyGgp83mI4EwX43Bgl5FvGhMGQj7LK4mw+w2P8EYJuQFBaLi4SsgN6e
ZesMkKa8BXjGzVs/XnMcq13Qp6Y+QvfHXqCu7ZxhNhAnMfCJSspHwkMKhLZvA83i
RscBOv1zTIYtahVf7pRNm/WLgrPhSMZuliK1Q4NsnimaJmeocQLV5SW+EUuePMKF
QyWDhxV8IEvVrH1mHkONaGN9A9wI7ksRa+W4ifwRFIDCna4cW52TFAkD+GxJXSCX
KbcHNfCL2lkpDgF2DYRxHKkofPOcKgTOyqe3RZpVc8WuIFCqrlhX8DFRm4A3JddB
aH0I30mZIn4ZBbJdH/mjt78IgLgGijj7RD4xNdvGCMbRBN9SvsNVOU4goNrx+11G
hyfet3UcdixhUYsQWAulAqLuiFDy8qW+JaKksAxdY+txMGMk9Nr2JgYYewr//XFJ
AMLiZw5hlNMr6qX3LlOfLbUDJG7QWhGUE0BU5GzGDqUroTSwufWCE/onYeq6Jasq
LM9dYyBGT7R0Y6fGcCaWc6aMG8baXwjU9/fgrIWv+cQ+rFtQP8a0UDHYGN5w9eei
Ixu4aoEVDNMG3OI8RJyIwUK3NVCoiPKRcrtMbg1YzkRKt1PnisBooiPCouD0JN2R
zYgVOHipIgXsP3X0Q+0Ec6B3o0I2R1dWBQ28RsP42arm06yUQ32lqJco+Y7791lZ
hyCgeapkzvHsa2rE30A42vOfPbgwL9qnRS5qRib5avyOhGO+mbBTpXSPNQgHcOmO
pibaO3aVECDA/NWFG6YP9OtDiUYDXIqHlBVQ/z+JfIWIVtqRJz7OALOebS7CxLqx
PULE6yRwlHDtP65f4ETJILKzLdVNIoNVMuEfAMNJWpF1mWTDLqxZB2t4PAnKPn5j
QK+bv3wEYiuDZRnLKvNlcVdScgebH2O5O8efCbsMwF/6rEepmNz46O0iRtFWky6N
TQHRNyj3CnNdABj9TvGtaur+xtFfEUUtFv52AeopjX1/gapvtuz2GHg7fl/eNIur
0ErUxn1gMAchKqndE0efGO7ad5tR81bgXTkYeOoGXwhvNNVU2eof3ptYjHtjMeHY
Wy9ofh3FGMj+gA8/HpekqwKIZLAexdu4Xn1yPRVjXDpWK9cA6CwQ9XnfEg4Y4c1j
0FURD+M5xhQYhlRLu+wEWcYiTM6g9uRkhlBjC3E4ImL9K6VxgJ4GNQdlSZu9QSeR
IdMHQk6UL+3IvyrLHtkVvKgPEup/282oWfCZsttGVwrnKZoa+tNymzY1HzDXfShz
bxHzU8rkGqxXRWyjF0xBIwk+GoSnPs/Cudd1UQ+C1jxb03pdknsA/ZRvamNMiaKc
bTlglPOL65TY46ipuqMmtN00o3BLxUYv6lHQ0tP4hFOs3TXnBbO3kin/ZJCR8ZkG
nbSiUOP3JZ1D2m85PxWBLkiqfLY7sxUHSQj/JHuzGrX/+J/BOi6l5qtRZFlRax9w
FGM5wf3tjkv7sfUn/iu0hvs7DMmB8CIPFU2fxUlDWRAUZPCFMnVpxdvyaTin0i8o
2sWcjgxcIXrf3yxQoU0/NJBi+C/X+D8HKjOvKowv2RZnFt6khoa9Ie059/73GS56
xyR2/Yv8QyRXkiQClMO3MofV8xCRh9XbsKxn6BOHSYx5bJ/e4GQiCSUJZjvuZXRu
RELnS9ScORgS2xTEGuAMvLokDfVyG15s5sz5mq/D0M0k7R1P+DJB2qMGK7Jle4wU
W315wIIVJCxnmKdPi/ZXiUWKqZXK8W0b5f17U2ONWI6g4kqKiGvEQ6t62kZUNPbn
+4wWrhlP5iZjevr16bToOOK5z1GmSfFi5+nWtVkvPEZtJMZSuxNJPDsR7I/U/CPq
ke6UsHOBBx2+Xg2XUUK8pvbAQ6uqbd9nV94c992XLEliywufrtC+65LTM0WQAoXe
Ok8zqbhR0u5qZVPydwUiENb+ZPpv6uL9itwj8kvNYYKfhrLkpVwCfAWIoXYFvMHJ
Eb6c55eCH8rjNipRSi6GRMgj2sYW8tZq8KCJknWTar3xFfXB816vpNsyUXcnulTa
r6C+oHm9A3Y2bFFsi5VQ/7srrs6jr7i+D5qEHT4Y9fuHehbiiCuLielhnRslQqZ2
USU3Qa4f7ezo+ifCrqBZDFC0VkASvbypP07w4eX7pR+eHOEhLeIB4vAk8MWjclsK
84KywI4CCK9EwoR9RSCyPka98U0k5eC1F/os3vUhHMjc9Pn66/M3rspIYgKk0RP1
Sc2kyO5N9XBZ42go6Dhk5TjMlc0IvKmxhHSb0123H/pnx2GXBYDtsqrTLyUMM8va
sjGGKFYmcFk6zg34PhF1JnT/pRiCfx/5yf+uXpIwz69WxD63/UOzgmEgdQw1w6jJ
5e81IH3l8fkLTZoVH9WzKkIF/wz3l3YjnqrEK+6KgPRkArHBroGLZEQ4MTbkOWw4
TmOS1kDHrtDyoXQZ+nnfW1hhNsw7/2lrLkGwkHdIBxtyKFNBQaFf6VlGEsoG2jgO
t55V16pNMhpuWDwp3J116lcziTRn7SwktSEkVKuBFIYJ+5DAYkYyMZueqSiGS8z8
wkn1ecs0bAqruXmjYspQbu28TaJ8c/7tThdCy3FuLRBDYs25UGjFMRBHzQI5GDsF
+phDP/gzD60Na0RIyU94EOKSkF+v70iZuCtRwsucqySseKL2ijpo+qEqrwTIy2a7
ZyyKMteEIrU86ntHKqfB+esQ8JstDpqUDpEZWgvtkOEwpaUpR2/CVPpoBXKE7Ky8
34SJhNaM2IjrZtTY24qETdKaw2SX04g8GZPBJ9CfEToiwfK2kMcUtXQDTLmj2M7t
/vcB1AolO9Sn+ojaSzbageIM2mQ3sdAoBwHjnA1ah2Nc4tQtyaZc9YmB/w6DwZSa
XCp1FA72PDTIi76jY/Ew9uCyGuKohUqsh8FXzZ9Gpcu6e1LVC/X9B8Jslp3lOw/q
VTsAyJ+iCh0pyJ0QJvKcX9tuTCNkFckBvDMTBYwfL942PBh+e0jk5JpZhL8tskG+
CTGObA62oJldg+Z8YQkWphFccTK6khSvyZezzZaNtHWRj/g/XjJmARYGYlLjAIlk
alkImkHwHxyUNr7kgkqsxxfnyEtpAOVon/WKgLnEtVLLdy7L6Gx0UmsErnWg3Ofk
VIM9JkYhEH8VwAyZOE/QO6w8+hYnWF01R24U6iQOXdGmEwriyrCfoqDFzQhfJln7
3Owep5gu7pvImP4w9NPpoGFV4+Aza8dVwRy3YteYIDjSSWL4GI5B7S+prh7wTPNW
WPxmF9EIDyzQE9TQeJ7PBottnJzYO18viKBzKmQs3FaaK6aU1OwkhxGldq2vM6ru
un3HZhqUY89pMZb+3YGPgIuk2gugPniNF7dt6lswEFs7hW9Iwz6nfhufj1WJkqfY
V9FuAJ3Y7B8fzIaIBVZA5bKtXvtiWb/r+vcN+5pmYEqz221bwYINQc4uOiLNHC7R
+mPXXn8T8KOxW5xlap3DKF9hthQmkcLDMk11Tu9Z/I2utkZPx9LvWQteibP2yhV2
VtySKghzUxNn18w5DuhkXTYnaWdh1G8y6NNMtW4drEKAM1gWEyetvrUg7QZqEtN9
NoZb6a31V849w8C5Cl/D3zY2sbv3PXwDNsTXze/ajgxsQcZCjYiLNWn1mszHVyeX
C+KHqtGus9DXwILaKqwM/SXN859t0t3AsuwwBA4LDruBYZyjz2icMOSXqDIOT7I8
gVhm9oxdj15Z7TgzRoew2x9VEEwqqZUrda3U/mn5YAtsC8RfjwdH+Mld2xI0pcAx
QaXECqFeLmwddKk4ju2OAFVzlA91FROifHSfpZ9Qa11JqLJ7qkKglxsG5xdoiwcp
VzzRmLJw3+LnJ6MI67WKXsYxeeNTQbzRm7jOyhChEDrrsYv0nbfjEn/Ph/2GB876
l5s30ZHnJTBxBZSLUEKJTYX++HF/xSmmfYam2zkH5yi92BcJOCOtkFGKPMv8wCWy
6TPkeaFbruQCrq62f13p8EpQRns/qptuHPLM/qXiKj5lgep6PzzwTB0a/Eoe8EKQ
VuKeAnD4y59bDONdLkwzLFFRaA1mAY/IKPsUZzn6Dexe081lCTlGbMm5cXQrOBgK
j5whYTPTuDTNCmyQs24/Kxq1RtUh+e17KgGEdtCxrdD0/v+3ElISBI3I2or5vDso
gA9XdWbqIVq/KuJt9gD4wKWY9PMeSbHPKgfPJ6IrOiY1iJvR4aCHgmYyUZ5egjYu
Qc0dv4DthdL/8Y1wjJL63MWmLuqoSZfQGy6Q5hmcBLqJxjk1fCG9Aa3JyD1Y4pVQ
gHOWD40O+jlecg/a2cs0xl2UoXVfVL+T6c6jJg8iMTS9GQj00N/X+l8ySZgil/L1
RLbs4xE2n1Gbe+k/ptB7tdV5lrCPu3vsnRw4qYXRaJrL/cbWWwVzroyUegTD5/Bu
8nRQSvElPGJ8wKmXFRNZNeI+c5HvXJaTzo92fSQTCd0QIhzdRPOl1ngjfuhIv4Ry
PsLsOXy/vvOwL9CPX/4t26K5xkocZ2JmuMUJs+nCQnYDoJZ9XSR3tOwGuKKxkv0o
9+IPXC5C4bp6y3+iuR/Ag1ZH7F2lfo0f01QvOt+Ugj1a0/J7iYRKJGghX099+e/Q
P9p4qJvvcQnHZJ5Erv4p0B/a9QoJ9yGvAtz+ilmpz3RUEBeWRcxIUAuE+Ar9PtSs
glmyoePGtx6G9ww2LhyzmxnWTFSq7bbIv4nZkvdc5nDfU3drWoJ2N4HdRnmJOTuE
autZziOnLKdGmdw63DMr/dFn9gmyqjk03pkrB+tFjh+F1XZpf9ut2SPoPB8WxFjc
r6dzBhqozW3PXY6TfZqx5rEO6Ugu5ll8OWqxSrJPVOQKg+QK0qgj03zBmDnzz244
e6pZQYMrUrhTB0bx0B6EL8mcxtaGmKFwiHd+lusNYCJbqYMYHr2Nnea4YcCqQcuJ
NtS1aDOs0MdMALH2Wn3FddvhAa+d3OjWvpvacF444W085X0dtfqnBdy5Hr7tNytW
1RueY5xx1+A/8xOtuep0VsZu8xzlL3SlodfKnM5C09P8dBxnn1a0XWTiNQOL6wMq
3FXijyIV7naomSVdZOplpEo2GhT8v0ykPZotb2vB+M7cTTOoe/HeWS4zi72/41ao
6Wv4Z9i+wVLSIzan4PBgNEwZkLt2jhMvHrEvBzS008bGsS9NuTB7MZfStYBwlvij
5Yo9tEGF2j/gj8p2u7ER1qB6P+pKbDItEmBmaFQScTEnMU8UUVwaqGwGOeYj23uo
2037p+CU7IW+sui5HSGqSiONEnk7fY1+lbM4VPQCkP1AjGA4Y9n4SizWnljomWyV
9tRhy7Ud6Ow5CK6nPCX02wnWqj11tmWFZqj9CFSwqlUMulffLAOlqVKRNqmmZspZ
cneB3DRFjPKzJCnZty9LA1Flx4buEn8xVpZ00vYBn0L8ScE8z2raLbc/M/5bJdAY
hqUVarQi67FmsyTldPoMwG9aYoSjmYjJ6b7qxjTZCGSk/iptBUlCCkBXebbfWjwL
JnOZhXYmfVGUdJwEx5quRytiBARf0u5ATxpHAh5b/8jJ3BVE9GMGm9ZTqOQkf8t0
nPxXfKsOSFNFvFSC2K55829Gk1evv3kk2t48aHACdFLK+KwNChJP42WqWeAoJE3t
Ith2QWbeQMLNWKQrv1JgGolQ7j0q3L6zI1GDwcGTOPA4AwdQKuM/7el/yAWqZ+lh
TCDSHF/rBQFz0f/DDxWCBo77EbFudNy7gJ/1ipz3fAkZOzIVceblEOgZraQ/AdSJ
Q+fm73H++zVzuib3kXfpeR7Fw21Jnp5EWWvB140zx4QzCVY04nTQz+4Ia9TuqP6L
PKDL4ppst2t1gj0dqJ42zEmIw16hrv4XMdIj9k2axHAa/ecPXUMp65tu+RkTRlPz
LgK412C7VIYqYNcNkobKxCkzLG4FmIU8ihpQl/ik50fbMdd5VsHSQUWcdnnPPm62
kgbZO+B8Q1t0KSz/ebyZd2Nk2Wv8HqvMQR0wVE5164zOJD57NThN4Z565+rCzMO1
UvJUOuPoIrxLUvCH7++BA0d5eNqsx2S3aPT4bOfTiPY0ccT0EMRm/qPSh/n/0esv
Ys91IhK36ee8gfPjSVRKVup/HedM0UPOIup6qUzikaCXlkSVrwK7iqroVzr8ZIcN
VgsrgmmfKmIApnOu0qVqvM815yTgTBn+RPwkIcWQqSsBdo0ag0NJqDxesc9jx92T
8ZxnrIaj6SyG4HdoFblucV64fohYhNyCDRGO41BH3MfJHFBlTHzT2EIukaLqkUvU
IfHn3LgdBPCUvPziDXNz7COGp2vSkaBDFgkeXgdMXr97gL17pqg5FQ1UjyJywTPp
09tLzFMMfx8tOc5BDG50MIqkUMXjSOp5xrCB/sJX7z1bHNIlEtJ25c3BxLumCcYR
RdJSSWXwdufSwjU0ucY0dXiTAFfoVQYSTFYadAz9dOY+T5rS+dTcgYGykGzi/ezn
NO9Auf0Jzb+8r5FBwAc3vRm6ZO0OEWoEXmz2UPxTgM23uPxZtA/8MoQvkQv37YQI
dQeeASh9ldjMGF9GEbV+NH7jxaJVPrlC8JoYIvkD8OfrG0TYjQLbbIsVBPtzzpBV
qq/rFtWeRv5DwTQKUPnP2d7FsiXrde3pasXkihySfM/c6myAV29oqkAAgociWCYT
4fvs/2HlJAlU31CwHa0nLdnm6Kz+c06Rs6hkQvmLjXkS05Q4Y3OXQ4TnxIQ042Ew
7Y9WisAMVvcGf2sPbNBGlRMX+UUN95JQ65v90KBIKqblJ2feGzpyUIG9/6By6LZp
fZPJw8bt31lKNSVKY6E16ws6eL4iVxYzpSi1EcHHxM27vyZSVBAv37SIKgDftiAY
cSV9wfFA6kq7nvcBzY7Mc+CCFa0YZ+M3ug1E/TFcx/B+K2dbazfHotT+SDRfqMNi
Wk2v6MEaB+ZbMf+csJi6O4vd5GrSu+Uz+C5JM3Q3zkPn1kzRkSRfVgeuBpPrdQ04
8pb4GVnN6Tm5H/Tv1S/h42lwLh75JsLCU3oP0B6VUWeb/pVeMli0FrXfrLJp8hKi
MogRWrawekbL75o5SXx4eTr8u2hYuWppZX53hn+fUYKDZFUvC9MJ+2SC1Vqz8mdV
o6IxJwUsdeP4Xmw7/19kxi8/yZl83Szw7Sg0byeDBDmDtcPTG1GAJDkPlHkt+gH4
spg1Fi/yj7OhIT+qAimNpzBsu7C8bXSPkmPgPCg95LdQPHJJ0Xs2tifr7eVP7qcV
6y8rzISrJJ0Ef+ili+3H8fF28RnIM+GqppdXvGLeth2D3+zIIVbCMgwS+lFTdLCr
ffH9BPMDCfNm42WEjfBT/IaD0fdEQWva/o6s7L5coQkcYLQ6Xgn9OygLMQUFJput
StW+iBgImIZHq0Mem3bsNE1gO0vzF/rth4FQUW4DXTOeBf4qRSpJzkMdO/KHAv7Z
24JskqUL8QSyZd89FDPksT2uIexTK48Mke3cO4mrrEdyqOvVecAsn8YJ9Qqi2hxL
roJ2BAU63hG7HzAwPGR/s6CinkYZqztdF2R42LYXOJ7dm0OFkamnRh5QQ/lHigFz
Hnvxf112Aspe2TaFvQ7+bU4RFJcYY1reqchU6gS4gYBZP8Z/yh9br/RdPXNOoVju
13O1aiy9el3zWkRhBgv9SY5yPfdDpefTJDV2fpDg3PJ5GQE9nb87ElWm+g/KIT0i
kbdODM6yyygs0AxCFkw2Su/mIoWTSjvCedKoYYOHHWVuMujec9VRpirgGTdBSvyx
ve8SJZedcT8i49tmyd8Mz11eNujhxK9y+Z5S6xYHAbpoGX7xLoCcolVurD4dz7pM
qMMRUPDvta/Gwn9nVK4znMrGqkMC2Hp3GdMP1Ou2ObafuXxTGd0mOaQ4xgPO6zNj
L3Qr4xZA7ZyxE5WjJjZYfUBQKRu0NCS5ljChJFy3IA3D1RdefzlTfJpOLvYRnz/O
zv3voXBHybg8GU+fNG5t5ASVewCa/5oqhQXxKgFbLxqAgFB0ZqvTEWeaOH0WHq00
XBZVpeaPYYm0JrKCBHgZdkeUAT5oI6BdOdVLA7UnuRtt54tKyOPmSSJy6WNEx72J
zL+/L/mQtp4HsYhnktBXOgWi2e0b1cZG1mwchYqzc7MQMNweGtaG5CiRWnO/XP/l
lfYQ4iOnu6IwYNWnXmDLiWQbciDbr/48TFl1ACugL+gVWgVjEUop53pspox5oXSN
Dk73C/kxZCsRVA39LF5O+pf6rue4DR6IeCw+nPAULkSwlJaXnPkwEH9JP6xzdXKN
jrqmcI70SWlEDUrxr19doaseO+4CSZQc+qSLx0cSDN9TKHrJhwzXeue/ngC171fa
bBcdsJcRAZq7S4Oq9O+D93NY23DhF7p3lDoe523DmTEHIM4EEC0M4rGN1PbW/LNQ
51qDSdEL5XSkY7FVOQCyLLf3CHM2I8hoVsrwAXScIzkaLzxEhd95s4Vb3zhfoxMn
InGlKMUrc0m2Cw6Y4EbN7oSX8mjfK/yEeOv6zoxzrgnwHJUAx9bJhFaef57ZNZTL
oQmre9e3WlOZVaFv5gABrus3iA6IqE1EC4zgDS0msAxe0Nm/S3n8RDSTss5SPm/p
fw/2qtsPMXH4uXfRssSpyTrSNbnVB1MMa63n1FUF1IGpyB3KJZxxBYGKBywJkiP8
QfCfu18G/pwWfskrIHncW2kcE78IDFeNR8WYPLWx9itCYp2mlNDlnCm5jh2VqyH1
oUwaC50V5HDOX0z24rjO82II8kKeL+bEf20fLKIDFFb2OL1aJTtzOVy5WB2Y0x9i
EG665s8GB1GRpH4xJoruhCB4g6m6+S063fptvf+TJM3NoL0A7ZL3UhuJW5CVTy60
NEsx7+8onzVsfw5dj8lom49dvK1YlXOM3mETxYCOH6ZcUN3iXn0sTFHFkIUukub6
wNz2opeY8epaVaoct7fPJi1CgbMdXYWQ8yAbAukVgfTmquFhRW1UrBcrrW21CCvq
rXbtg4ZI2npCHJ+9TkECBVx/6QrsAqXV/w+JPZ/V6c6ey+a58Nwzcr/F2U9QVkFy
BNnohSp8mXlAgwCwaLl01doCn1tJjoTKwZeyPM+Kqc2+B+oHl8/5V49NLYbr1cj+
LajFh1ACLjAzCDs0hgROCafXAvKa3Pe4HtgsIvRDjusPUmp2qNAxKwRCnq8Js7L7
lwznXk4Vcnfp3oPZxB/MKn3YCuLGXFTvoZxS7cWomvwj1ALORIjadYvz51aBlnkk
GHKNHBauj+6gW8jVwfYqF1IsZtWdIDuHHSwgwmUXwTfJuIc02h90zx2Q03uX/sXs
HjAh0X7XYXwDYIOLp5HYLl0sm6xR4UljgY9T1v0vIpTWRClE0OlRu9ZrvKhDbuMt
QjBXuVXwcZk3BdQzg+gR+dNwO724iqNr++9Tzg1jazBWn6huZmAm7e+BZQ9AgMe0
1JnzoQ6kL/zTPbFi2VcoMIJrxw6k3bFwFx8b5GZYxTSghkvCVHiFl2Nwe11hdvDD
2UAjtaXelLhKnDl9IeMk8+l2Obk6a2Zle/y8LrkeKZUSurYOM5DsBT4EaeEwC94p
I0ph0QaKBcdzl1NRrmdN2fqtwpmFFiubMQV/LRU1K+v3pL8F2eUQRcVny46YTUra
k8rPfwbn+cPegj533dy1lGoySWZoWPnrhxLGwXLkeS/38l+LF5S3JbDKcb1ZUnby
F3X9tdcfHRejjlW3pYVGAP5XvpxKMqml6WVgltejEDe2PDwcIUwgB96dApl72Itv
31btyHq8BQ274x8CGz3i5hQ9LNMK+phVDql/daxmReEspR5nhx0si9RiCyzGkcS5
vZCLuac4zjtmAZJMew8CepUgqepvKFhemxmERj6u/IUyO4lxmUr0j+zabEVttnzX
fNVqr6Szx9WWhtX3+Av50ppCibkskKXJORxnl45PEpIqcaOSxzs7fzSf4cM7m/l6
OYS6QHPlADlEEfI7rqFERIcakFc9KF73ala72FQK7b39jLqsX4RftiSnIDJv70dq
bDnE0mFAoecqXqukl/UGhqa2ydAneelCVq2YEzDHhwRWzlgZ1SmYgXyZN092RHlr
4/QUD1bv4evClQbdWTbTPu/C6uv5iGF/319sVRhteuz6gCgvdDxzwpayZOIKHb6Q
dpbO8Drh7icJ5ypfI1KBqiXf2e1ZPtzzT6gMFknDkoDhYn6MnTDVodV5gbFHSkIG
00IpIB6buwo1L8lWhjit+S87maXwjhQUCDCOUw1lJLD9pT0gOroy4FIMgQc2P6hS
0UHH/ioF8SIkfK/UeZNIJUdYEgEBS/G0HX73sKCdWAfNwLCVbvGghoXutcv9z/pU
Y8KVeKKKn2ouJF8bUxHWvEVcULtCaSHkqxdPWumKDw1vliM03+dzvgqn88htY3UU
yWzjkLfiyzh5DBe44ANsqspAU+8N17Bvq/VttTP012QVX7Ra1ytoJIuyafaJh5nj
vZB0p3TMyuOCliDlylXPFUpKhmlNjWlYuOn3H138b8a3vkzFkxtTm1CPryU67m6i
Y7WKKr7lO9pI9sEI2oWYWxyuzQEkClfkLaxTy2w6Y+qLv4WElwXvpTdt/gRjMeCE
9oaaHQ5ASnSNR+pmCaWszcznzhuyLmkbdncr4fC1TXGEIhIkfu3tv8SmSshlYUaO
ImtLSebR/eygijw5y6ZzZNH5zkH/St7PLhKdL7n2apSdFj54I7nYx3KeJkYMm9k7
SuEZsNMcQ0nlTTIkxHdwbmkW0NveOJ8nPH9YmS5JMaqkGr+8W44DrdeK3rJ2mCk3
5qAYGfszehWlIKbF/RiyhwMZTnfOzJQo0Ed/uJG5bZ1zHdPqwgpTrBnC6MBkkQ6L
m2hq5/V1L++DVxrkLnijYQTZbNxdetLj+3zlMs6NaHpNLA/Ve6pscoBSmfnDHCRD
Rlr6oDVvJf6LzpDhDzQqarHkYiiTZFkGLljcA9ZuJ5WaV9O2fUi2mQGeWQFRr+Si
OXTwoM1I/uMWonHYLxlqD7GFjUGcPBn9fVTpdTqSLl+7GdHXG+/35S2x0W8nSm/j
OmB6yfA4/4NCh9kOlHa30NNhIcu2q2nKVxyTdhgUP+GtHnJTJIEkw70Da+k2we2l
gepAApmlXDtKB9pIv6r8+hO3ZgXE4tLpyWQvncJCWbdIeiM0+XEHqo3qZUAaC67X
yCf/3ov5W4hgQHWHI3H0PHbCN+6Qi6dX5+DZa42RFSgde7aEHzyAL7CjDc5h/TZv
jHpQTHW4LirZLYm9qgqvgp59HXaLtmijpfhYNC4s73e6QlwQV/0xscvUsZZehWUK
GCcPchrYhXIPRdG4s3X6LUv7qG5JuejqlaXtNc6LYUAeuzD68nK64lkWAxtnEmAy
fUc3K5Itr3jQ4iDzIjHjGCd50bNVF0bT0WJaiUGsGtGF36TkH7TN3UF9r+q4/wXF
R93zotAhorhbQQzdwJxQW/nGvu045E5lxpnmhZNn+Pa0HjDfPY8nO3nW4rg3/dCV
8lh7H8CVARLYv+bnFHKR4oq3sPyJFMp9BIWRv0vURxeoZGEGRRAw/pAvOq14krgD
ijpt4yCO9G2eOvm21oug1cYnC2M2Z5nNSagWyVvPlBQsY3rSykWfVlJE4pXF+yKu
8Z+8pnsXFslZCNbpsLr1iEJkvfksaQBp5tG2+u/qucOYPHPoHL2di6PC7o0T84wF
19SxRgmAsTyHRzBZjOEQ/CS834bxjbI7EadMK9SaVWDjB6nxUkNeJR+fzYITjQM5
gbwmBxWvtWGuUV+sW2Dt6xylrBCsKQBHmQ5WYeBtt1CRBwsGH6QxhDH6aSbZRXOB
zgMQAyxNtzNSqpDO4WsVoDNJRSCvGgEpfPRXBvclJ+m5uIRK/qJkdWDh4aTiXaed
eJ+T4ZrltWNCDbf5k2I4p6kGfidlrZeI3MFC+lriM2KmeENAzkB96Jv4nTiWmy5L
3YZ0ezgnMCy3stvWC8ZPifdRypdiH1++qaK2m/n3Wl4QOAswPf3VtJR2yT4CDow7
BRSgtx16oOuWh/n8lwdVTw9MpPzu6l77/5h8qBVVmF5HhNAUr1r6APRIGvtAYJmT
E69+URzxdJWNPD+hyUR72/25dk7UX3AaRB6DxnLqma2IaDGLPWoROPzivP93FhDf
ACUZOZYu127eKSPvRPZiH1y8YqlEcUHzC1tpRbslND1JGeRZy/17CcPcV7bhb1ug
kSMjJcn6OBW9N2+GPCzm+5INz7PJ/DgDCqrOXdfo90K9uOQq4mGzVK0pCbf7J/d4
FjFZZ75Lc7aAGzuYtuTP+uAOdCAQhhgYzzzmDrHEbWGJeVeLwDrBMv0EAUVea2cL
1UsAnPjHvDbTtbIgnJSMo/ZsxfKkbs6FeXfhU4n+USGNHBqMuLtes6RN2kNRxo6+
j1aYlvAeJn5pUEqdfBf8bHu81CecfbybvL7TGwkVsjW37g2Iqc5rU3OrvpquZhsx
86tHRELsEGTBm5ESgzNE604wprURGm4HbiNV6Bo3OrwuNUybtatj/+lZV8v9lPSo
ktWoDHq9R4sTU1JKqyTl8A7crrFxaj2yMDi2cTALc7wWjmBMHpeo4QLUGPHb3mUO
`protect END_PROTECTED
