`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A4sdDYaM7jjrPXIuCjh0lwdmIpXwV51Y91GE6C7nuivR4xGwUeraqRmZIubnd4L/
OG2M+f2rvQMSNyDSqdLJxuogJHShLfDKstVNVQj0OeF+cWHlehPh+iJY7LajW8pa
6W5ZJPjmTQcTTIOyrPTAWB3sNcDQYy/O4fSNJVh/4TDoGGh7+kVWLbFC+Ha5vv/U
31hXypKL8Hdy1xb2K9QWfqcwr8CRrIMyZCGx0WSLYksZVqVWDj+XgQ3lbFbozjrP
6AjnyaIrR5tETkRIfynOZkXPEtVEaMqq6q5Xa8AO6iEWnTg2y9bovivc9Wy+UYs2
Ht2QgDEeSLMPYxsjECTcGkVPmIY+pZPVVx0hUvVzG2cR2ZsVzGiL6UJj92Oyhx1m
HTACGOFfSp9qsLfTYeu8PHQqv2MOY7z6bMbA1UNZ3LdnE7Q4S4nmF7GRMpKgQJP+
Yt7oMpBigpyE2+9h49ere0ODnD6x1kjymm7oc3lxEngUcSfoSrM6B+QpcOkG1qvG
Q06xjB/VkWbupTVTw5sm4U84k/E82bfEKaPxYL3JJejFrcNnsS1Qe3SPsK4x2Rfg
lM+6DDBREEiUjtyQKcADHQCP9mpbOaMbXvlxei2FA7cDr4b5Q3+gWRtyPTmo6oKM
6Xj1PeQWmsq/5ETx+DrG/9gauPSBsvYsrjjm4jO/cFVhVWn1DIGpXN+8hTy9CrAP
3mukz5em+75/ZIb42BgtOvKBeIIlWLNxoYpXXjXPwJ6XZKiOzZNsEbp/SIYkphVg
/XWyIE4lVMg4rdlaJBzvPK/vbu9Cp30mEVireHf+IOv2d5RnDPBf0zDiLsNWDnJw
YZ/0x6u00Evm/PE5e4QkstZJc1UVJQZKzF4Tg+zpowwMgGAYlvVWmuu435AqwWci
`protect END_PROTECTED
