`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDAwVxC8grOXmaouoRQLhc4I/k0xJAbQ+jLY0eUQbPs4Vh7ITsbF4A/rLN4c2pBG
NiOitIsZx07s0+NWJmmwQbA7RN5Dte5JhmQkMQieZKyUE6SnMJDuAyMEaOJSmLvk
fqGglAlIKeYdiZMIq0UvTk+H/zyUbubbS5CJXw9jsged1dhBPA5CeZZJJActnwh0
BqHu4Xh9yN78Zh6KKBLN41BUGj+6aZqg9AHL4idKB8E9ONAS1SZ3lMLlYa+ab/iN
gY9uXPVej1ofeMa1E5Xw/u56KfZDtDCzm5Flod/T1lb5/l4q8HqowkP3i26ZLV+t
8CGOkMDwm8lT2zB8m67z4sT/Suv3FAF5ny7SE2nk1RY2DXovdlXua7uxPOhR9Udy
AusZYFjMsSTghZYU3amCHkcFa4+C+FNK98Dn3mxe90Uu0vuCy8HhNJQcdlCUW7oI
fjYmqLIlxREy5A5vvnopKXzfxyyJ99tyabFChB295d5LCHwbSZiVCBRkgQ/DkKem
IFjy9rrb2OsME3CAYeaxreM8RAH2dDe/Sw1mfESx7kp4pFLGtnb3gcDmFdIN/xkl
Ug/CFIEWKY3F8SIbgbVLcftkuQMRcnqr6jzdQUnpcwE=
`protect END_PROTECTED
