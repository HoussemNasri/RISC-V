`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dVbUJzS0/as//DB8F0FuEbcAczYwxTqsooyF9Ka3xWOf/CIEx01Wapdz5TUucvwK
yrWI6dd9YmyvIIr21C66I+o9vNB+W6Y1d7ORBnme0eBVL6HA4GFjG2GJUJJgZ1OJ
zsdh0UrmPddnhMcZ2gg1FVgDQK/k3/8CvfHg+TtJJ60P+W7/7GaAbrbuu9ZLmleS
C/Z0rZoQf1NwTUlM4fdluPPfHqQe8ICplxaFZBXi2J+24fE63x1tpm6zaCPynWOW
o6qRBQ0kEfLaJ4JqyskgKQvn80tYDKnL6/d7C8XBe1KW+L6hYONhlhNHhRD4Et/g
uyJiEfL0PdjiINqz3O5A0R3c1a3nh5NW2TehQtI1cUIE+G73RXdinDgh0pVCx766
y13rhWTUicvLHW4QGI+Rgl8p7briQhJHdWk7p1LEzwCb2RH+HG5I/Ml/cdJyuRtX
qfiKVsqsWuXQjNagn03KLRiB7N0F3p5YocIBMK4z44pl54ginAe2AomsI35SWflD
FVnYT8wd85dbX38wajCLFfJVXXTVsrW8FjYr10GKiZDyfbwpJ39M5Fp6atNHtHgm
vQhI/4pTqEKuMjdiGYp3oRg6dB5vVp/cNhWmYy7Pv+6xh4cYrwEi189yxL+4cZvQ
VVTutH69def9BrvNEHyxHBPDKUwQVTSpn7UGyzRhxWH7xuLvHn448vDpuvqpssD+
L+s896aVDQvFHWVlAG4Bz9C6SsQ1Ml4vyI8fOntKuT94xvMF+yDDZl8UDcb8wPRN
VPDeZ48Pnp9d6dJcQkEuCX20fZgv3TB/Q8V8+p4K6/Ks7HBY2c1BS3vUEiba+WV+
XwbQ77eRmw7891Vmwflpam/w2qQYO/5p7xm7L4x8X/GMpxgqNUtDpZ3mHo3FS0uf
ZWqiso9DuxSd6kBm6YhK4siULleDaNMKKzRxlpyZR6urti7zsqCBfvVV2+ajNLBj
ZKBpwj0bhau9HfSEzjhjCJ3qzqzDWoaAD9MZUQfOpKnzGafFyhmLPJnxUhgZwttx
S1yDYQx7RYiU9u3Xz99EEon3bmCvxwUgHmXsJ2Lt+zhfFJ0A0ERc+hSi2/Mgfo1/
UUV/ztbil6ShRtuLQ79Xs6h2DdKXVNnRNHN2d70pCfgVP3g4kPTg8V8QGZn0OAbj
Zq46Vet/LjGlNumvPPWIHLOGbBtA1BuRhVOyZWcmSWrjibTOBOW1fk7qU0LqxYVq
fdAvdGfrVTemMP7oXEqjgfs66j9EgV+vDpfOX8ChkTYElFxMl3Viu79EgbrpFzRq
lT1KGpyJ3dXXyRKDwEv3Q8nF5HB2u4NzZ4YsWuQQFwB7ZBXZPHnPYiaVVegvrqQB
cZgrNepkraWpnRUTMZu7k5UTx8iqOl43zprge4SKVVt1wK1W37rXQpxyQPNmSUAv
axraI3a8yuhPl9uPukI/pC6n4MnIEv1YZH/xDMT1ymukNt3frRYmUrmZuBS08eNe
qcHfs7T7QzXpvf9zbDq+auRyYen9PbjDHoYoiF3JGZSgRSVDk4zoPJt4Lgb88r4g
BW5zSgeI9lD/Oi6ZV+EIbZlPu3nddEz2k4J5xMD4ZdKbcqY6X4vjc4gXJAU4N/Bl
MuMHLyTTaQJ301KXvjFqjbhmJHc3Q6Gjwmt5wes7rSt6CWw5RdWDOY7msRNYQYz8
2OgS56rxo/opHWXnY8AdLwQz71FWYkNDMt7A8MUw0QQjFvwCRmgz5vypzdhrcxAZ
50QaQHOYW54uCskxkQxGwSLTRUpqG4DAFuQRAey/ZdbFaNw9XP1Q84/7CitrkdZv
CGosZBHlQX88cwHJAWwhUPehDBOMKRNJ8GKvY3b+MJy4HC+lFq63kS760qTIwyxB
7Ie51lxyqXNpy3iWoaDUo9pSM8Y0hN8xnbkjiJUceNbAuqs3iGvl6XT2bIylrNLo
3OL7VlXnB1GJJ1XFlv1bowk9L5Cj3322OPst/zt9ksFDVXbq5Z0L0ArPjuS+ojhw
wnmvYlRRHQVHklH+8kJGeRWw2h6fBPoltn0c4q273oJNwPhbuqcdzeJRthpWwsjo
zx1RnFe1Ze0TkxNepNDBd5ZeSaTY5Ttmj+KIX1lya7vLZQ41qnmkp4aW9N0hPvl8
wh+4KjgOlNdCJ3UWbnxciArJ8udy04SpkbcGb0rx4d8rzDa1vyaMmOO7eUBJnkrm
dWO0jWvOs/QrKffn6Z6es9fWzkKjS0x1RxNtkl4R6lTWo42T+Fn06N00iUDma4kh
1kVGs8xTabOj97n+FBSEJkFqo+xNHiprIS7e21trZNCnWHTe7r9gzLUey2mrRHS2
Lww9TypbMqbPPMrgEcUai7LJY+OO2o5Ds/MEvc9LdWGfZJ3WkhqMKTnWjJxfyJBj
wmEzn/HlSzVBbnXdzKic9O1DO8MNmi2YNXdlZSagNUp8iDyKTV9XSK5sopXpxXBW
2HVxBuzfgNYinAu/eVnVDFsIs4M4B65RjMUMMMX92lCcVAUG52ujOy1Uc8a6UvfD
FCLv/4ehjGwxlabJkOodiYpDQpUSVTvVNicd/yMS3WAb6R1CilKsDWOwyHWXOrMq
lCYH6lefOUkB17Z5NFKn6NxxcxaclepDrzrUsSafb/wMVcAbxI0aHyalz9BxXUib
A1nqrKGThfCbFkcC6CfPvCjoVX1I8vaVdJYm4qLoMTRPOuetrYZPaT6JM0MCpDm7
diAaE24tWw27sCx9BsmR0oA/j2oSVvAtMeliuPc5HChzRy8YbQvjjR+5eyRRDNvs
joAZleMgjP2ZUtDy+P+D+G8Nho/6cqp4qT+6rLeMLZk6SXa8Kbn4asanGI8TUvfF
yRQHKC2O9MFdhZtOLnPCQd9+R7MXs0NMbGsNy50g6b4NwpKnWaRTFa26NktRKUP8
MjUMiOhBgY9siUo4kKHH1fVFo/MwAN/qykBLUBTwY3JGoaymIpGAUVnUjdgmz7DV
4rCDVXUuscmluiuYPGSbZ8vTjeGyvMtmKgqJsJNd6dWZ70kj0QQqETDrhjPGw8M9
08hNcOE7Lqjr3G/sc1Q/mk8IHIX21oj2rdilgzTZjEHLfRg8hl0SRhphFrlhpAvw
H4OO5Ox/CuUr2EzG24wzD+fYt/McvqVw/EHi3MUAdll6+bEcJtd+TpsFj+RK/YoO
dAz6YUj62NPdLY4QiQNm12WalcsQPAd277YC9ddVzNEFarmmdYiKN/8jVp0qWvW/
iO+ALIV8GZX8rQ1axtGDdNRpIHpwpaZ0kH7PcuAqmwzbX7nSY06Rb3Jn2XwPCT0Q
05nnrbHphuPZ7GAe9f9pBnfR4yXGYWd0G92aa1nYgxhFzxAvuZxH3SwqKHwgjg7S
TLCXV+H8pp5UMjoMnkhtbAoJ3bvhqHVX6qzwhS+p0kFIjg0yCPVP1RxAxVydrX/X
OtRa0VFrZxDVF5I8MLCZvsN2XgvrZP5p7RHZ+dmOGRiJW+ArZ0CA9AZBVEwTDBFo
Av9+dpAeQAwoDzYhtPPEBA2WSocBKn7qv6rrSi937DdjnEF9kX5HXsgsv93fdqk0
XsW9jnyIck1Fi63jV8OfWkrOGl7HxHkMxmHoKv3SgRx30rmjXX+0wKEn6ttw2R7y
TBzJR3TIxE76w2yVo05PUA7qIaLwYC2/TjtvWL/jQm/xlM7F0rfIhPVLUqh2p31E
Um1BuPu/n6jMwr2rtVz666j8qQYFKUjWGMiGuBQ0JoFbvvdIIutiMZTLTdDhL4NK
9+CCKgOdajKZmZMJdVq7DBl05zs+fYcPVtjqV9VIhZnCzwD9bsrX3C0L1tw1TNAw
DBQwAwBPqw7empEL82IHwZgNTqS4U5KPG6A28fChtlPfZnHuUpp69gtXSv2grPZY
Wk9k8sKEH2XxIUGB14CSW86lFwzm9VJ5kjIp8kAx2VRT6q62kJWQxtOPV1GXO+lq
6WEsm5ng1mN8xbXsclGWAOfYPsGLMn7o0wr6SAATjDgmKCRWxmDFz5truaOE+WH6
ED8/S0Kg991eK0kgQBXFBzd49cYzNtckQwuWEkEncdKSawGedqiMxdO+XPcf23v9
kVUVlcDqlothIatvO1NSJjDygdUSyKFGq5efcDYppuSbzwoWq7xUQHb0kHKkY1Gy
mL13L+tzSCn08ZAfqosQrpuV8/5iA1TOH2/Fpsl8mfWpJANm+kL4JOJY7taZWrLU
YY1BgTdZCer/dgW6A+0+JS7qk2CNQq5VNDXi+iJ3Jt2NIt8HQRrZLnERufu7OI5m
5ZDCpPOfyXlTH423HTtA/JmfUetp5ksv9z+GAPDZc0OwNn1gPtIGZ0/J2nCFqy63
3vw4EvayJC347fhS6E6H72SujTpSSgoB1HWXLoArSGyfXGyBjCn6n0D9KGVYaRRN
dKLr1hpmta5BUzJ8ihm9dA0B2/TnoRH7sBwpPYRWn2eNqCUaUBiXUvh7sEv00Biu
Omv0i7aBBfUyzoNANF9gV8KaA+ozycqyQcxUr3zHDvhHRfRd2UkCX+lvFh1K3Vea
wWxUccTKZFYI/2RPSiTrGlUUrxeQWsbRBXv8892RNoQ1Fz0f7SvC0ac2kffGPPfj
1XUmqSxtj9mi4zQlLh7qOqTAwtrghT7sT49/0vWmyyDZaRYn/aTDkTlU7shLJrc8
B6n8XcQ52zKWXrnZEPr32NnpiDv9VxYOgGT0eCkWnQyBMtf64lK2u5eNmJ26n01b
Wx2Ng1UfO04slFu7LuVBx9nP7rNZfSm7o70nrIbRfaVpC7S0CQsYmGnuEdf9oIMF
hYLph2yndW4WrHJvxnmfkovSUgQKiC2mx9PXBY7oRYk7ieor3C2gl4JHop12Oxml
eSFSgo71j8u3bPlx4e/eOlajsq00H7knpjoPpgwd7S5Ziq6PlabhkK/48oGcQsYl
Njm4vhCGwxGWHS7o4+nSvFgsM48VhcbGdKH/VPXl/Vo+ZhG70hZzKqqFJiGSa8AS
guYeFGZa1NF8VVz01+KJyD0wZKc8ZN/HMDwRTaGgPGUDDvwUkMRqTcWTrDJe1K2F
odNQqLPzcxVVJ8wp0NLgBmYXveUcjhzOOCGPjOg2/tSb0fAQ6OpuyAbEAVCtzG61
fy1yrCo7A8JN0PvEtR2k6TnNckJqu2qtV4V7o7e98Rq91hITrKvsLsZWD7sSLXGb
CVnX/o9bG+FohC4F+5/219aOWE/7uQKZgbBInbICRS3kOQ0cCUX/PpEdLiRv3XpA
qB9/aiKWNyf+6rrdluDXAGSqPVkdf9hkAReCyyys8FNmsO64JU8mZjhMCtQOEIy7
UjYBdIvoQqIdRMPulvSykN/2lSsN+/20P2SbKjqg39y7gZCAYnI0VKU+Z8Fa7yM0
dNaDBsI9CLUQG52xx5C/I80J5mrKPMao4Oy7YaPjEs3/D/lE22M2GSmIVQtAHHjA
pzBO2jGxUX0qgHlAuMkNnvq8B1x4EBXXNY+z49CBP3lBXWYuBGYQzk7/03pzP4a6
zO8wxFn8eCFe+KuHTLB4jhij3ynpQ77sX9A8p+zMJT3XrzkS1qUwel4Cet33cOcW
ruabtYuKABdC3SPaLlvkxsic8ofwZp6INEWZ676+wlsQvUIAKH5g4W0UD7kqn/tn
FsKydZOJAsIG5r/3JjnrWV9B3VsQJFD/xk5+DWfHWeaplT2gMasPr/bYCfmaP4q0
XNzDMRXekQmv7UDewo2kbASbKwe/NH26NS68lR9QXwHT8cI3lkbdivJE1Bz5fveK
LK3gudD2lz97lKkIne0UfsyEezrc3HlFnIfHINvQUxN8J9XMH2kmEigRvei/M5tN
M2cGGz59wiC3zV7niAqz+K3JiyW3ZoyXd7m7XgymwxWgknY6Ts/VPB3GFcXfmJ6f
9EEX8CcAsitPUfDbXI+AqeCbDKevVKGjqjm6gn7G9YHl3YFGP1xyvbi2wvy6fZAb
JKFWGtQS2UNgUiIpqQPHgkVgp9dpiR9wTA2o1st1ndVdL5OKoM8/HhF6b4Bm3SNe
zjZH+/qgT7GYG2KyeJ5AcXfc8346Z7/P7H6O1ciWu2nf5fHLdhHl/mUOUxdsWiZO
KJz8RAPmSkQmYcsgKSyFLLM6A403Nw4PoSPT0kgcxfKo0AQZNYK6Url1Z/sMYsb3
MYvIxmLrOuIaD7sAhwRAIMrTsQefPl1JU0+kkmuys3AITxPoVgq/TiX8b1a9qU7L
rvvCkgWarA8x6kv/Z46oFrD3a5aX5KmQTUTnYgnPIEXym7kX1zBnTYbIAlcOEHcd
RBWDv9pv9y9dNm59rf8KU64YjOqn7CgtGXK8YHlIeNLsBP808TdVVJP5ttikpdSf
WsVIGCp1EiHhHASgAl2ml57y0wZ60dmtbjC65uhmmpwXyzlFYqqwHUWjZuWp6IG3
SoaSgCke6vMosjgc8T0icuOdZ3xkF3GhjWDmF3kO1cM4cz+5x+Ub/gK4XfaD5x7g
1iF3/bIdNN2pZQqC8asC73FfYcYLTxCDLI3t//+QGJww+h3FoCFX4iuk7rkTahq3
jDNbi6TKzdT03mJH5SjiUMlbHu60mRFH6pZqujEwgDx5FEu02V1dlPg5EWxNR7eE
sWB2uGvJ7tWBAGHKmyRYAz51d4XbZstKhUUyKVb+aRZNQKiydf1uPFAarAyk3s0l
iQ5yj7OOjPnBBEDxMvxGnJHwtEnYEbPnAY8X7ZbjbZCAA3EFHxHixYw/FPzYf+YS
fZWB+SVKF5o3ul/VMUGDiTTcmEHk8PAgQX8LISwl4nhVSUGcH8UgSSMHOcVSGPT7
3ssHZX1c1yWcgsijVylkof0Ay5//2kqKUk4fEa6ff21IunNZ1QptUw0p3v0Gg8gj
0U5HleNNCIafTBNKoHUVIBkKlqQhDrCx9qXCp61xnrGUKshSzSMTKePpt8QCbsa/
xCfuNQRsu5lTyjRI/jH6Gm3Of6bAoj48HwEz9ziJQcDsksAKSM1DrTY5sig0Pyya
ZWjb0lsUOfHhmyUhphKQEUn50qHYXjVEex5C8w4iKM4hqW8+OrONgaif/qgQhWV7
+Eh05yFJebXJU3Jq2sYFWKelcdNCroMQ9SFyTQ6+/CSoUlX5ICAMHeupTwweB0Xv
9+OPg+2CH9hssb9c6kFBXXr4HdzkxQR9kR0Nn/EsSZ14x3YpXKGjmdNy3oQu02UD
yK4/82xwyoLYKuj3lsFyN23GPmSz80+6+V+reVp5STSjnika/sQv38SOikgV6sCK
b5gE3iqeRfyNng9QkmYBHBDrcVK4iW4hq51c+oa8pKv2iXV7jXnnj75B98kJfDzF
F/mKia5KpPBuEPFFTI+Tsk0yWhG8O9cXfgSD4/zYW700iUfSUrb89DHUDMpRoS3L
KPVUWcBctX5WQ42wvgyofqp5DbyUSqgmmVJmnO4YCWGtjyE3NkWzupsbQLXQtCgK
Le0YiG0oZlbPqdyEgEkAPzfXgZjji1hZeHP4YbOvpF54wuxktytFzfy/Z3YWP234
j1tXVKNfCm+DoYYRvBCj39uiUM92w63NEWoIkFO+RymwCLyt+L2FmOJmfJOKxuuu
y7uTn5HuxJ6wLatJxP8CipJSLkFEInvSxBFX/XDpgLxEa79fZF3OSVOnf4J+7Xhm
4GFVTgZUxs9N9XxxmGHKIFdWhaJi/qj1cIunyCevmX/JCJG+irjF3zuT6JVDZkWk
11OcWEkQN15NlzTK5tG7OSixwjjW1QtOdSpyHRQUu4+3pbzNN7x94hQnSG4EDCsP
8RBLM7n1ZmXGFgGqOgICtcAWfZOfWhrp8PCd+XLmr2BJ2R2Qa5pAEDCvvWIArrUa
6n98+pQUguy72DKkT65e+JR4K9fVg9Ff+SpNCzT8nZrzkjyR/iJH0sp/VrCCKrL7
0PTtvJBngmy5pOzPW70hw6RAMs7a3Q4ZPLqR7odIlfzxeeKFBruz470G6Yoj8wiE
WLvAesnKLWUECJznZHE81+mXk0ryYn3ORn/E4xXMCc5j+kRUwl8H8A0xIWdt9rVs
wRECgEFiT+d/i9s5RCNUs+PDjSwRuhsH5XGoZFyGXb5nyqF0PCHO4cI4hPtYgNTq
5JtH1+BmOnbqu2e7sQ+rxErfVHXmYgzKjiqAWAwj6hZ0OG+kTrJmW9qNfyjUt3I7
91xxG4b5oGGfUhv1nG+rxQ46Gj4zepu3zrbO/hanIaLGIQTBnK4eV6c3SylT0vQw
ozOUDqGWQchoRvJJYROk5NSlE8wTWYBAmZuuZBLhtUuNOgHKD+fuY85WhhwmvkxI
v6Tq+74PG5pAy7Oi/ikVnKjNT2LAzSsBPBXhH7dzrzR8G1b7iBwwYNpzApytSwnA
5nyXPe0FfEqXyfuorbYPxx1j+8wQNYkh6RHE8C56BNbQiQyyMjIuLn5qtRFkgYFx
epyuicQ+DELi9c1E+HwUJ7iJg3zL/CfRxS7Gvbg6+EiU3HPe7R01yZqHfQcQZi0W
foqaHADQfwOySUqKe6p6SZ1JKXkZCWzoI7OLmSdmRwezOpwXpYeXTDLZZyeANw5U
dvsFTD9BWmpyvZlTJB+ecu0kEtuR2yzqvfeUJJAbosFVf8YJBxBUHzg3l6Ut9AYM
mPZnBSAIvFY6zJmgc//X2yc8ASosIWfijMcCJxoLHljBoS7BwyZf9u7zFHy2c83U
CYeySGwqMK8DckdHXzoQzpLsweoHSDi+ZYHl6NQRa56lV6OSp2R/Sop/iGLkDeaw
Y/tUmn8535ze2h6JY8qCXuysqWmL/JadhfHxX78+EzCw2ir1nkTamvh+C76pFjsz
68udGd4TjUrT2TBGucoUzzJpTUDMK5kmZOM3sVtO3tOfC1a7txeJ7g0ybOG4Jnxn
C/HpQlGOPniukLeNqx/LeQ3V18WgpQ/JCBCcl04nNV8Vw6JydaQwcYtwm3cL7fgm
mThdnRK8I4UcFiHMMG6eeS4Pu0aVeRU6nKuCuDW+CSgXA1hWr4lWEkAu0czF1gX9
oeCQp6W88/DUB1R+KE6jyqslleaU5GdgvLyNYppV57Ggpfs91L4rx+flMq0HV5mj
L3FaapwiNJoqjIlJ3KeRES4A3SUxE89uhHHaRj2+m42MwIN3FK4DRHBTBgZcOucd
AfC7LP88jCRkYNbaI0FJTc/T3TaSokQMaeliLK+6znByf0l2NjPlKYNAzK/dDlYv
U1PDrqSsfl304uJkeKXuyP3zeRD6bKRxAh1sxzNiNlLXz9hNZ/V95ogID/axvXIH
ADiskryiKs2iQZuk1XwEtATJ6gVGgIIU+kJCWG3vFYXY1mTjaoUMQOMraOUy2rfD
fVly/bRcCaO7FDeO4Rib+tkXlf2VDH+fuFKahIAY7rN1TlLZKVaybncSr+yKT/6U
rNYVt7G9NUbuHLI8zApNFNQdNnMyxSuA05xgXC1P2jEbc/GwBfkcmWXZUt7eNE7y
1KZ2/V9V+LlrMNY/M9xgh1aB5Ba1v0ryodr38NwMUiBNDW132i7ONjw7JKNEpC3X
5cjVZDqAGkmAhvMAcblmyLLKnFAiquX3DiGUZTjWLLzVNgQJlWV8N2FWKeIqL/9L
XMeAB70kMiJXsQmrik/v8/IQCX6U8Xo52X2ZzwOnUT0qqtEMUVV92cRvZr5heNFh
uJXLdEiahumNLLLczE2nNsRMEr3YmpwNy1g5CJWrdP+K6qUK93/XFYKQ/ZyAXrsg
+LIgWxqHS/M8bDhOfvmmXMApjAXFlWvk7kV+LaB/8BEsFSLF6Sgvv7ABUzJ6Yj09
1mKOkHDR9rp2lcdRq8ok7XBGI0+WuP5x3n2+GM3tNQ14e4aFr6vzJZ7FeT66dbWQ
VWAZAW284wqOG8ytjiLAb+9Bci2GYyq5vp2IQ6mB+RkFZEoMtZoFFoX9zM2wbN9I
kKSqKlZKBrH5erak4M4nrlqDbnKTdiyFg14/xKSzUrrTsxR2gqoQZxqtMETJqc65
vkYJMZoFZuKbTMAI1TZwzKLef7DgykQxxtD/n6o4FYQVVjbL3DlnJgRfOoTJZaWq
L8yROQ5lVBdPUxR4fjTe1utQQ+AewTYQYyk0aviXwdZ5bpV/YfGf7vOTh7wuJC/4
C2M7QA3dRIHzxv2i/Q2ofCZsC1AwSkM+wCAUAfrxGPh3fqWPuQdhGkz26NnH/mvW
nhrNSAjubYLwQPNjjvh+/enmu1BbuFk65JSM3+xVh4/h7sWqaNux9EbsBqLfawsy
Jc7XSBOMzrXm4yoUlFllT1lnijnE/5ovgoGmcWs2jmVfxEVqqrREW8OrJrEcrvcn
tk7wTOmHm9ZPL5/OMym4wR3Tl5CGtFAVLRP1JdSieEeFii6kjQFr0wmsuxFZB7DR
+2Ruwbg0qg9MmZmZFWHwaZdJIoUowa3NtvggWuX4GykMKRaCON7F9eTtO3FPszfo
I7owUA19rA33++9Wo7aFScujzxIVuLD+IoWhhNHHTny3uLE5CIUDZtgFOR9dthBK
EoePyZIcxpKtVkEQHpk5fgxooPnKvr08X07/NmdvazRkV1rL7aJUETGcLmapYHqG
Yxuz1e2tdjEkISjl0IN74vBqsvKCFZX/i1F5MJQYLf8VeNVwsqVRiOTZbt0v94lr
NE2GkuP9chzXR/TFRec+mGnAENGDMoXqWLQ3L9hbjTCfUQiT3uXvI0vGOzZNPRvr
4ZnTylEhQVziU8qexMelsIFrRhSJMHFOUxsAhvayAaMAtxCMk6n4EaA+VwKLsnd+
Em9MeAG0XhejQeaBhhZWowGpIAyvDudPsq3Z+t+QpDGc4wll7GkETBi7flgz3N4Q
xr7a9sdzAd/w9YQtykBsbcqCY9wB9/QH940XZldMX3ZnXoWNecAIMltPjk4BozLi
M9WKqMI7GXIDe4f9EypvKFt4BVbvG0gSeNcL4kQidBDYtaTnafIGamdxfJugjtMN
ao7EDsSnbzeY0IJmgKpnK4p/3T0O6AWeR/VCdt8eBjrWcibxwYPbGsxa0nnpHm78
NiUyKtMzoJlNlNlxQ1bimtaA7Ae28x+1OBF6MGDUCVOPgOOipoKsvinR1PA/xIZe
qvmR+cEaAI1LL1b7baT3t1JZbmolsdDnDmKicE6sbpuQ726Z+XUFkaY31NsD7w9d
wH7/fFK5x/PEpvBwYjuKCLeYdEbkEUjCKQbuIYfRGHpZRWu9X4ThH97J3tTm9m7x
3/AP6o5qdasj9QzbBsiyPy0NS53k9wjeCUioT2cdXYbI+usreIXkDNINfpqfP4br
o9UpeEyYX0Vvwcy1/pGnm90FGgssBD6k64bFYzq+xozQkclGfownAc/ANaofHjDu
2seB58PDX8nrWigemvq2gcE9aHmIXtH08TcQMOtjv2upjXVQcKNJTwURmuIYFsaZ
L3y+nytJTEfnRaFfDxvwRNGozhAmpHQlCObMpCiQCDHyP0tBGxa6mFeIcJ4HbYV1
qiG4E4rer23xwAX4yknUxhVTYPxxImsZ58+sXCem5+oF3oy7nr2kKDrLJ41oPDV+
viDlBua0EAvp1aDn0UoNg4hHMkrwTtZFG4Fc9GWwNqjpBW8ADsGxWjfuhecQ6Tgf
U6wALcu16AQ58waZ5QzjkHgcFOivQ07ps9VY5K01kyh3v+68ZXSXQHWEaeLaKqHm
8LSBbs1AeiD8GKNmw564CQO98JLHxGjyvVsur/vW2UKmwGoXjlVjM1R+p5UXsXMe
E7a4Vs834rszgdnuKYi1IsOtB4QmJNNlvumTJuju1Wxw5z+JleM5gxkxHzDoxVNO
YNgWfktLoMFZhzC1eoG+lQbIaHdT3zqmD89Ml5AzQ2acaOCoBoUlwLAfBRxgD0ab
Emp+yyC8nTx5krLSqGXYOJnHkQrPRfA4sREtzKvkLsnDnuxzXoJuwudaqbnbDXwb
dtq4pxp4LQ2KiYBT/dxKtRt0hZyz7VrEkk3ew2HaXL9D6eUjdAbF/ujVZ/FAcq8S
pweJRcpbqQeSasWvYWyXs7r8AAGkRBHLpopvMHZpmX/J4G6eh0PM+Pd57S4CE7pl
20BfsZoX+fRajwLEdbz5b2e9QGdWCJFodFcRE+tkwiLtrrhnX0hpWOLgFW8af2qI
mQXrm2nv2uT++8i0pvnX398Wh0SKx0ZvDAcYAyJDxI1BeOpCf4z4eXb/YJzRCAeG
zgjPLsN/4BWiARYjSoLBaCOYLH187/moBfnY8TmT8A2zLR/Gtuyh430gNPAfv63L
QP0rUMlQyMDxb7Q6lwVBVmAZ1ye0XjKsvDZO4ck5lNxWfncEf/4LKnWux0PadsD1
57AZgRI/RwOUFEaqvK4w0E6a+Y1M9fzEzp46RzJLog0Jgz+VwIkFTl1EMJm80/Lx
ose8snDG9WMm7Ek3/6fGNSZhBwCuHNHD2WQiUJapKXNArMqtpk992fest3MOsNMr
oEArkasifHN5eGkUSV9lfN4P1DpT06CAK2XJon3tO2Gt5UmUDMUwe+1ShMJsE81L
idKkVDS/KT1SVibMzQMifysgqX37m/ECGZVAiwhXa79ZMquhtslTWm6u4XhkvIuE
6oosJX1iJssGGkscR/Socm9xM2i08+XcZiaykZbI3BnXDI9HEr5ujBjc1h7N1t+v
7HzaVhEAwWjAwISpDbDBXg00mypy9+xJgsFf7lDORw00VHis4mBcPBbwYX9cuvSB
KNaM4qT6iVWlUbECSTTeo0oqwpsMe3gGWujPggdziNWzUuefcRHSpsKG/O6Trqs1
4N+zrkIB8WsWuyIVJKNGA34UVssUrlt6p7NF+VgJmG1ff/G0BVRLgXgIKPcAn1ZP
LruGFx7mAdt6wdJvMMBkcrIqMTeJgL8VHUUPh40ZT9ciFHibJ+3WluiWDl3mSjdY
UpDwuNGdr5aslXvAd7xIUwlmZyFtDLDQUaBLUZLKtCsTmlMFTLt8Y9Qq8q0DhC4H
mP7CmXfKWUr6EiRsCRq5r3hDWt8SfLvPQjqsX5AdHR1DgCr7IpJSHm4FSnhnre1b
lWhQLfCiU56pK5hqnddfOwwJJymmE9xYuHR65cJ6BY8x1y10Kv3jJPYiOgJ6LxSx
9IYEc/fj2/EBE9awtaDy6QqzTHC+M8bYhFtN5MK6DK2p+TQpI6lVhKRHS2P5+J5t
PipqGlmsNh5hllPTQYuzEjFyJD/QsXlBSsdSOqJD9RmFQrW0H+uiDLFa9n61MsS0
SCXkkHpxFoTSEkZjSp/D66UKzDg+iJov1csOJxWNgx606G3qb16lN+A9O4nvZ6FF
EUj/zvlxURLBXSzBp/T9YT16PRO/uyjivSztan7egGYke1JEZE7FihVXFsiycSWH
BQh5xgIYoEDmB6JDMbYmntnmcSrtax/OyF49RygvBPyPxgA+MP9US0RJHGkheO1Z
1TFCuViTjHc2tkl4/8Heyl5hajsVtIBuEcjnHaSa80VB9/tqVH+yWCsP/e7hB2XN
5FTFhk9Tmro36xv4PZ8Np2n3lt4J9WuQgYbE0XhjLQyizlwyatv63EoxNrGd0pFF
bsPosgQN1TVDcYPZivxCMxG5CiXHEgVXyCYvHfVs4nOujdoBr4sW5ivB1bP+eJqi
h9FrL+JCZs8CtGCRApSho65C2XR3Ey8FdqOR8M+3x6EpLwpVJ3PFSvWs4V2dX+7p
17Xhn4hroVqsW55AcPl+TQ1aUnbX5PeavjKd7l7oxZ20y4ODpaeAXv3cZCRM/G1V
QmUERodJbTg5zt2DVdJOLAoxwta/fHlPIwcas16P2yNbtSW+CdtuXtqFJjyienPm
sspFENwy1BfXjuDeyKhcfravkH0TkD+ltAEcigmd7Peb+uh4v6L00Dc7EsMxYp17
Sln28kuJTtrWEAXit5mT1EuztHeaHBd3Fe8DwHKCIZD3MpG2p2FjtIW6CGbWSIaO
4pxGdNO8VRJErI9d3hCqRowfjp0+phXhdyir7iQX9RQMJS/O6EIUemjgU8UAj+x8
1ewLbqsS9YnV1AAbVysyY7p05GKr8yPhnISaYt2TUnQ81kR4ikHhCqOUeomyiAMr
uaEHdbYHIRp57f36b75VGtNz3xMhgI3QehbvwjnJ5lwAeylB7G4XvJz++HOLBbA9
9veMQ2/zlKn310J2rPdPSscFPLiBxgYynN6OCIRgzQxWhqrUuy4bEWazqYjgTE+f
KxR0DgwpZjoZfIGv0a1OhUOE5JbhMygTgmxdyVcYxuOjkrgftijDhZnsC/lBt4JG
QW+7G4C6uisGmxIXFnGt0HI0mSQ1N9iRNxPfnLbFSCXmaNEdthngLqCSUV6siLDB
Wmb64gzblZ2lgcn8Pq/i5iaAVkQ9TXd5+NkZ2gfjU3YqwJHlqe88EafrF55exLcO
KIu7V3fqSwGdoxaEhXPkEGAda3JneHJyEKer0iRZoZXxIdxKJT08VmzzpskcJA+M
JCIJ6fAd1XFoFb+wsggsip2KRFhgfisUGf3qwHplpITmcPL5ORxUqTgAnAdu76Cu
u00Hw42EAq28sgWtdOhnqQ42YEFLONpuaWW3grpM+xEUtkU061fX87rDLatxWWl+
/KGGBqJOAphxap3i07uXXo91v+u7ByFDhTXQ07mRxLIqHWbAFDzi3TKL3TtwC0NJ
WTma8jRvmhAPeieLb4OYsYTIX4/3KA/lmJ+uIIOTiJ0MwlNGaW9Fz8IGWH5inoCA
rV+BH3t8XxdFsqN+IK1tEgxUxUPiPPoncuuFr/Rov2p5kWiGmrM0k7dsMY3vVV4f
sDuXIhnpampytTDS64fjkGt8a45JJlxQQDXcFpaz2zmIEJNmJpg7W98tRL2cKdEr
2LEyXQGiCCgW690d6QMyEqfbvvM17EKNMlPo5Ozxcag2cf/EoLWACtoL9oqmlaV2
A+5cYflJVPWRnfHQr7KUXu/kujQMn8HzaP1dwXmr3WLS1Kw2+WHy+RJmP+20GMi3
VIzH5qoNE0uBLzzV3kFAIDyh50WMNZNhpf52thiv1rptdkDo+GsqwymSs+o4Sjwv
XoiUbQRelW+ovA4eY5h+0vxhZIZvRnMZcGdnF+j9xA9a3A7MJ1/nufQujzdclQqs
wYlXPjab6ry02zhRoUSTS1T8M1HoqgvKs8m9Uo18JZmVs1TMb/ir7dRr/0VS2zan
jyb0PJFCkqqdH7F5sfwJn1bJqjgssLFMRTrPdD8WXe8epif9At6tFtosaP+ez13o
6tiJwzFbIzkB3nE5DOBv5lUbD7ertOWANSNt2O0OnWtRpdlO5wGu5D5/lFCZcHKO
Y7DvXEQH0EKEPSiKGSur9H63hFw3s8meE9ekPVkU+qXT/O84AxvaH4G7ZOJBN8q7
rUe80l0qqY4+bek22su31/G/DUjp7MrMl7Hiu6VtcYL1vPzJY//W4uyiawjv1pKM
Pf/vD7B/Z+GkhUB+wYCC8xIum9pLySs0IidGfoTG4dhOsovWJDC+6iBb9rd3kg8B
ikygSGEiBdbqxUWtZV0zslcVMmHc+mQTYQW+vOds+U38D+ZdSAOK2oReoKm1HFeD
MapvS+Mzm0X/Lq8alRwLevBn+o/wGPCHbKhranlFKYGXW/0w8o2snYLwAREBfHk3
EmxeRjEok7MFA15xfqfDEJSBwQd8MXwTlX47aqG2LwdX2xNG353v9NpQaSdxhXa8
dgr0/mMV6TzhVeOLzo3MdOJVvFePADp2ZdVkej5HHVU1nvteatqTw/bmmlrNJb1v
/x3Y4YTEwLq+QL4RXnM9CkasZJeyh4y0k+1JU4eBu8RZzcQ36swlpu2HqEuMh8Bk
JHEgmmJj0EPYAnYy+OHINKabwuikZq3i/cQAUnHowAWP4AHT/mPcACIyf9QlzzWe
LjTeMl5V7xZtnto5+ypVR7l2lCkfQokgu5XYNH6kRCdLx41EeoWwYbSpAvLLHZsu
Ifly4+Jx/GlYeL9dnea23KqbONz0KDRQzVChoJPKZA/sJdgnP3x45qVrTESmCsnw
DJ9q5/X7ck8RB6Tn3OwJ8AAx2MitrnjC2GwVEzFxv+QlI21MmhMC0QBsjsxV+oDd
w0uVbMvYDVk2CXNLfPl5aaBFkIs4ONatqD66iNt+ljlYCceySUXtnhAXSesL6jwd
BmxssBzX7YM7EDBjj82ICU6en3W0S9mqEhHEkZl+jIvyrU5vbo+74ZFGDbgqwv44
UwcIGVNQwBXKRe1YHoYKUzKvSH3dd6piSrLOpwNbilP9G95QUyaFfS2gzOQHp08p
4j/H/QwdHF3FKCjlXzOwNejJBHMH2v4WwTY5dajE04MMSu0j0+qxTP2BlChFviWI
IiMz5ALhuxLg0ie9Ba7RZysUd6gdRDUpxCvYvXqh2v5/9SqjcJVY28pzIMn1tc3I
UE2LeQi12wapY9wovTAewP8RKx0juu/eJTuAAfILdH5y0YVr4/MNGinPRzaz36lh
7LKJDLKgMVV3h8tubssr5Sl/WTi8vu42H12PH5fSk8z2CDZVBEfqfjHhIZMZfkG6
gdzBoflXrUVxpaVU54r9eEoK3XpM3MOoKoyodtoAWuMdif9Jdd7xinaqCOkUQaYu
S085oaqhjbIh5FZYzyaVGMxSpDEVUJqhgBgX5qyfg6A4V+en/3Keh4ibsa+WDlgX
03BMdSntrSrro+bOtEyJUKoeFiFg7zS7tRabyc/f/p2ZfEfp/kBoccb8tCUyj5rO
p8Zhz4VlcCC2lC8i4JZNK3FgSAJX8I4+5fkOlG1MjUiZ3l3VCwM0F1AoD8g+Dat7
jQPRT+rPnzLWP60mpg/fTiUA93AsHthsrrEbyiRAnYB82ZMLjzgbW2DKgzmOKV36
FY898yHOU19n7EF1xNKg2+EvKvlaP1ERfx3xTBd0hTVtc3zmwQPnvQ0nRfvoEyz7
duiv8gu/OmRg6YpaaVA7lwgHXSlalcbQAEFlwCOJuUKn7uHjmSOBE6k7JZm4LBku
49nBw+z4b0Yctfxa/86V7V2TEuR2WQ/xGfsjxbEOJ0C3KH+WlDJF6BwsGi4s+QRr
5bC1zdNMokGL9veioGHPyACedvXiX7xeqoJrWCeJBOHRr+E2AKftJcsNWe2i9RZ1
X9DbtC0gzlOp3pyK5W9iT+Jqv7CiNU/4aSlTjHoQwBVWJrSvwE8qELHfjN7Iyu6y
h6uJuNcTSIyCJe4nIFQunyrf+0Zn52lW8LS3/jXJr8l/QDMxJBh2GrfHYH/B5MBB
8pTD+h5YZKmd/rP2j5CLMVsKt4ekwV7GMHTZbElQdVtGHgSre9uIBEmeDf4nGVHc
SMT1895a72L/5MPaEfpr5sxkSwDT35mwOI1fwQpkrCuMppu5F9yzyTDVYaOMDCFq
a6lWA1Y8UAzVshxlcjPC/6FvCaGwgCTqae9tDOEOeoF/aRc+b6dyH3upOUHNaKwr
HfmwBvxTGXjEEJKDDhOiUUFlol6hptzxEKfTq8qzCdrZWiVe3fsaL2YBcWomGI7N
l5SlrStqp8YdFu2qI3qHEKIoaZ4vsYLBRBwqG+wsqE3lOW544snLhmvS244SHJ14
Umsy/TJb+OLjP4BPYzIW7vHZ6qT8w+LBKUjKa2rOvlhAV2Jb5dI7z5LE5jnfKws+
QnSwFdm5Lx4g+R/2p3cHaVxkpQnLHszVTwyvhfxO5hpVJfXaGlj35ddUPQCQ55zP
CQ/4HJGiIqu6pC3lHLPf6f4vAOnodync2PQr2BKNEesl2wo+nztBs1dzd9KLejze
9bC+0yp//YdUyAoXu4ebdp47BD9bwasZUt2IcNMDquJMsk+Itu655M0vm3SPh/7z
8GKXwUEmB6Qkbxpx0bJk4GBKuMTO7FP86/LH1eP15GfSq7xozMQC9cDTiCDtckJC
kAlBjEUnTmw3Gtm5xEoNW+eSevY2qTd3cr6ibBqNzMWHoI3N1LiJ+slFeW66d8Jj
rulnxH2RggaAnyBpr9x/zlcSyu5orsJq8oHiVgvM4E+FZAXJ8tWU8yoCH2GXky+B
Q/VxNSNYIUDsKRgKZSlS7NoQog5WmlNKI9FF22w0TGlzT9fNnz085D1jX4tCcak4
ndUQ4osQ8FCV71CbieacfRsJFwUj28/ubljlg95OEzajZO0MoEgMXGouzwrs03SE
8b/VrrRBj/E/wvh2+qTjG3cipfO1cA0zupdHCM9sNs57EMPrfNtzYrDzlAVlHgPN
Xk+K+YXsBjRgDJs/oSfsMI+dR8/SJrlK2hH8PqMYcxam5g669auFIdyZTGS3gKGF
3zMmerGA89UnC37F3b+YqFFctzwNKfqH7w5P3EApnQ5JzYhvfnssIjUeezVSjCv+
bK6A8LqxY30tranTYSHukICWBsX2pQiRy16HtuQgH6VMOgcvurGTvpBR0tNGapXc
7Nac+MNn0hqcTQLXYgDV/m1fhFTBa78Fl0GT4CMMj67+dAnBg4R7ty00ddoDUNe6
BY1UvoLs0hkWppq+zQlmLqbdB0p3SSkNUhaf06zm64UEXFZf7oyKhUUvsVtouasb
KvhWgDLquiP+BlCAkzm6uB1danIlYHhPGmlPQMGQUM+SmlXNjkpl3JHTZmRaqVAz
SgTvj1ZkvHY8Wveom15OueLk997ysIsHE8YUuVHdxDQOtHI337JDvZ2rrYr3PD/A
B+koVnUzOp/tYyRJNHLECnTNfd5CrMoXHENCcKhmatcbTFG03jVFM3hbSEaXElO1
MoQ61pN7d1ryrYXd2O6nHupqlOCnSgFmZvgzTKUXO5u1AKMOgIhWnD3jCepenGpE
FROu/7xueqflTaEhbUui/85IsDmcXLYEMs9diZc5TGTdIiavPPigO1mUGCvJpEIp
jpBGid+tKcNSQRlpbd6ExDUrmNOrjDpTxLf5iHz1LnjI3wnIbMLFbH5457XXYi8G
tXXF13BrRTr7OmOBiLhqUOQ5Gnrfoqi4ur9lvlyWhgwSI7sMIOKO/O/VlYqtGTZg
bQgn0RbF5oEJ5pEYN3ljV80NlAGTAVwhkLuh8aPKPHYyYUXgPxo0yyBirnKnCbFI
dtAuFWD9eu5b0e/LoKvXCSESFdm48vob0rQAG6figRgRwPCovTDF/Lawgf2+MYKK
XrJtOJssTzOHDzopdxVDugdYeLyUZzCztNm1Xh/FUjzuTg5Ezdev2OsVXaXzx4Wa
j6ouHUrNDFauj57OuoaV3Cq6yS5sbxpPamvWnN50RLm3XtEHDLMtUjS6d6PztnhC
ZBRHHb4w+zXMKUI1znJAAsuxDzrIs33tLk4RCq3wF/DBRMVCaTlImfog8PWbcaxK
OhUwgI+b+EkbcHaTSLldX3SZSjlwpgGVDhXXccT5WKQW7SYy1FaCynCd493HLR1I
/ZCm9mTtRogzz36gaZCQNcu4TBeey2smIBxREcXeCQ79ug6EpaGgJFAs9+xwc1Ov
/Tq+d8MhrQXgbBTkECrMIUdhjDoM7LvuNrv0gTVLHfJ5aeHtnNV+cJtvKGMY+lz7
LL/qlVoRvYJSbHSFik5Wu/QafGebnTTA+9z08XA8LIUMqg4Bna6OxBr1ACHBZnJK
badIXI1bOP/BI0bSq04UdC8cCsRqcHRDiUDGLzAzKhLCfFE9ICO1DaPN6VyOWFdF
4o5ITZg2okUmuoVp2Gg76XaOPzyrx9eaTk2+5IxzuQHFT65NTmM5Ofnk6uq4L7Cr
HtK1zWy6U/ksaUl75DnPlWCVk61asZfzjvORz5f+yOdhAzDo4QS6gEd72oJwZzHJ
1dk4fXZ0uYgq8xlEoD1vEupjXcrZTF6SrBRqAndpFkARtcC6STUWKJRophjp3Fr2
qMT1urFXxsEyg1hF4DAFfHe8gbAb6VoSCauQIak0Kf/cwy+LDTr75BaY+wl/o/TN
KGglwgUGAHNHni4ezF0S2gNW6KX0p2KYEDdUgHtZ2F/5yZ9jjRuusn/HdsRQBjKY
YqE2ME28nKjBnVSq266cMnKk++fKDU4uF/s5B2RJtIGkqds0HJRy/+vQiBW9bO5o
wcz+DE4EuUhDIt1SC0K2VqKnWE1tRcw/vuNL83ydn0FkMkArIGyml5FEDveGz8J/
HK7zAwWzPnelJX/pop1EmroDBLn5UuA3/tU950F6/Pn5KsFKdGe50gTRW62CBmzP
j1qAExk+Zez+sOLoPb7Jz5lK1iv83p5O1pf2GIXvjdld9os9MhdSsDddB/vQNLY8
8VcCeSPmvykYgwKyRRuhBDdtz0ykCrnz279IY1oo5BdU5FenwKM2dzxmcFuxQsSL
mC8Kao1hGmJRZdkKpnGElKBK5RjMUSSm/KMtaFv4SndMU61AHbfjVpJIBRKGfyG1
uPMBwCs3gpw6osAkpnmBw4+9Wd+ANMzkHmWgHt/6N71X/+FrJmyQFpNwkl2TyTPa
i2hb0BR29wHj9gsAyQl3O+FRP0JVIBiwCsUFwOBioTtpALsz5+qzeDQb2eKLaGh0
NR7Jc5n6/tMF4V3iQnBOu604obeYD8e4bRu3NeUpAEj8QI61Xx2cbZHJLqkWZWEy
DX1+v/tV1THhWHyKapMN6eMZbKy1fb55ULfcaDYOHLkqcRyFK9VpZhbJ06WDPqBV
igfzBA9856K7+7pKeLvyRgt5ldxQOsraAgBzKAa9uUWYSi1qBJHzoi8m0hv7Wv4b
wtPxNPQPg3E87N4+mnHorgUjwSmXqtbT+ryVLL4vFa/ZArO62vRQMa7ARGAXIotR
PehkXNSN+pykn0WjWjGTxZcNCzz6lWoDA8a8q9NbxQBuV0LU28l/IZzUNoXydKDO
77EQcPyyjoubrleOSZ6FD+d7UeXaoNrA1LdgUbLDRsMr3GxThW22USlQk3ohPgrP
lLK7v2sqVdalH9ofcLXZJ2LOYK7cfFd+Hrszr2i3grt/+ErVaFBVvKAX/atWrZf2
vTXW6bOswUooFY7AxTt6AxzSP3RjBDdeUBSWOkpJRxJO7a2Ydbxr1m0JzMTReVfl
/T8uo1LGMrlHCm84O656r4o3afUM/U3cUXcQY32pBCzjVo/O4KvBemBU3JwT1qF6
HLxHwVU/Y/D1ki3Y7fY+SOF4QLpLMWBGjHBDu0DREOmUqcJThxC9T4BvWE7gIZkh
k/VNVhEDzqFsRYu83Bf1X8Y3xNVVpdBPw9YXOz5+eW25taNIStzq9+tHcw4FSF46
//3hRH5zvMxHl3CEMSXKLRsM/Ecvky54xwJwlGMPnpm358cxlO7ulk72sGvCDdH9
hfkHPSJh4Xn5mVFlu5NbeLD1d+SQNAkUlnx+bKdg338OxW8uqFd3FDMeSWDl1EBj
RGyx2cqB+Vqc5x/U2iVAtf48oPexcX1lnO3Zu3vaT7UUgGf4GSNANLcyQ9dkcC+2
xcr44idqBpCWR6zj5weSAnZmKbXXq5qzy1/laRSiCyTrHXrCneQ14WEEb0qZJ0Wm
jEn5Vn8ZkM3H/u62jtoPzA0iH47x4hG3f5mbpGjXbfUV5Ip2b9PyOUCoFRFGrydG
OSZuBjkOW4ny5vWb3v350epuyhJrN59Frh4tlZhgi4dit75VYQpBCy3RSkl6PvjQ
ROTov40upsV1H5eZ+9UhRnaMJ2snFTKHLw6VSZUcAK5XdneQgQeT1Ir/34ipUzUZ
j7CGJHasn46UNbPPu0HW5EJCKQVEK16NtbSOdILPzE/kwTXaAulnMT7c/Ax7T/eG
5mqLVvlMG1GZ3RxLhqi5tCiU2uSMQqYjtSCSKAlJwzJD+ZarAc5xg7bFrooh8+TS
2GuUMHkzaYn0auZXya47CbU7bnJbtC6jTcOqSaRm3AgzjKfsM6lPqTNaxWucFnLh
ZKVvUAugRjKQXvGhoWcThOjT3yObNo6KuthvamNvaNsAegV/75iNbKC2/zXJEK9U
Ujft8BiyXyFhvyXEGNgD8Id5RGfxT1szbHAxPR3bmvxQ8H6B4rysm5WJW30DsXcY
PN6GHXnlKt1XdivmQ9Rg7MABvfL7cZtQwVAmIyq1JWQdWyC3ouqD6Iq2PzdCdm2f
HAKcBg+eTowvX4Wdi3UZQHLuN+PUfbSHq5H6TbXcvceAagdaHd0RO1O9itbz6JV/
rWYig2uOZYnSqbPzn9k7pLHwPmNws3XuSOvGbQgEgancGZjjChZ9e1j2rQFgAxTH
5uVOcF3CrMyUfzx3I/iMB8vdbO030SBiknpYJ9rHk7hw4iMaMeM7aDWhoXNdtUNu
234/Ov4u9BdQ/3BvK5Dbhb54AoF5U9s2Ze51OAYJQzECeDPELjC+/+1Uv0jup5OH
jUz5r8CRFHMg9diiSMRBb0ihChYvgkkFR48Af2+HZfbx6Coc4UNbEoopS52zyE+M
XJlh+OaSc5B2BFp8q/y2WPVotQd4njB+Vax91VyJQSHr7bKccLonjDVnqkmqdLnZ
hHFCGBR4lZ5BzNvzH8JxaFBI3N0tSOXqtz3hfTeFnBKuRjFhsAfbu+SA8bVgDME5
wPHFTeyAAfDri2dhsn5UhnzVJsqV+AmZDCvncUo0kqehf1ZS2GD5GfSZUVG/kbTP
2p2o0Dk7t5S9rYrzwZxj1I0osanJ012kz4o9J21l6Fcsaz0zS6telq6fSkmuDeRT
S54CSvUcBUNTUzbDpYgb8X8qkdEzjLaBvZ8Udrsu+7plH7B/CwVBA2OjJquIsF0f
AI851rlCq1rzPrMkb9MDs/+rVUSaXg06WDMyPpyundNIM5woXGrWYL0/YMv4DAU+
OJl3YSXDC6N1+Aky4zojnp0fmrLWsQw2qmBRj50dqg3A0cSRh04ELWMqxL2vzST1
hXAi+yxILt4CeXQaZoweel+M6QX3AoW5k8xnL9I0dKx8N52lbgKfpzBptsI1FH+w
IrKr4cs4e9AtaKGWeluF8LK0cwAxyXuc46PSguVcvCpkdLr16pjIyOLASn+Oe38f
RACAYrFF/mH2AbUtSVKBnWlPgoG+D7TCg7M7osvCfRr8vg74yP46E0CJz4EAvJee
4WGeLg4CKgWY8OG+UnIsm6anJ3isvKJPQKztIS9Loxmo/4CVO1jytN2vS/z8H6Lm
Cf3uGCXP8NLIuLTtMVGZGd/po7dq+Jx5mexs7bNbFKJOxdQtpPpj4knEzDuc3CNs
KIl1Um29Sxd8oqnWDhaP8Pa5gc6hICFcLNK8r2KTOI8Ig9521L63V5gp7itc8MTK
13Eg9iZ2o/SVhLkueRD9nlOPqK1b9l1W5c1vGCEzAOLifJJKl5lvWGrnrwBb53WL
USaYbU4c3fGuKUa4/aomia1MOEbysQh+9PWx/yciuspFMezPSJx6wJd+W9PIVZst
o1Qpqj4Mjslb8ELhdplTjXAu09aq1kpzwKbUYpsxxM3Kc0DfBeW2lObRuSSytjRO
7JvKdFizxgpbKfjA6dm2MlV2Lv9lRISrgDpisadSODxEtqMa/uAwmys0aypnJwki
q8u92xBVVb4dbaWGd7gCVKhODxIx5H/PSTlyvkTa1MmBqOf+wyP9fdkYfXh94HKk
3SmNohWoHFJBdmFxxr4kDbWEwiWjhds2XrxBLqi6VaOnRDSGDg+66wjmSuY8ybfZ
TyGbEimoc6tx1bQRzCDgIUUMpGeJI4L5siJDUD85au2earE+qI2cCTT3/asqxcWH
D6t4iGu1Kcz4cX8qUP2bpGlJNagZ2vw5Deh84m5t6hjh7KvyVOXcRttXoEkx1huE
7DiWj2maKzhSNz1yyvES++Csw4dtWhihOnrtBZQiCf8v7wp7mVpWEnejphMCF+I2
LYsxeKqVkF2LGutbJJ3SKsp107y+UiRqP2ajdgDDQIbYzV+eiH3Qzl1yrAUolLO8
iTXuBoqa9ctEvg9CuTdtQKwC3yFJd8qHAQiLw4I860ow0OD0k6uDyzVwpVj0iKdv
KvR1218lhzi9ZQe2U9St8GIezQPzXkNC70qybV7+bzFjPALGpQFpISmQ/Aqf/p0W
bryJWPZhWU9TaD6BEQ3oHhxT/N1dlb36Sty3J3HSnbtjLypsAZ3lLijibqZmFGtx
lPP0IzB8K5kd3Acu7AIr9feFyZPrCWxcHHod1fAxLHwahUu2LXCysMRCepsRqRZu
ZEkLXO5g92IdIWRwvbc9T7giJTc01r4nHbdUpChWvJlxEoQw2TCh+qOSq+ANoa6x
nNCNLMp2vAx8zzq9J0NsoQMmdRcpDMJQeIXwAmvghF3s1odjTym3LNHZ432ogqVJ
xFQ945MHYHqyMm/rSj19V4Ts/X4Q++9cL7ZLvYOWjpQWQe0G08+FNXtz7Zm4LbY4
0dzAXbbnLGebK9VfdkhfMi+B8MeioWBf5Q9SHfNBISnvF7V9+AJDb8GojxHB1Qmq
ZlvnqYUquu6hwzcvaGwM5TA+zIhxO4x/NGxeQE2FYMOiASsPJubglHZMGHCp6EBP
wEoFkrjPt2JFy/285n4pgvLmZsH8VunEYnL5fReOHhnuaI6EiQ5rU6L7pVJU0BZ9
nSykGX50O4HoBtP69ucLgg57rL4UhMU9V2INxKv3kej2y6VOh6LGh+bwu0bUQ47E
lmDpd+y51tCr0Q4DzJiCFU3TXGGW3yU6EH0cgDdloq3KTy4rQBB6LNf4caMPKTx8
uN3sR4I9odb2TRP+XJnM8Tfwnx4WJlQgS4VpPY8IH70MF5kKiRsl6VV1BjBniAU+
T1SnFHQoZ5xaRMNG41ijmA7QM5QFqa3r6Of2oX9yoJ/C3UoeVFFt5/pPZ3FSXixn
cx/Pc6FFsjgllGqp5/Nqo1WS6+hcW7U6+c7LE5VfODmykygyNpFw7s2l/ts6sS2H
ol4CTEK2TKfuZDTeVnQZkEwynkvBwV/x67Kqa26HKnbQeK3xe1GNSAAYuSXRYpG9
OJhJsIKgo7Wc3OotKPPwNCJfgYotwsU1SPXXqnoGyM0MuhenUR9cRb3UzaqeMnAs
UikEGGz/P64fF2WkJAqys2Z6kSu7RCsCMfEl3IoQJSvdwANL1lUBJac6tpEyEmAP
DQNeIycpGaeohz9OaBhc5JsOuIXYojNcFKuh2vEycHLKYqO9rHZp/2q5MN3XqDj9
BcZmW//Jcq5oD3zqjLCZR4ffZYukOo6T6EoKAp6ejmLnNBbhehbvpDBPNb3iQ+YQ
wIiP+E48Vme2a6hifKulET1xn+xQsUfLwF3jnrUoBCcuFxZYzKj5gKbIoVB/kKCf
P78XS3ILAzKdxSrpphm7yj7uTLHsIdu4ncceLnZ9INtB2bpkbkFmzZ2yTzWlBd/N
kuOiGLW9rQ7Ffqcrok7jDDb1AhOoS2IgYj6er7dEG+PGN5SuaoreZ2/VyL8iDJ3m
MgIdfgHTC2amD5XBv8weVxD6oXT6MTLinuQtUftW0tGakS4F9tr0eRvBS6waeMuQ
NVtSuOJni59p9IgnAlHgInMn93LUovqiAt2uUx6gTOXbXKBBwSn1cIUFZaUTlggp
s0DsdoBRYCEt75WLfU+I6Au63JPFH9EBikAsyQmo/cpkLDe6kcml/3CeQWpT5PU/
4vwt1xnvKK+MWNtS1aixXuzS/lHEEZT86Ya+v+PP6H4xQlygtelHrjMxnflq869t
HUXuVNfOEDWksLfIHnBP8LMuI012m9CYD3el6imLjsmFyBiOMeKUV7sgXuoso8W4
eTawhNw85IcuEuzP2nUgb30QYtCgH5FbzClavsiwbgdmUZefBCjMaDpWZFXyCjx0
HE29xYxLlUDxfjK/iuPVSINsrLO6Dq2zjiFX10649oS7hH6shVD9DaUICWJUCTWJ
jmb5KLfGxCBY13+vAFlVaYWN9HZQfhgzLli9rD+OqRHfyXXyhq0zPZij6pfw2nlt
xXuyMfzQ9ENEIeoahu6NlhT9DuSeVYOXS7GlaLADqho0rN9hRAZ28TdqUiwygxYI
aIIQTdbse9xV4duy0Yr9qfMhuyjRhf4fJfRK1w+COwg6D8zTWdgIfNSqQaRQvlZH
cL6XAIRMBGqpz2Bf/rgd82N2ss80WdNCNGY7wAKG1B0WauVCvbybtnNzf209Qn1M
v4/BXX5TgNzTxV9QSr3WlF72Wk38k9JTqqc5P8Q/6aNBu/0aEUWQu/LTXJjempUs
bq88T+C78SdIr2nZktGw8a1QESrwwKhVxd7lwKqscvrQ0iyvfBIHVw1NqRSEMIzP
n4Ox3ePR2xE+5//WxtB8PH7G+4Upr046vChrdQX7WdiHUyf5WDIDOaDUQA6nkTbv
3g9kbhr9L8uVmF7ZD3Zf52NyK2Tmt3C2kk7Ewzv5tfEg3Wnnv/Z+YciaYQsKkvG3
ihKKkKle3zyfbQ2FJYKUmCtGPbuIWfXhPlH4FseUhmS+xNitsNvhfmuMeboozduD
27DkYLYNEzRJTQjpzc6AUEIoFnsv/F6rZajT2XC5WOUDcrMGwh41xWgepevUQ8Jy
T6P/q6/oxlk2IYLp03YgF5Ptp300lazCVWMREtVxexnKGSWPZytWv/TSSpM7zSbg
SReDIZtvhZKBdNsN0AS8HzyNVzcHczckFBMwEpVCx5WtVyWH8v3+N/9mJP1fK2qT
oVXjGCDnRMW+Wvi82AKITKqKDESRP4EMxup5xUC2pHKJjNcKy7Lqx94Gm1Z+qK28
BeOFsdTpbE9xoXw7wfGx+zKJ7/kdIKH1m09kGUSux9TDqVYdn3mK2hfNJ13qvw07
TpN3/q0onioz2fIHlzqdTol472W5C8TBsD9MS9tkHPH/A1Y0bMYFtJMdEn57lD0C
SS+BY2hLeYDqcY00aTiD6S37jiE2IPorwH1xKxgrL+YmhYsQOlGbCOooDvFtyeWd
KgeacCghFLxWYEJfBQ1EOOi4vMta4Tt03iTTw6NTOoeFtRF3dr8QJEucGWQlgdbS
/omPWBXkxHdqmioy/w7ojV4DF0iZl9VQfb03S+2mHW4p5hxuowxj8/rtxK5oNNBL
CqB0p53pKfodJByOnN0FI3LgVjd5iWh4RH7bnYl9G0m5lqeLqFHcfOjt1UuXCajG
DePFubs1wrK0VeNdGuocqq0SVzM6oAN7PqMHPyz2ytKhXJcQkd0h5ie264MMPCe3
2YW1BvFCGHbbWf/F/SL3ZULAGLNrqOdvVxRhe0sWEajAdCFBDBADzA84h5YmzloM
qADHEu0CTtSPWnS3PafMqltfuIfo8xQHxAT5V3IK8NndNsR9Jlmjj3ePEsPK8x6r
lRyOaWb4pu8MfULTrDC4tKb9yaHBkTjSNy4N0AGG+GmiFm4PNARTJHwH0zgMbRwp
AukpJqWLIuxw+kzGqWepl+upIYNcvOdjG5MDenVkcsC6SWkY+UTwsqgz/H6O+MFq
5gdisWiuo0EcIITZbiMwm3i78swqJgoEHl4eRCPpWEF1xKDQbBRi2N2SFOxbPqyp
ZywIWmgEKeG2hJzVBiMJxSwhiiYy0W+h8MRZpO57ixSHGDKKc0cCrLlwlVfvQ6kU
Q8J1DX3MTaYyLYSr3Z1IIbLOxNUyEbhI79R593ReO6ygo6eCiigVOTCpvC6WqUQp
s1DmmJRE8c1teCAU2dxGP6llqm8EVBZVKTdiSnbEbV+qjqQDTqD1curuBJVtPtsc
Wst6xeFVVrFyhKG8sO5+mD67XDbue3ld0mO/+lNhJc7dPt4ejSDZQhP84g5Xg+5g
RC59sQiyPF8LvjES+0C6PB9HiNIkAkFSE8cg6R/oJ7vzXNpJb7yO3Jeckpdnjb+9
QTYLTBzU7H/XRwKsk/Ih3FtfuwC1wcOdVPkBtC/D0loWdkciFEX3K6mpdXqGSvsg
Ml6eMXCDasLrJ239fLSCQbRu64L0H8aVRFuNdy9Mb3pQWvgdtM6+fuA9SHwh1fsH
TE/2OGiWc8IU8UqRoesWub9VAqtmqq5xh/hCQxDjQCDk4IXu/mbVb99IxriHWDC8
IHIrlGXYlmog0KkVWiqMMsl/rMlWBb/bKR3DRp2jvPNTaDjuGZMVb4g/tVUxiZVV
GT7WCLcUWUK0nVIDtRcJtoP7+49fpJkjOaHydviMrK88s6gggelFQIIiD+dSzmbH
zNwzhyHcJ4tgYu4VP++X9nKVYQOJ2lkDAOhonE5wPEaTNw6jfj+XAAruLZPyaFM9
NO8BeIwKuLJ/s+AZV4gEKSrQ3iZsAC5N7SbWJhp766kZyRbgmqWbj75ZpcYeRDp5
+CvCTMvBi4ckRUc3TzUEtCqAd9/HZXgSsQ4cA+hFtMPskRlcA2s/LjKQ+w+va6i+
jaPpKChpGOiq2AOZyid96XHntsnLAi4O+7vd2aMMDwwNmlIVstMhPyJzQs/8oYFQ
WaNoF3u3XcrT7DBLo4Hh5+T93nPBJ2gYaGFt6OAMBN9s9rVg/04Vq0pZwLX4JuLY
Sun6ie+xArKnbZtBAK5QMlI3/h5gnoT70EU5ixHuBllLT0evsHzlNSbKccOv5T4P
Jjwv/fOFtCz9UHZOqa7UHKQFvw/MJrZahlw705z3lA2n1m4Rl2Ba+Lv5XHm2N4jb
mGz2jkeg9BJ+gGu5rtnRK3GeUZwCLjq1RSyxaPP1JRxaCKn6r61mGdmZa+uI74UD
OaOqfiB96KeaVyKUCySpm+NL8vO7nZWCfzjCYhpDRMGU5JIh2D7gMhfToBkWxX+/
MSSrgZlAhYxNCPJ93p/JzLAuUfoK/E0FaiDtMpKKCOsxXS7k2cs1gTarNn7hOp/X
8qyqqqLA+9ovwF2WRnYmgAqvVl/KWl7EC05co6b2W9ZAVM8xCFgdlxcKCrCuOAPJ
JPMP1ucM7gJwjIuMo8EYDJsrq0m3YKtydvDjZrYsHZNPsLdYDkXVjclhJT7ASR77
6nwD2GS6c7hvDy6+MR8jFmhkIjdupnwBdlOtZNYjPhf24NYNfRhedkxzrOizWh8q
lH/Hau1w+zSfjqYY1y0eh+x8xIuKXYZ508XrcOfUvUqJgzjAbYKimXBzVf2jSUBx
6mBXo5Dmxvs82QqXz/FcrK/BFh/9ltLnlF7FqmHxQW+acKXmu3ktftz226lNoE8l
LtPDoqWIwLXBs4QdJmZjRI67AJ6p0uwM8vfW+xSDHvAnzA6M0UHlyrUmPd+XQgBN
LIoiIDK3kBXzB8mTpPtryN9L0BQs488Ik99o3JZX/d2EyHZuEqePq17zCIbvCefB
+Zmej55IQRIYUzGvCI9t2CinMs2xFhpEvh3H0UM3gbq7/PZMKh6Mebsxd2GPlKJ4
XrqPrwincFWVcCJWX9TcXtfHjjm6qOnZics06K1I1gCXBsDIFdlOxD2x1dMGc36K
RZ3OPPvh9WQTRwLERZT2OkL5qE2/opB1jYVzhv5AKH1nKFYdPta+GHcZtBVNZ8Vu
tHQ/HSIrBxuRyrNXyiLNkSC1BRDP/sGd6Y5Hh5vZySLokw26omECO9JiApr6PBaQ
rCp8vdM25FDrwh16NgqocN5nISiQ1YaHgcVPW0DhW1+F6ozf6bpjThu0SI4bKuI1
0MN0J34S/k3j6Ory2+/BCijbgQ4gCUxt7HfyD3usNbxk/NWq7hE4IveAQtixKi0k
+38ukYuDjTMtUnzHpMK4xItu4pzyv5KQVo3Iu4zBr4lndEyz6GqoG40rgrdPDgGJ
XHGBBxga7lL0Wnw6Cuukd8PH2K8NoTg9w9yttDeVPHeu+e6Og3HJDKl2JCM5dHig
ysxIRW4DkyItc6n4nloPUJhbflae7bU5iL1VruB8x9imG8WSDa7XKUMONC4nxLbE
40KkAyjGzvCAzfOEnHUdjTyCqQe10RoYv4VJAILkLXcLP3tCcbGhyr10Hjxxttpb
yR0r470VGdP7cmDjgDxdeXxIJLKW6OodL11Xb4AOKgkSYARho1pUFJUzGxD4FXka
AjIj9Umgkd8N/+gFk+Ppn3W7Z0GmWPjKnuaK4zLCpXqi7zFkLXJ7iblIJVVcNud1
fROkUgZg2QWp7K9AAnYYma5nGNF/FvMh8wXmWRShaTdIV3hasmcb75DdsLYROcrc
QNVttPfKp7CCjfOI6znsWHbWoIv2C11jQqubVNoAebxu6QTFY2rBj6xOIesQpZgi
H3R8RWZN92g3JXsdrAYLyp6wkfSTJQqR9sRwRnz7gmZkA0CJ7A1UvT3Bgb/bM9EG
4ET8GFi6pZ0fVQ3L5s5CSsTsEN+iKOL6El4pU/Ey2YnCyZ/mFd9P2ma3U9qp/YQy
YoStIii4V5Tm38slUlhQo5sepJR5iMXszCmm/NM0BQ6007tvNPIu76mL8rq6hTxx
g8B8Kyvh6sVfkcFojXHHgTV9xn8dBlhfaTt6wW7syEMtaDwo0p4rxWMB39V6MLEa
zu6BaQznUAfjOzhdKFESmq/hoQR9XZGdah8gMwawUz7lfepDAH1fvMcKXa9W4L4A
7lObQS9LzgqR6tO2aUoOrihAkzFgRAOYMvu94qhBAidHfpe5MycoI1ZUcgg1YZ+7
53bDMDng8fAg0LUYQs/KrKHdo0CMI0Xyc6c7/TgCdS0KSqYY/lG2HLu6n9nPzn3o
xJtXy3Fv89f8F+GUKpelyhXxPDM29wmpmfay+YphSqoqPHcEkFBimT/1kCbF1jLR
pLlZYXmeRaMHxw1iHnZPnCdZ9/b/yoF1vyLewKcDYfA6Hj4mbOhUWkaXb9vfob2T
Z+b8E2gDslG3LOeynEqMQ9wTFp9avHkuvp97Hyo2c3VMpOLHDHolV/Y627OgaVEd
gC5VnmQvC5UhjYMpyA1y8w2NcWhOzoJuN05zevkxndDR21bqT1qUjGDHzyED4YhJ
GUMs7RL1imlkNppNScfJBRAzsFPWxFHrFW2TO1+qcn39G2lnefP/RQoAiyz8Weva
CVd2uvu/VVJKJ2sgbew/y+bgUJwyuJM+QaybiYDyrtHaF5Cc1Yow4VoPi+s2DD1D
W0GdtLl47+pHiOcGvicKTMjmV3XoUmsTF85a07uu6nMCTAeqpA/ZtH0cKrAh4LZx
/E9etSadNCYKa/TZI659+4PA5+KDSpYPG1MpBqFJ6h5/v0trf4MbbenLASvE8eBq
ZFVYlBPFBdm/alUKi2o51svBwmzXl1/PjO1VZO4SJq0JPjlMrJ4AcRqAhTLM8y5P
NzkMQEWGnPc3JwCuJUS62g1LCXWw/sWkeaboxrV9nZDRE0ZIIHOawDemlMckpUwp
Av+QaiyG51M/ouFJ7VzFEC0sbzOQjrB73ps9ifsQblrU78gkwS4pmJmVnaY31C/+
xjknPIjJ+bjvfTyJD/kG66iifN2sjzLk3aSvl+8YHN+gE5ozZ1LQKtyJFoo+7L0a
ezXwybq1uGgfFg3JU3waVmmN+CSb3MKv1nGURDpAaPy8IScQAesOcky07t+FVYlm
sbVAaxjyT576sfyjFiMSEC1rO6Idp6gkpKk2YVftmrAusA2h/0wQmKqJPeQCLWen
yxS5aMlqJoXUgYnx2zuROvMy0w4cCNFBZUfUGgZZTCRgbO8+Ylmn8Zlvkw9RamJB
WaJGeMeD3Nu1BgQSHf3u5vPAWyL2WHCrccKXpi4/TgwzJrm8ly97u+5oos5dURSh
z1aKVMoEhe2TINzidIUWnFIRnzvECNlrb7b7hD2nl3lEC7wOMggCBRyy5gzE8gZ0
/u8ihyQayG2W++nlg9z4xejv6aFhygsTO8SuFOxc99DMdWnIRATLABg3+Kn7NWi7
oYUU7pS5r6YTvTQXAmZPRQ+bd1ppYUNx/aVphFZpIV15fc066ML87q8N5aNtZgjN
DMIH6It32dKFc4wm1h6x1SbXZhcZypqrcjAcIIkIo2g6z9Vbowdv6rrOFDd8Wasu
UnnCuRFdziTjfMDomzKMRPe56iiEKZSEo1I06jKQcotQw37krbBznYAhRo/9As+E
xfhivQt3+KxRXhb/ji9K8Z24UeZ+Wc8lB91ps6iaaWf/fIThoDHEfSohEC4dLPPo
ztvYWCM4VLbsvEs0RB2Vg/U5yEgIJ+u+/Mhw1KYx35pl6X6cAzklDSGk0pDGVlGg
/HE51WX3ypbLb0DWcIpVphs4pWwecfPTPkHqixizTwwD9EGCQeyMh50vI+lYK16q
3AqhBRPHlkiYplwawiSJFxVm0XGJrWURdRmHZV0CJzOsFm5JeReyyWcKRe0gbYbP
q1I+PJNECc2fCAHaKW4WOGGusx9p9UKQV0xScOPcQQdEhTKng2Mo2+r8yXpviSPC
8MLrd+7jmZK+sHuPXPdtKrU1GbBVPU4wKNy2RsGiSAULOhQuY6oWuCUEqC+BS5wr
zhm80QbvSafg3P8PS4YLvo33KmRsJh1oMQedPCF4Tt1Kc6Hyqu4HzEMFN1g2z2Ka
wiNqbki5oduMYa3jEOKzMRyMIcKg0V+gNMQAx9F3F83Njre99LU0oW/cHdeKYjWK
W9ccYitcC4/V9qF2iToUwA/bl5MUq7CzcjPdv9MMiT5Zk7BOYNbZ8wzU0aTTN0/v
9EH9a24WPUhZakq1Y1pH31i/XNNhSzlAhUOH5iVbYAXOaY+UO7bJqsfF9dWYWGlM
kIGqGb+QZTOQk6NMEirTothICbfD4I8fH6WfZhJqIznAO2ok1y08976ZlT2+5VE9
a82slqk+reg7RUHoTKInh1UAHA/bbgZz4cObra9q6nVTkJYOkrHWZfKQsTtTi1PG
9FGfHJZh4L/DmcgUXS0KBcj6Ov202XyFd7oQhDlDYGgspBCfOx786yU0U9YgawH4
RCLQJXDekYwJpfm9eTZ7NAdj/CqHnOu+EOEP53VlA64XTm9LKl9mIL40kR/gixds
wQEVMx89kSanhzMkaOPEuu9KSZBlm8KydfwaNjCVDC6WsppsUX5XHxl4SyfCUz9b
svOHpTuF6t98YWllMjy4oZTXoZOVOOoLRFgIHzXfXqPUmx5jgfu6RrjfMRFtLeIc
j+dKNZ+PdZeoDlB377w5F7MatX7V5udZKRkyByw4RU+mRxd35f1tAxk26sNJ2cE9
xM3Xxm/u/LwOuw9wPTY6nnltxCuCL22CVlW5NgB1PUmJEu1NUhl3SMu/wvqmshVy
vrMSGQjSAXsqeVXiLtEUmtV3GJHLdoJmiJJ2iARnVkwAYBtkG3RmjF2M5hqR4Qr3
xj9wVMFWuqVz685leacI15NS2WtTTMiXPlwKn2WdOG19vA6FESGtnThIeO5V3jYh
ntiJhrbZAkQYnhDHZ90u8XY9PgbjiGOSHaSrtPPeTnvtbBr7PmARBCwjTQll6YWh
HddPHTnmXiA8RNgk4zje9tA15NXBRKSeCadkQfpTEIMLp5on0NiCDYs3W6aV0Gjz
XrA3/fn5gcAuFPYNutr6f2FFLspg/B5/+z291N0tCGFDkIXMCfjbqQE2nciA/Tux
vwNmgk679TMqz+nSq/uXUK7/I/a0RqYQ2J/g379lgB4vYkNbOwlRwiV2hRfiGj0L
oKHeNuvm3lzMU3Rfa538icMt9Oyd56Q8deIXbpqp7PYpgi670/po9OovtWs1hkFD
PolvX4Ns0AouAvs2niSeBaw8KnECdgd/hIv82D2zOMNtZjUiOtShUxc/MAM4Ps7F
j4oIrYuBe++R23ZFB+OBKo5wgMZVhe9JBl9MGNzEUs8C2b4wYiKjAsX2zJCGvmqH
qcTrEztCKfXVDyy8W2OSCX51rtosetCbgee5OuIh+fUl25NhPR3cXsIyRkqxIHbK
7iEH249Rp6ZVr+GmqDISwbvAW/dlny5I0dRbZiq9bqJ+YuZV3i94xXn6p25PgfbL
7Y1sQHPkEb+RPTpKz48Xvi+eAeSwK2MHdb6ynTmY7xAGcr5+GYbyUN+i15bYP6jm
wTbOKeemhSYBaGDGcB0BPBkSryAvORmgCgki3drh1hQgHAp197vFJwGKlW/qpJcp
rY8DnKuWZCL678A8tv21w5l78qo0N4JbS8HGA62Vbg81ne9GhYRqxyFIh7yk5vzy
VleacjmtPpVuvkbMHpq9iyRrWNABPJKXFXQdc3hj4yhR1i1CYyCAwtzwW4ibhaUp
5+BwxCrnnRKUFBghtWkDJgeeQkAIwE1gLC2ml96u4acsqZ3EhCnKDWqBzwK/8pzx
qrmkja9wrXyh0aduBlqjNUEmXEsbgEjBdVvsteLGJU97c/T8EIPZ5R3STuyshEut
ijgdU+R/gmnTkmr1kgFW2t/dU3Xfw7my8gWkURJdkXBw8mGC3VLquMi907T0pvfy
aPuJbU7+hEozdx9xskE4bHzUVE4A2z9fekiCOMnqoeUZdn6D/sqLroow2WjIms3X
qrnq5TcF3d5gltNmhZyOVIemtgOjUNVbdqY6PeFtrlbhk8ETh8OD4YF8BT/HlylG
lWXao3zPF+wwdkWTXrXJpPneB/EWl+uCF6D62hQjWNWnUfSneurf0fyArj54BZSj
oaEKMarlUh5fYAau50ybOliSLH/B+bzGpzjbpyguYIRfvDsWC49ZJNHowkki3ZWF
0G7dGJ9qTBfaA5/CyFzRLYk3YGbNigpVX51vSOJQavcjSFmwk2bamho3CzGDvJOw
jhaqHoa5eBE+FmJPtdvYS9VdVNWgbMCyrBYccXfoZgelHoRkK1lNLHM7ekMelmlT
z9y2kcCAvWQt7Srll1aq6ctWKioWFdXkhyRqeftxuwIEhzqSVf6WnlND7W5dkv33
aMMrVmCuTGY1qNVE/HfG3sbJtpfZmhX4zKA8dhsZFXcA9qm0jSlfa61bCyIEfldu
6qrbal5WZmjz2fmH6MO7Y3XMtu+qkTe3jXvp9BXDk5b8IbKRr4mbgFtOlibMG8H8
3qOhxKDWU8XFRHsiAVjWlaBscyV+Zu9fUFWyvBzMi6MEIxR9GlNk/UVf49QIUd9+
iEa0adKz5tIz2l2VpLaEdH6a4Gs24lPIC8tedoBny/FanJaUdwKedgdSaHim+0au
9C0gdu6rcpodwBjAYUiLNWPbEgCLIdjM7+1X3y3wnlznbHMq03GpTIkyKumPKp9X
Uujhh7YqKO9pWU58iEB1KVqkbD6Dcra9p20tKZyQOmHf+gm+scvkcVeLMAVLF0LW
ukP6AMeyKd8q2GQ1V/ppAFBFXtI6EPwFEMnS6TUvAgUhYHmobOoTE7L8pE7BzA/t
MDdX+TLzEqs1tnh9b22GKgqsuPrKTfn64kAZtsYENUJwecMwmiJ1n1jf2JOYTNdY
7z7utg1470la3rIHl1RGhaDnN3CEAc3F/rfluvWH31OADVb3Y18ZbxoauP9eWvtL
bYG9I8SJmheif3GJ4y/KutiEsTdZ8tBjnULf9LuseqrcDlKluze94pDQjNfvOh3f
+W6HOeRSBFJP0RJK29/R++RdlIHc7OTfNk8zuSGVqoNGZIVpCh4yUfG6DzMArWg4
RL7JUk8hmaUqF5x7eRqFdz3aQVMibRqIvZ7KzwmAhpK/LIobyUBD38GzIp8dpcmI
e/bJR++5FWCCvBL6oN4KzxQpnAyleyX2xQq+B2xFHUOaNJE7mlhsdryfn0iX7748
FZbAmm5am3zLAcMIblNnGKQqL9o6Mqph9rQktKUKE+Auhd9bNE9ZZywsGaRwRECt
P4ovg4YGb56Au04bveWR6vA1jYCmKo+IEnMCrR+lk/gx8XNomYKhANraRNWQ32UT
xkq5DE58obzHFpgrGEmysIqhuWg/B93x0Js34DTqZsfSqNqGzYlHyyG8JHsFvv+H
e1czqIcOBHpNqr97DnShjPyX21vrtxmrNvu2b1nsPMN5goYQLqFhzjnpfOm36tt1
Ru0yEkFqNBWXYf8lUEiKj3+ABKLLcx3or5I/lI3vMi5VHI077CK8u3zyucef8mOQ
rvFqHFHUBTc/MLDLPXqKXDdOfTbck8r6HPOmW1e8dwc1OzGMIJEc/fTPS0vYZZLc
hQSCp5VuZVunn8GF6JyEQa5DFHFZmVPaTt19D7rwN/n2HtBxnG8HVJuuMQjB7IZ7
7C9G3WYjfAYiIHtVETOEIVQuB2Z4A6d6mIuJ5t59wg8PY194KGJsGzYFVqWB5TZe
2BOtfDmpo5rlS+e7Ud12GcpiSwXa63VMNy0L0G94LNwIpDIzbwkYwyqzOVRZH0fn
dOeXJvrJLZ+EOm4pGV0Wo64FZ632UjZ7rG8aZXrdT+Dn/etroDFKJn6QwThmmX0F
+ufoEWnXBCS0vFWGD7IDhkwApOAj/dk5rFvfmhL/B5QP89DP9w2N92F8z6VEiXrx
pJWXbS9ut1VZKBiySZ5SrV7GfhGS+1EhqrGcd2UeZLp9nKo9MWHTSGl9vhmTpBVD
dyOdiZkiFpmeNdKbcYj5rjRAswkmAYJDPUvntwquWY9mYGI61CWckI3SGiMeYt0n
QPUA/r65td0AiU6v+KyFvKf4PP8hEo9IqT4lLVja01PRqSPSIGLD80m2cIGyRpDc
unDHVMBx1EY0g8YQ0TdqMuUhqTumBaYBKZUbataqNryxHoSjFpaoqtOZLQpB+3bq
xYQjbXl+mgSZ3nYFZZ58EFdNY2i8ByH4GjeY/eXAUOjuIiUfZKyToF4qI71raOwf
Po1R4Y/n0JL6GHpmSFkr6PeIOZa0m67CbOoLYSRSONNeYe6a4GsqChL6eAFfcW6A
ZVVostwqOFAoNgwSJdQ8BX6EVZsTOrg46RiFfXU+vNnjgXIrY1iSwtLm515ivseJ
qxuTYzfRdxYi7knIVzXcDwuMZnem8gWtWN9AiY4nrGbal2nSlGmpZVZi1l7N0XeB
l1h/UMwZUJraC4cnruiYVtNFgaKiGgpGa2tnZ2zxDp/DZ67V3HKD3q8eLOrPyPF3
lzfDsNi1SZh+oT0uND2/HXMxLb8hQUixDphLNKnAli+pmW9mPDG4X83J51px07Kh
QBXZaPsAU4yu2u2QC281SRls3lKxyeCm4vNSxfLJ9DXQNyQvysI4YoF2xah3sOuD
MND9SZt2kksRt18nbfZ3vIsrSXhuh3ZC2+9VshbEdtp//885LfC2yXz8r/2JVWAT
yzGh80hxWP7rYEaZZUhS7mKr8LMjHE5iUwkCISLZaLG0ZzgFk1k9Awc29WLQdFoh
f9rH0nB0sBNYvQZpmc4J6idBmngq+Pkcep1DK/q7dLieKKuDPCij9kA2o6l+GHeH
Ip2kYFi0MIzsQh6NVqWZ6ibw7Yv+RGWAcE+dLNghbaSWhCQHMQHOdvPv0AqNvw13
WNaAfIYl4QAklobWNRXpSe3kC28M9cyT5IQoRrFVqjcHjyPnL633TfsstXcTFCOq
i+0juJR09Hu7M2mDPjpO7vNOyfYcnXWjLufoiloCVreD+d86qe4q/MU2Q2VQ2msC
d6SbaAZOPPJ2GyFEdFrr1Fr7cfD8IyiicNqbKkfCaDJrh8TBJ9vcFuzsECKvUWqH
/wFXX+++S3nQNk8qfK7WjMOask3H1Q+WQxaQH1oyMg6a8dODFVuQ9eCPgjj3hpZ1
j4KptjbJL3n77qXZ5mhu0DnFVyOIw6sV6cc0r8Pb8H16tK+PAILsyhlaU3FZxVjz
5iwbO92BqbO2SN8P0yCoSMvImkpUDKnGuENrTG/NKoYX3Nz3wMuUUvFU2+ZI7ukG
xN2JDoiCdotfJuavrocq+OmDQTNt9j74xj/jv1lSWM4AGj1pZakYI8yBw80LFH6C
KYj1D32HUigik1mU9xE5wuaaUMDGNMPezliWt2oJyj/7E2koxaa/ho4hx+GUgpNm
2tEICqiTU0tm7/J6Ecq2y4nD9Ac+QgJJcOwRwLTHM9r8cmo8avyH6DUWQ7HqO7II
ijRRh9fx+etV4m1IzoKV2vwbu4n69DUl41JkXvR6uQnOfaD0ENEeiI45kNosI0gi
6NzCdpQKCi2BUWF2XhjNJR98Q8Ym+aK7GX51CCGA6/OsaHNXl6pF6ppSNVWOT79t
e5tVnfqhocTd1X+LE7kVINomcJckFQkk7DFfT/+C542X1p6xx3VLTQ2D0+f9lEZj
NsWbCFxc8HJ9IOR6ZehzPp7tapG//jfu8cFNrNsQTFjNexL3X+EaRlUQ+5Md1bPC
Vetn0ynK4MgkYxLaCnz90WdvoweucpL0yOsRQwWDXJhf9XaGHNrZGMeqQ9LMQSKX
UW6eCO8gLLCJajZ2Tbgk1YThZrcLrUDMtqfzHMS5gxehFP5KoJoUYsNdj/vYldt9
i8PkAaNTY4v7bkKPs2XOcWkMTGSITy6rJ3DKfosoF5ki1XjZdOaNt0CCbqSpJYDT
WRN6mzs6UimHCajUiaCnXqR+0h1MbLZlct7WtY4b+Vgcxx02rR26wDrrMbtPn8Pg
+Dk59ocdRV8I63VORB5zX10PwwRyAdiBYAO53DoOz697aCilFWUy46Vme7h6B9Da
8+EptVmDNgHF1YNVw8DQjgVKCICidRloMxU5cXZjsprOLd4/6fuk8lDVZc/8XKJT
9NGjnZ221iKiH5V4JmRZ8WV8eEH9ZLUwJOJdMlUmKRc23V2VxJV4juXb6s85QBp1
R07BIHvlmzE8lRyFMmya/q/Ua//2qSFwXwy9H657u9AQ6Wo+1mkKJ6h/0zcg4twY
mB8bgGvBcDFEUg6GpYBr8ehEf92iU+4XSleBnU998SppPcHhQUt3LTfDsaqg/1pe
GesNNtRKIhzvf2jSQ/pD6d8kDFJhLynd8yYaNkkcv4E74w+Z+ZzDmfmg9j3BDxLo
ose7QiR2RzbOK8PBh4LJk/I/ucxZPMSF5nGmKDGtXb5N2fWhq88OIlKi/mpuvaao
fTylqDWm1w2hacC981XgYHkM/4IDdqnxxlSa3/TnQr7Ze4jUa6HLWyGiWLWk7CAI
uSlwJykYBJVI5XPfKbZBv3wOemarCT534bnhRqvDui/jGptWZmSO+12sdMn3SBkb
LQWKCFURocf3koFoti8Ssiraazl5U0XH1RrV7aGnWRsncLL8N22gToRikfDMDO4I
3SnpZ1+NdzunO/48uhh+cJaPKwbPLC5go099laVYixnF7hvolpUeJim/wwB3bjAm
APNJPyuGC8mpK/D0Zaemur/APmsC1DMD88hoFXm8ZpeVr7MQGaeMEN85k2gvlrfw
6bg3GXBNmNR5of39FYo+bolWn35US7eUdN7Bb0ohdgKcUmCSe81J2rgMeeJCDai3
NhQSb2U1Ppfd3AUkj7b3lbZYXOa7jGZjcVwQLNQNPu7rnJK4ZYCdZnNdDtgFlghI
vnWCDv4UY0I2IcCStzhq93u7Us3Fi/6suAHhrYtrA1LPtglzdeQSC6kQHeh+SwTT
tlPMH3+3hjmN+XnOWrLGRvr/EJK6m2MYUjaHU0Lp8seP/hSS8VY1PY168iFsu81l
6Ucuxup2nulVN7iQdDWGC/4qCn3SazyB5MsaRKtmg9irsaKRXMp5HrHzovmTOgyq
Sn5mIJVtZZwIyYuHWHvdVqd9R+eq08L9LPnfFZHqCTPV9ZV3V9oKIe3c0DIE+vSd
aToMngTvc6J/2HZ75Y/zJ/825zSVqPsj6fPYRov9uLW4Qs7ITXknq8dEcXv/2Ch2
R6ItRSUToQdVplwuvaa1Xv+A+MHuuuimnA27KmVf9LODzZpsLHeBKmXayWjzaJOB
l/sEAqZ+KCwr9xZ9QYi0Vv+fBo2perrzn75x7MWpJhUXd2J6G9ZkRLSVQ4dJdPbf
QcDW1MLfG8IUODgOK3jwBa/QU70t6WY04OwxXnwLIM914dSGqUvgoEesoRW9WwWQ
B2NzfZ8zqdJfXGOfMIm/p2vubLmfnoB6P5V5S/WRBG20r6/E4FeEHt38jJfdfdIM
i7/5mdnnWc6o7epy0oaAIF4qtl6CI0zsIjFuqzH9rgQOa+x3t9Zz7HikG7L3LnV/
BfF7fnVXtH0qfzuJAQUGHsgRi4vgS2/10w6j+Qste5ztYw4UpOW+zupVep42n8Gr
4uUZ/WHKHfdqi2Gizl8ycMeopFoqWGUn92KJcosx3pxDzGLcdh+Yu1vZwZ88KDD9
2s0oom4p+DNTgld6C+wj1Qj7wjzOgbiJQTqcvoXnvxa2aEFSWsDObUQNOyZHP630
KZ1PFpmVTdLG110pzFMeahhKRR3qrZPACnwVjmFOH8XQWYgjjv5pcVUqVw3QiZHv
iZir4xeHbDQLMQiX7ZDFvDKZWQayaz6ILZRhQD/ngT66FOq74xeLlkjW2wZ6xzA6
HjHbF7hDbpweOMMs9KFfY+iDc94QR2BQ7uj2VgNo8g42WI6qnAYoG5rAUZpjybDd
+l1l3bWqkzxwH4DI3MQQtSpGUB+l4Z7Pd6pk1+TsfQbhgQPH3XKy1EFdrAxE/rIM
xilqpm/EWnKbIxUdkaQr1608L7NDYTyU9Cu5MSjvijy48yt7TQClP3Qub7NL2Ss5
7eq+VrCsVdo9lCCrIyRfl7tmkXevnlN8QLg81ueKfjqcaFm3WJ2LO0t8fv6Slxgb
mWYiK9q1rAT68UKjM8yjfpHQBocopTZHZ0L6Z5wrJmNtaltFyjAWv1A5GnP1fKab
JHXqeBNwlfXUYmPWva86yCVFKlh4PHjfUGI5KVJ5ICASSCThOPl9bBKCzQtHnSke
KugJqlNx3/iL/38fPM1yknJ8v2HkiiGWI/sCF2lIdlx1s2TGsLgqFhk9VZSCpH5G
8WaZ2wZxu/36fU+hTsdXzjjXqI0iV7/nyhS/z1qg8bZgLLhrc+93scZFPDXEjfNv
7AwSTmaT5kfz63bLlEqfY+jwjNHjKo8GoGz/NWvo37qY2tfrvXYNcivE1g0ZRqGU
GMOtK/CNJ7BsxdslEvL2wa5wpqYQsZV2oktl2bc6UJrmhh4vkknS1yWdlp5bdGKE
JmpdHV/z2+IJYHAF4K5EWaV6+nTIVEBJ4ASWYD/n3ctLepnqK1zjXZ0s28/BqbMs
MVT+4jN+HMFT45J/kxtJJdLcu9iFWFUIwdrIn4adgRz/58JSwOAy5PZO5WP9QzJI
Rxpz372W9wGmXlMMhbL3+CYbszAQuVdbFiAgVpoxqR3ea/3lWOIgF0fie1PmF9IY
KxsjivHusSPFf+FnjWYXhBXYLkHeaMkGV9pxkkanm2Ixgom0r+78XESYqpeUBhim
UANiEwfLLl5/ir3jsDk+8jc+l+nITshCii22B1sSj+Ta8NSZGiw0aSFYhggz8TrO
7B6H6FHBOxnfSE7pgJN5RdvyiLeEqxlV4quY1sqzDXx7EPR7MFgwu52U7uK+tEwQ
o8Z96XLc3Ynr3Ehpp40M40Eaf/RsFCyHKsOr2u/Rd24MeOAOHW958LQsS8o/usRl
kqg0q3BI60yC9BjR1PvzlNYmTH0EIoZx/g61I9A0w5iVMLOLcakHGcmLgnnIrGoI
gKCTPZRT1uUEHMxiLt6lnMNx6gZjXjbH8BLv/fuIvykwFFuWqr02bv/9XGymXQfY
Xf/xS0wAhxAz3X4YtheEgpLbau5XC+Le4GI0w94NUyu/H222FWeLmt3Es4g57+eH
6TAtl3O5nt+2NTalDbov30RR+ZGhzdSTHwb868DoPaNEs7dcc62QGcxhSZ9XEm9W
gbF4vi9Txzu1jWE/7LvCVknh7R7rJl3YUv8xhkUC4IBAzCmKnNDm7y2EOmf+HVWV
HZyTVXl/2kykb4Rcalt8gMbwvQQbhBNM45sBUFixJlsrLrw3eRC+vhM9YylVmoTO
bEMHJBReu0upOK88sI59VUYMwE9VWLkgeKWvJc7hRdGnbkfR+ZItYGdz65BUUrRY
y6dPfbpyr5V20Tq7g+mfjQqwztPAO6W3ynv5t5Bq7+ewrdCz+mm+Q59d2QEZQxC+
2UA9BeDBxJqsppocUxGZKqT237pdSf6PtjX+Va8gMED1WOewEHEHYWk2sQq1RJWV
pd3aXlBgreCt1ZG743HMLhWHg4jFgoSl+o0CYYLspUargXfkA16n4NPDWeB/mB67
XzEFHYxqKN+enchM9A0cpkXy0uN4gOAPzeBAZCDgTtPHL0p1thrwqZVWG5ejeOQf
JKrBUS1EfBzq1vgMZ69+oW8yjdwLWKdUBxw7SVr6yphvvc0kH671z8/BGb377EV0
MGhqP2NbQ3HcO/Qge6T3XR6E4JJP7I8KS4DPGXY7QXIKbSKUVNYxLAr5Uxljjq7T
h48P2pOrsF+zzJvKnVUe449mV9ljYpZvWmdiOtUZHb0Hcj90rKGS+G8+h7rfmEo0
YiuZL/Vp7rY0ye4Go4chAmmegZliJqwXVcImvZtcYz5DUhB9D0/SgO/cxVjDc4Le
5GsFw/2evHY3UpdDXLSusnu7D/rH9WnfVH0iXH3VQkw9jtMMgxEITU6DBHADnp9V
tgMO2HYf5p+NWmsZYCM4ba3y8ww3o9Ilu8HKTRJ6lckA2ipzUFxStbNWqZYmgDfr
5siH8IgyNqCnVdbBvlo25sch7vCnn5EsaiAALexWN1LCc/Z6OMpkwaLtkASvzjUe
OsfpsMPhpExNBp73jh2dccrLZIGu9vzkx9vQHFKFKwhv2zWftK0A1+4uvGGrQ3hH
ND9XyEcNBXeZoNTWD/qP35Ka41h9e6oVqLu1Qg1eczGk+ro6PFp+QfyxVW98czqc
UZw/qXxv2OIM40yyxe7+vF2i0MNYYJGupM5+22alFPmF7WoCDPL7+fX7l+wKj7sT
OlBHVxPv0kMsBB667dQZ2kwKJCkqu3blG9QoS5eMvCjy10zzspkXikzlnrqXC8YT
6fwNqnT1Cn7UGeyNJp6ysYHMb42bQSGZbPv5eV65PRUIbuZF+pFxX8N8o0We4HFB
YPPB0XAt+bOZxJdYRjfWLFUp2dG2gcxOHBvm4psUmu/6O1WvbQCSXuznckzU96gf
35OuRS4ySJ+zPfROkOwnbNBOkO57gmEk8TW6x827fr0mw96HLq7+CMdnHgwwHsFz
BSR5kr0M2CzZSz0rDNiW3VtFHR5e60hbEm8ZPNmWzHk52I223QCvazIvi0fnCkLC
yfT0s1m2sOfD3Fh63MZ6dr+eF4GmJ+F457L9QCQV3PO4Bc2MY4FiSNZvS8D0erXF
4sIdvp2JFsAj2QnZCFd1lg+hQzleYqgiE0BStFWqpsZGF8QUK3PahFU8othdE9Xn
yzpQJC0nUWD3aIIlPwpbekU1zejv33yUzAZAOEHVxOFr25eVCPl3LMfSQir5N6V2
Jc+moqaY4n9mclOFZFsDSWfTv6r7teXXASg8EikbS+5OzjLSEf7zxTFJ+4ikrAmf
c3fcU4Tv6zVdcSLho+VXMXjEl8A0sSFdTa9Li3dvrTc23ZjJnsV/sPjKncD9psgT
YXZcoutW4+L/9fxUdeD/Tz7WTu6YQN5nlNh7Io2ExiJD883LWqGFKMPguoTqZtPx
HNsJeJ+XBA1rHRgtQ0rhdK9KbuXkqX3guQVRr5kIM4qVA0xSBWVNsfEH9nslA7fe
2JHt7+8DoTrpo0saN2cP4zOCFv8CDBdnOhiJBbdJrJuh7VvOQp7fnbAptn9yMaJS
xIFby4AE3rDwYxTQ7f2CgzLEEO68rfRKAELb+eBro+c+oFSgXlxe/qKhQQIj8sDh
T9213Dk+3nz2uX4W31Z9rL/rjCP4udAgmeriD0CAeJd/bcD1bl0BHd+2vTegn5as
ja4G0C8lLclyoa1q8324ceqpLmxUH63bLDlv0u6OXzFzT2yOKzOpCIkPg5hoQ7+w
Q8AU7g0eDMZRak48G8MhnT7LaOpu4/F9uOqMk8AKbMoRzcqdG/Vef0sk3DN4XdPM
zC51BY00ATwEeyew3iWF2eZOviO2OLjL8L8fL8PPShYjOP1SS3cPko8IM6MwiAPB
kdKlSF7AM53H1p0eZikLBxqxNmgMB7ULzC0R1bgwgD+BSaMNKBLOG8OsdWxYDlss
J2RyTzCtAFdfQVTyKG5B1Ou+Q6RTHw0JYoV1CWj38AGPBW3Q7EuGTpLLjT/178gU
ML1q07Px/x4VWNDBaT40iVizrVmi04BYd5GIWZy3jDPnuDeYNLeOixRhpnURWRoP
zZnxhwk2WtSCi3PM8cpKB5QcxpPEAYHT65cs+31lZGe5EBJxx276I8xU/dNlbiKY
TTBU3FtDYKKwLMXwXfTo713F/KG6TCsYy8CN/A7hM1qPlNMcagZ4ZiRPlXa8z4eU
5ka0S85HiThja1BAicqypLJufTJyLWGvxqxYaSNLyck5QJJDxhGNjy7LLDQw9Ey+
JVyRt3wXA+mEPr88ueTBp/4obXTVPJ//RnOeIe/OlwSP3ir1PMueU4hkFkJpQBh+
ppFTqLfbM6XQmDBbHPqTv7263qqjy6d3hcTThzYGExI0Qp1oOPC13FD4axq/2rq6
6WCtjFFEU6Wae+TZfMkhwcN3o/KHM4nSLvh24IQUnA1O7urePseSZxl2khfOroWB
TJuGn+MhqUMpVJpTAE10DSMY4f/gtp+qkXFwTU2BI16BuALHRkFxZuJbnceNUoI+
JZT7PgaGtobMB8InAVaouc/+LKh4E3YKjboMa4MSikq/yRx99wtmaUhp2bi2sY66
UMuSsUtUJvk3jXF8x4s5PREhU3WlOPAbQoTuXCyIWtwn7Ky/VvKi+7vSOaPZz/qa
jxP67EIHLhOF/IHaD/eJ8hIoqwrJfWkw4e/ybPDdw+NobY9o8yOacBKWdJtrfAz+
GbFQxXlS0pQYY9p8axeOlbVE3cY9v4z0EOZ9qm1tt0wEVw1owRukKmsjh1aS3JxQ
3ig47atQO2R09T6MBtYlpw==
`protect END_PROTECTED
