`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I+LoKCPcdNoWa1tW2UQ4gmgmyQNSAgcS2fqOarcLORL76miLxb8cp37C/QbrYFaz
6rDntP+g/dM/VpIiCX+uxFfJEo+8FFR1ohvpTOZSMwTq8FVSFwr7/dFYM1YD9MLO
nt/69CEmXYgJL7BroSI+BV3iiBctJAAhLaic83CN8xkxGHw2Wi3IK4xawTgfldZ0
8aFJhUlrOO/oQKM80EWO3ddYQ8RZAZ1DiIvI15/Ctcp44QD0qS3xmj+FL1qmbYag
c9Fmez1/saQPZmsghSm0+uFoehrfJ4VqWdn+08klIdnvWRonTvPpQhevhUcmvu5b
Uvvibxgg+LGEagrZi3VF2HFoT+HfidTjRmHMYA2Zq9dvPhsEksWpXKAFdy8yu7MN
H8FicahChDMWfGsU6zI6lQ6KFUlvmt+2vFoVr+4IjuUkj/Tnvj28SKyyaTizLLaQ
XUUUXW6xkZJOKETWCMZdcScTUSfvkAtRLtXk6OKjmQtJlz7Z11pO4l5TUZ/gMp27
kbUWEndDY/1jGDn0K+djIeWYjI1uoHHM7+INGV8Lv3LB1OTRzW9TB2o9r2n+Mk7U
sOU5MR8zVqya4pV3/ssHl1vbdZHJmz4jLEA2ORwRGAQV/iPXSsiE+jawPV0X5798
48flafXCTvUbWFxEhGDTLDAB6bzEFSeyeF9/eiBXmrIImJy/QkZLKgtmx8VBv94G
uYHPmza20LXT9xdSr3xlKIYXHBhKUvLOzoWMR3S1kVmIyWLR/q0KvFDOqhIu0D/t
1+F2Czw9cNrMAHt7J7nicvSnsx8wQiB1HLQBOEZyMlnC5lqpARSjP/U/raWSZsOe
Y+WWuWB1Qko4JMkma3XP4yse5SyspRZrkDyf7a4Mr+CsHBDSkwoT+dzsmdkWTC+9
8SM7dM7vzH1trIih8kI9aHV1aRk1S6v1sq7YsvFFaqpZWikxxOglbERBBdK59oqw
RqAnY0xjrkkq55QLgaeypAoT/Jl0IXqbcovEzgLFdwDO+T6xtVSs07YENoo0E3+Q
de21ys++23ZtbHx27D+hSzgnHKjaeTvhE6ljjExipJJtrcPCUbTzfABf/c00EADU
uEe01qeeOV1USPsCD8wzxkSsX6CzNl0K2P9b/lH/tbicPB8o/Owj0B5butyy1dGy
zWiH7KA+F89ke925mqnEIWq7mVxFVWfyDcUOTE5EG2E5tPdyZRrjBFSj2AJSsBpf
MoIeZGRRLcY5fu3EvMBT6SkAKg5vQnW+KOyZ+sUk/bpixsHuuPCOAJfZ0gYlgX80
BCMD60AcB/5lIhdzu0vIvss3hi9Uln94fgiCGFNHBxePtcIc2TwedMTz0Aaj554A
8Xh5nWJ3bmnBwReS4UJWL2/iaaiP+TWzt0nR4sUu8RUZwagj58nhrIKCnIq9m2NH
oq94lcZdMv/2kS8a9nX9V60dCr16UDa5UOr/zBRnN+ZQDfxvj2hr0vhUkYI4nzAq
NR4BWQ0nqiFZU7eNOUhFzALoIR1/q+7s+SNoqnsD1chA3bSD6O03kl1rq6xGm2Vd
mhrfV5cNEqKUCW5NGvyZqr+3WL0cW9ExMvUT7L+a6cAJ071GQWUGHNO2Adqvm3BS
THd+Xn1LMav2PwxGANKFCncXJyAYIkwUsLR0/sHD50QX1Yj/XeFocRzc7eMBODfm
2IzCmkIjDZj4tvBfBIg0QSObEZGBmJtDLFeMN68p3zJJMxi1MQTpUztezkJgCiTz
FlXsSAq6b81ctHjFJ9SdW07uoH1Q94jKUYgMg1UWUSMU9gVg92tP3qJT0lGQak7U
pGkjd8oZxxfvQqaeFjmQfXKZdHCwuANAnaR160U0+4nTj87THiByv89E5/q9DpJJ
Maquyb2wuGZMA/5DyyVNlbH/N2Vs7X7Hz4l6C1dhOzMAfE+BUCX6BU7fV7Y6VDwq
rfxcCQ10dAg/uqke7vDxzM0RjY3EXPwLuK2abrDxIvBwj2BVGjglT+d7vCMcV68l
XHcE0QYYCLca6lvps/DSzPCZjO6v0i/tPjTGW0APvxniI2OFtq7jd+kaDD99CytC
hGlHAKvTiJZ2KWZUhowXepcHoPBSOlwkbsUIiXolUPU/TmZEl/216XXi5bKEOIo2
iSp0espKvN+0Ob/0VjVlcxRq8cfxWqOCz8GGFFF4aDFUYqn1dhHgD7QOBZjXZbjp
4lEW1yHrtYOh8XnIz2UXWeUvfD0IljA8LsVgWk+vHxDvq8JCU0Dpbpp9rp+r2TnR
MIlK4VYW17j+nAr2o6gPpmdB8WA6sLtZ3ZUuiQvhpEm16pN0buB7VlcmbLuw+sMG
JO3DBwhDB/CNbnXvbKtgCJlXAXLaUTSCqLOyGxLqzImxHXoMBUpow8DfBLp/xGHV
BAokehozBRjeimty1mdKJocPI6OJYGEUFRMI7OGhkeJqvvLjtUGcQOGgpBHO04kj
qC2waiVuxVn42k3XUn5hJ8TW2nf4CRLKyCIsQN63u3NSk+alPTFtvPfojHKtEFFa
CSV5ns1NoPHBP5CcW3CvlWng8dgAOk09L9Uqjg71rGbDEyQ6Ly8CQ9iUMq1OWP/C
9eGtJlQ/36iOSsvpuMdUkP6Cx/ug9bzQf1L2ylOMNqnO0SjynLK1ZHFNOrSZxo+G
PAw5sbXjI+IgbHQGb4UrnJi1oHCE2WEYlSgm0Ku06OuvFE83cQ8dj2qn7kOn0Zox
VU6Nd9Jlg1JteL1k6VizIUANJB+P+RjWyl9RW0VesCQrvyUeJgNasg+jpayhxW2E
p1Ex4wIPSCVq2ZcwzXT5fXH9wbyC8+viC5cnDLdZRqS0VFQcedFAFpm26MW3aPnN
pJLHnEyGVKPAOLPk4Q3p6Dho1/hYchUq3cMSHXyuLBuLek3F3p3NtuFQ6mHw3g/M
W21EuafT5j6L9yPfKCn5sKbzTq9A5At296wmiMySk/ZYw4/oKu9OL31TGVmIyPBW
hwKKEDniGSPEiAvcLGzJcFUapnyswKOvY0uYaKi54DGstEbxDZrIUhW86VYkS80X
wDXyCLJdu4w3Cgo/35rBXMYk3dZzO6Z+cYQQMDDPXJkb+T9sja39JWW8v+IVdJp/
18ZMsrbWKyK0uNVkUaNRD2dtL4UgIpe39jPnq7lFIHNkUMSNsSaLQVkkkaTPnhKZ
TvZ3c9XdDbMLf51wEVKkEg59qRDm5BD4eBSf4diMhnoGvRkNwu7yqDyVaZCmiEbG
5zORmzK8vlbg4r7MHtkeXgRoXb5m5QQMolgZOjxVKtRtOqk4kPl7h6QQ7+JtkcOd
z5jAvWWggrqssPBXkYElzfl2NZmZHHbTxr9c/sFuqTuOHNtRuygFj5xwNPZwktpr
4H5b/+UPG2g1KJwqF8D12WFySU4AHkvFzE4CjbdfIKPvqq80TGJrIHeec+RWOMwA
TTan5FKn/BC9WqKmM3N4dB8o7mq3XiVraEDRJT/S4v/9+/kuD61UB7SALbZMyrTm
sllvMO/r4KXFcBm9pOeZpsZ9V6WDZ7rxoG5mGzv51vtEvxw1QgrrGEGO5evosed0
s3yZZNFdfWbV7dU8XH0ZfMbz3nrbMyDKk3Lx+0Bjj6mdgtnXNMxgtAelvxSAOD33
L8O4NYbnCs2NPnS79hSJLeSOF/6SH5IQzTjNlshf2j2f+cTl1TivHgSmxPBf8208
qoGc2+7G4KOeD9S/CojS0S+M9BDQBRuwc/CIRub+oAUrq4yEa80kBn2CEnZYZ+u3
j9y472s2p+MpHOeT7tdg3e/kXbi3aHn2SqfXLgTeKhJaulJN2PXoi0YQr2pq5Zwl
7oIonrNxeYiXQf+bQzqrog9ACrxlsDj7JbMpNMQXeLWkkVa3L6UeGynmVc7G4vxW
v96hODDbjWePYz8NSFzbm5jhvXSU6U/LYl8NSBLLTJMS1ZkICDlMcDikhDt3hU5g
7DUk1/FZ3w1zaHl8/rssCOUiJXiUCEpf4CnRot3e179NTZtomcSCbOjYibCIjEcN
Yuscm4saHQoXfCegpaBvVZ9A90o9xjN87T97+F0qSVOfAnqlyhY5BsFcxvNojkbZ
JIBaskC+wAxkUdw9hdTivL7oPUNyW8Tq0R8RLhulkxgqlPRuR/9OChg5yQ3zno+J
comzWDbmWscsrn4sP5Lm5UgK5KdSr7Qz/g/pSBE0d6+tRt9MmWsgHJAPY6hLGgxY
XKTysNSK33SHY+onxGB84U86yJB20x08lMo2ZcMvrsuEFNQq0Ee5txUIyPOInyJH
mLfdzD/34thwOftktC0fjPZagk4A5WGH6xKQUhaqU6siXmw4CojjNkgQeG47r7xf
rGRJidw1TWzlvzU/FR9k1NjES9HdB2pxSQWlWQpNyvYyNjZ23iv4Z4DwVN50b3jT
03zvvdNm+zF8CG+y7JcKAWWyDcW6Ew+QQOeSRnu2vxgBGo8Q405UW90yLwbJ47Ka
qcsW30qavh0m3qnk9/2cRPr1yxlvBAQqQwuhUKXcYcmiK4k0ddAXSwG28vIxFLkt
AmCDtRsrgHaNRHt0QyTWkmRA4Y8ScQ4ELxeDu0hZrdbD2/U+BXysX/bGXzKfRViM
P120FpjL1ti0EZW9DBgTWgo6fqrnpiXJVv9TVAw/ZXrbweeR5h8ivS5T722kiwr6
OnZCv/jGuRtPyTkEdM9Kp25+BezSQSQpI9hpoMf51NqV1U0xh4sPSdGpKFG3bbOq
7yhb3Sb4FzFRSx4sFP+15vrS6nKBlMO8kP+9QwIkFF/esvQteKc7mnNfn/jcvrxo
isF5JAUwAqtaOxiqqoI9FcXrtPUgsIhIsa2UwMwDfbQ2eQOWS9Lyu6hNO/cK6RJi
8YP9OLn7v1HgvQ08FH0giErw/IOIu+nOTJcgV10a2tgIDxMUp1hWhaldKrU0HO7/
G3A+zYYyHaaAS/5Wd4MdmDPpWE/vekIN4H4CI3Xx3uV4MFLz1k8UKHQ+wSQ+cIgR
xuEryJwB8UpexSgyjlnvcnQgOyxVVdlvD+8RUOB7SOkEFSt3pmSh9WdLv4J6xniP
MbDfH13TPxHYwzain88bHdRnlcJceqE+1fW+hpJlLNAcOz90SwrjtC+oTdi918ta
/MjkdT9YrIsNwRLpHIWXAN8d9v9bhY9n174ObUH/1df6W16NvDOssr41fGbFHqkK
J49ASMwyVOXOmVCzoUZltvK3oTk1i+TiaTftc8nmUToZH0Rfs7rtV5nlundLo2GF
EaC2hlYSCIocG1TZKcw+JXyHhGmL0vSuFbsku8tFyj0j9+Cqpaowja7Ht+yVFrrB
zc1sZUBEMg8bfbCjZaFENKLqD2a42ELFPkUP5lZmnWHDSz8OR5yyXPAm3FDTGlo6
P+K6hSum9R3DdXFA0G9PxUgWje3cR0XDevQHRxY+6mAp6MZQFgb/G2m2r0IELXAC
KC+wL8fmg+K8zIuUshVnsq5qewiAz89g2WppwMXfcoRwBZdiauUBFFQ7hzfMywoH
P3NkOPvNZ7s9Sf90Sc09wc5f1DfGJLl3WDJpUPVhu9a2bzqo8crD3ZN9IvZsKmnu
mJbSjtxTIVE0LzYCFk7ZMPP1qmS/Wx8KQi/ezawDMqdh7qV/Z/sid2AcZUKSitB0
F1Sj7PI1RWNM1khqtRYJDeA5psLQQKGAEo0lv3ydwKOBOB5uxMCGCDfqOExSSGG4
F36QKcvtdXMfKQAF0tUUl21RJ678zfWYfMKDG1hKzK4MkxJf1c3DDEJIti1rFK4e
VxVgAo8T2yQyQ+FrClq4s6R0Ac0/G+1eL49ZShvJ9wB/PfR86Far2p6tZfNZ5w9O
crxO4kImzxCQ0ZOCEFiPR37bAyAGDMxe8iGi1sUieDBX5WUjKDZ/qB7UbRnfy3+B
s2LEVCDOoWcg6tU/srv3SXns2dsggXEa1vgp2ffzpoHaS/tNENutFXHvZl0Eqw4o
hhtdYUy7e9yvHj5jTUkgKcIXDLecz8yuCAdc0V9KghXBTEqONEevD/Chy1PWqoaU
ZuSTzdNaPUr+heg1HeLcpeAQiO3fJ2Ey3yBMcaQYCqjQaY5V4pEdTiF2wMyIjJSj
DU3IJ4ce5WEl6V0E5v3Mo3igVxhYr1HZqN7VslBztTXyGbdEE5elMLluhonvS79h
c/uyAx+2bd1SlZTjmhgaUXenu/3BWTaRQQ2KNPWQV4VeuQsFu4oYqZRsGAOMZ5wL
kXhJDTIQwbRD8HjynlGyBs/V/Be4qSZZ5HcOw8+Q0m89EN0rZQpTilCbWkYoUF5u
6udu2gzbtKE6zX1X/LQzt2HN0WpKq76IfUNwRoFLs6U1brdUolJ0Yg7b32Zy4LaO
p23B/6tphgno3rXIHTri3HsVcXADTzWRwfcG7FmrulMfIZqplt9nQhAcGo1irzb3
1FxoGiocQEcPMlalBv+2NR8S80+064VPSz1mvw/xyObt2zfLnFnzA9JX5VugBDzX
ZDA9snOn2E+hpgTgH3iMlS9iNQ3CIwfxhEvFdqfPf+2x1IrWByl9jzXtyMco2PXh
qJZaWdVsQr/kmQrMKeeBSZ4vYRCFNnaxuHpdrvyLf5h+xfB0GNU+oQdYKO+cf0Oe
Y2ROm3w1/StvqWs7eTVYFVhxWvvg3W/FeqmQcxNjqD69p0vZq0f+bjK0KRmr7hM6
FuxFq4U2yzsVlveVyXPOQSN2VmGzUfpBV2EmHX2UT/+mV8TvfpCAtdMdg5TPv57y
TLLHZBHLza/8QmIKfPszW2l5gmWwYAbzwqW4ZHMG67g3RMJYIG9jD8a7GX1wg4wY
MlpOa8B3gg1jReToCkG0W3oyS2D571a+LDTegD60PPlfTrNiP9LUEEGcKWe9cIaP
Ta3lvh5NRdq+sxPnY2H1/zaKXBiVS0513QBE/3QZ4EjB3vj53kKnIelsABWLnyiC
`protect END_PROTECTED
