`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2+IUG8CpGVRXPejqK6OR3m50QKApGzQ1k7WrP7DDgzzKJzYCacBdqkrb2VfWbqg
KeKo+1IkF4WBJIBgDB4yQ84BzrQiveajC7psSLGC20wu/7iCCqvk8vD8TcGohvCq
3WEzC1FCByKJF7zvDzkXhmLW/eLW5Vd+FO5OyUUhNgDQhobPE5xqeZSYnB/2e+fa
KzYlx+1v9XVLgLVroe+yet5czYJ/QglTpBoEHaGkS9g6mVgQeGjzQNjh/V/VlMwp
DMRBGs7xCn7tvRToGltBiWCX/zXHgstxq+/intAWBol8a9dd738FXzlKxbEI3VJI
wH2P2qVTUOWfFjFbJr96bGs5oAakUnYMUqK/5jXEDeUr2WQ7LInRsRHRwA8qthXK
8Lnth9hW7C6K3L94D3bEoHfeKbY7l7JJatYhtpFcIejgV3f3quGsyR6PuHInGu/x
NIoqdVjXSvnXcZinS+m4ZnvMnnA4HzhotBvOSy7D1gp+uKfAcmFwTs341BKwEbPg
nnIru7VUvah+7p0wx9kLjYpV/VnsTBuxoCIEHjUYtWa9fWL4toAaZX8ujAhOTPWS
wwxDAwECCw2GpYOP2P8ZINzNtMyBZ3hgIfd9Y4i0UCYjHwYnp9jbcPDS4foaldiC
yL7D16w1EFZ4KgtBH/HZH7TY0CCWnXeCluZfJnRjjFY/Xv5O8vSOONifbImuhZXu
ZdQiivy5yF6OYP1k4fz4yMlMpTTE95aPtEdH3F/eNN779CkPp2Um63COKSzLKirH
tooA4M7aRmMhpsmr5qhB2t6cXbC2fVwKs9DotPNNkgN4Zaqb7xJYLXIs2t8Y7VxT
hZ3x1JSes7ujKsdAW7wPSpZF7uk6v3fMbN0KjSqkgB+QEBkjUnHfxMUsF3kK0/Cl
tESfytOCKj/YuSph/VooTfWF4jl1bJ7rOMx4ibMjCuovRzIDUY7MQegt35DUv1WC
tuulsqzlb56/Nxuj4oJB0qlEF0trgX9Z2qCSNpChKeEOdYDzBuIyM04EW3wyl8Yh
p6CSQ11+8ll+2zV9GQlaE8CsNgHiycgvuG4RfLPUPKng3GZSmDrS8y0Z+uDqe9qL
FakgZwqBKG/MC+Q2Gs0gzWHoEFZqVJ7Z0RXZcbsVjep+H0b7pDlUNsjjTnkRNQqI
0EAHf+c8Jy2zlebUa069uGw78CiYrED9lHqkY7xkGARgQjZjoW7KZtcwfXI9K13x
Gn/1TZA5axxItEWa3XE7lAtQa3Zhdyz3HtFVqfVu0DbiznCs82JdQtLOPl69JCTv
udcVPMJBfcrhjORkHgYWugDjDICMBTu/af4EvjfqdiIrXovoRtWr0siCdtyW/e8i
qgpy135A2i9NWw7hunSXUku8y6V14Ni+tni69QOhB8ndWDBceejAY5cm1S7TSono
R9hg47GiGopQjbaLTRQkJ/syB3YWjW8aaXPIEtFA6ylLSl/PrLgIOvHnBn1V8bwP
YH3msu6wPYwtMNgXnhQ7rFy7YrKnYBbiKX0WNks5CugMO4VfW92XsfxhxWJdaEUL
TqFT1MBFKyZ0W+bmImTx2wowNLtrro+qtTxoXE8/L770CfPPTEdPbJzquPENrh5C
pApxH/sa8aOGI3hafU08Pg5JkHIxLdOcceYS6H3DS3JTFTL/ipTVH4ykFtclFqqU
4mHl+ZTQXH5n+LIZVWpmTmZ7rMmXeiCK2UzvdjwWW9/bKZpuKPVOWXRxPj+KudjK
pPGb/Mran9FMZHEESJPukexaPz/CRqh6d+puy1VGOmWvl8YI4ISMmk61PN57im33
W3ELiEqYnitYbTdVJ7NNS+gRhCNsO9CCopBISrShrCZqb4/CPakXfLIM+ban2Xgv
AZ2VlmmreVVp5xnLaI1rO6JYhKdc6PheQbl3XZpRtgBjT2lVmDGzekLm+QOLKZ2Y
+2ckOVU0h6x50R0OfU4j5ODKyhTPl/zs32coX1j+VPzYMr8fhs+oc10NAEAmbrIQ
lEUm/41J46hU/m/Gz2tl5ks81y+s56CQZy3X2/PIcTVPWNQPOjaHK8fZQFF18dev
q6FTugBe85a6bCkRN+e2wUupJ+GLopK6kxmSerPzpr1KBDYRJ3I4pJuj3krZzJxk
zHcpCvQT5TR2mnLkdYRdbXnBb6unM/u+Ro0KOX72873IKG+TunabQdalHPduOJbM
yMwU2RraduG3HQNqRfyCc5mOhOjcPGqLYifYhII78HcKK81edKQJd6MBIvdOquFp
sGDhhTCdhEfd4XbXa7TZlQxlXco8w/jG6oYtzRX3CuiBYp6ss2ePLeh6I3k971HJ
5qXtzLb3F/s8i+n8yfdJc3Ji809WM2x2UBIktBduqcw9EJYSi+G+BcrILYEwpazt
JoLZA+HbxVJ6EknsgM8wEBMKtiOWqy1KhAg1VO0p40w4hRZ64fGjNgwOeXKo4nYj
H6HojVrtSWQzwhznxWDJnrHjmVV11rSjxZAzdopEhPKKAaNiST4yv1OgbEE9IeM1
DH6HajoaX2jY8pfmTRKtYtrNaxV94tnJOs5qGUbdqSHR4AK78qDTi8Z/eATGKwDJ
Q2WSQRwp4a+0XFdLUzDplN9q3V1t59vCkRmzXUT6afaL1klK8ZDyYWiktk/1NIWZ
FNoCj8mn8Q57d+bE3T4NOs7CeD2uPoaevUH/LbZrQmpVIgs/pZhhPoHvS7bMNkYn
BjOvUwCes1ABoi/Jm5P0x0mXPkPdnEbrlY4gbwjj1NsSZCxxRXpGo51DV/AD1t4H
10n/0pPyuMmYJ81jwH80Q0CIDr4LGrgEjxeulL5TthLx7Eq052O8JNLTRXR4WPLk
Xbf6EvbdqNv8cO51xS1OfdW16yuRcfqPZpEiut+prub0U5UhM+YZhnM7DN+SyTcg
Rqt2pRAUaMLTdivXmsjwK0Qs+4M6zovOQJpDwgQzevjLJAsOjZZaL1tX8gF46z67
qQMETuNS9j6kvfb2Fp7q9MwCCMyNfBOThCm+8FDPmv0DPTiMy0LjFgkGBTMcdny7
qplSiE23JfUGF+6FW48c2jSqTFoB4KtsO/pvFB6w/UDLXNezmaEb5zSaWeIAX2e/
Sm693p1UhRVMvaPuA0Ivo3uyGbfIFK7CPJmDpz7vo8k3oJ297ePU+fTM921JJ0pv
X5L51M8xRPSE3EOGw65I8EuFC3Tgwht7OCiom8eiaW+4GWfLW1y03CUreaYjSfyX
mqhu+Vf0bM6WS8jZ6PJEg6xQ1xskrmoCj84XU6UZRmoilsTC09t6pKRsFBglIMaY
FQjDp0o7/zOSBQcDNyx6aeV4qmFZqBjQy7Xiy3QF1Co22nOEp+F8yGPZOmIkSzX8
6fdRiI+ugvJzZaRlZZP2Fm+K0eKsWE6U9j4hmVTEKyz3IwyMm7xVFRyd5aaV9uGO
TZPJTRlImtzaEbI6EpQ42rh66HWk66JPwjTr1JGidtfqAwQEQ34ErYWW0564kiFm
BPWPHbVrEdMSo7tS3hSW8qZVVpqdFKNt8vK65/X4tA+tuFlmLEAK0TLj5dPlozre
MG2IcRQvDWu1QH5ETGEyKGI3OCw4M+HzO59GwyU9TGQemTTyeDXwIN5uFOn3fAS/
FAw6BlWQlySzPxPHgEsXYLmJnbyaPG042Yeqys1DTuBY+ihUH3EZvd1runFmS7Nm
4T/GiycTCAjfd1pokJJKm2ZSh2ft81tau1vBp9dL8GILp0o5by5R/zm0rtTwQC6+
vdhJfA4uzDIPPro0GcIbUw==
`protect END_PROTECTED
