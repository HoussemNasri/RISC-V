`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XQrg+QwUMXatlFz7D4J/GiOOyN/T0KpRorz1NfOl5yus3CL0ItoP3zWz1zuOIz2k
Mw4busjVEe3VORyo5XEP77ZkxBqqTyYs6LQ9oDfVG5rCiOIwev+4BXRgBflaKJoH
tLwYMi4GOqvkyWBCHZxi1MZF43uDUpK2T2vme2/jnYz9ML6dSZEqG8fXMC3GGn9R
nbv2UZkvpdOvGG3KF9yuXm0Ns+1lJkjBVJT0B5/Frgv6WsOLyTA4EHZ8YF5xOunh
F/e20ZZHGJFfKmKXlNm7kodk3aV5nRSYQFQWqI9Vr2ktZ2ESuB2te0PlWEHP/JX5
puxTxMuKx6tviPEa7+NjNQeCPawWtS6xXy9dnSjSIluzBWUH2jJhTxTxHyTY9yFs
okIRG0+5WkTpElsFOB5RpgOf5xldk8yo5IR7RyZLwMGmOZrTnIZnZgLWNb4rgl2R
+z2j0C6e2Co8XHlJfLC2feomE4rxKIovwZtM5ue/cqwokhq0eSNobEP67m50zayW
JMu6wauHDAcuujDynBmuN7T+pWzim/0D2ZgWv3YRROzab2AxHH4gh40w5fVi+ul8
hWeEO2Oc7USBJgbAzLNc4MeH3aV+5Vf4x+XflGkOsspOHVoy9q2h6ork+rDqhuRw
sVnr+CC7mbGEye+8cQ7Nrw/imVg4J9JbaRTgL3VSUzOcWLJuzufMrJQmcYKsK+Jr
Xzgkv+UAbAqg8q4Anu1mWKwHTAJtPBsfMM39VoqAezTpxQA+E9jNsoXsvPw0gRgR
EdepD9G4WwFHVb+ejRG6nT/wUPaQHXtJPmUyHW3BZ2J+oBWDZxJ/wprr/syueROw
8gk6NiMzL1qnxmJrq7q2WuWrDhq2dp46eO2WNxE7I9FSPnBqi1PbyA59vQEk7pG4
sjwJItmPUsKEbRQnjxbBojhhQHR35Hbx9gdquuOF0XT8fuigj53K9lCSlOwYYM2m
2nGlQr14i/yurTXdT4l9DlIraMa3uJ9wo9rz793nVf09h10uc9CYVSEGonpA1CZf
dg/5BWyApI06vPj7nmK89hnkv9NVxxORGDy/9h+JHfGUh97FPKhHF8efOylAF994
ymvGfrLE8NEi9eQPogMSuxkpeEY7O722wcpSIVBL4B0QDk2vTscKd0GyrpQ90V58
3msCvbcOXRt872vQ+Hb5SXlWlGsdbuM55nkx53OBV1yfY3AqN+Hjeq1S+EBganLd
KOJIRFdqvHNJrrJRNEtI1usryczRM3ajmPfwyUAU1gMv8tKeVtwnA1GnfynBuens
yIAW9W0c8gPT2D8qrsbW7JerCbl6s1o8GL13ZA2FKcXBxWEBw0SdtLuiDTz/3RGE
rkGhMQRjedD1wK49Mh3bsQxC61VowfX9PPGj3T9I7vAEvpIDlHIRu3UCdY7RzZW2
jtSUTo6JxMd5o23+hO1ngp6+49RqupNgPQYXYooPODDIB57OQydun8hnsU0/AilH
OMdu+Zh2J4FHBqeBwP6XU3s2bESrVo6VvF/5xpOFFXVVBEFQFIzuRvJYwTPfy+iU
anZQBW7Xi5QGz1VYEL2/Zw0dwKx2oUPHQqPEA1OolEa3ljtJjmwUKEDGFJonJW+T
2VInqaPDy+yDZe371Iz6y2XxjOKc8eCm/KhEfVXdORk=
`protect END_PROTECTED
