`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDYlUGHXHZWMPHmSlyHt5ZbrcVh3OFrapZ/aqhqndN52UD11Ug0c0RpoUdvQqBEc
aqNp4Y8d6EtL2GyPqLr8FJOf1fObAydI1YCTr1f2+eCKbtkhWereD2G+6Klju1kD
TYuoC6+3cPicRKCp4RevZ9J8YGc5iKaY8UYGFPKi0ZJPjX/6Cvp869lMWU0LtJEx
iBVYgi82OIkgELqMZtYyIj7Lj9VTPgPnmW51KOJb6yzirGe8VStZOsez/h20jn1C
N0RzeGQFFX4/C+Sg9Yq9HIxVtCCW7f+HAh//5YZMU6XzKZtwNJC+uX3WUU36hCpj
mh7jDx5pCGNX/Sm1izgccu2Kqx1Xz7HZcoKlqOxggY6Pyb1MukjBUzl1XpiR7Wdi
FybwssfgyNFseXcicZVGo9+X0y/vliDpxN0bcAb5klrPBHP93oMYba3gweUB/V17
KmKYfCJQlIDMThe16GFejdxSpDZ5FOmuKYSG2Q42XbWFSLJMbg8ODeDxmViNjO8o
wuKfe9elb/6qN1D56oN8zXLkvaMOcFSacurcMtdW1JRc3sAqkmeI6aiASzoAYIHc
n+aWmDs5Y6cIf6Vkx06Dh8dBMf4bEUF4CZiXdxEg1zGhbw3/bb93nEG9tZT/Obcx
8bkMvxqSeuP15BlmfsYdAEQxbenQQOYXFW0euP+fm0ZxBhdH7jWQouzbxgnSo9bI
YreDU85eU0t1qeFLFYUQXYFfa0UR9FhEubshmmhno4cjkNJuGo5Hwy3QJwvV/eNd
RDKfp7QX3TQyP4XfBdZGSCnSx+4MuVxR6NV0P+Nn4aiiAiVZgOJtxhHwN1pkrDZT
6xUQuB7tVcUrDHT/qBUAg7joWdrAlVtw2tOwDDpzUVCsduswkk8QncoAeZlAHdtQ
Dewum/ZXylwNcmTg/5W03dztrT2Zs8CDNhPflJchGwn+h/a1RbTFsLdFs7HT+elW
ROg0k7PGkfrLUhmFgRK6imaovq+y7yw69MPfpFcmSTUB0K8ZzEpOlUJv2lt3m2gC
rv5JnNHBv0/Dpd0TW9U8kmIGetEkUxE1GhAcGBMbHmuKnmmKjoyDXXmkEHoxUEa5
29iUcv/FYnqp1YTJa7wOxczeDD5PjJhbic+TI1Nv92lRWGu2XGpqGzCP9RJVMxcZ
Adrr+C90h2F5JL06L+dK7w2+e9g4T2Aaxv864qOmUPNzOzmANCkkSEXDxnDr0tNy
YsArjMTar4eDpcqFsBc6u/5CYZR90NQp+TLWo6V7GRv7n4Rbr9flE18+UaclwToS
ReE6DpGOl0GcxygbL+nbYaGAfwsP9zvTWkt0WdhZLdpkC+Noqn/Zq7gHGO6H0GR/
zKddZRODEMEVWpDghwEeD7fjfqHPto+hreZriH7M2U7b9RX1H+aXuQkPjzjiJ4Y1
hdhMtrfUgyaC4V1H19VWeaBh1k1UMc1e1kvhQdIeHnGqIOTqlVCuVxHno9Otx4tm
zaGNFpWr7yNKAwgTpk127IpO9d/cNcCTtFyTLsseC21e7rcKzhQwrS3u5WCPQKaf
wPZC2QX3qwh9G3xvSirAEYLXwH3Zkb1bh3GrGa5HsTUDLB/uOoIZE8+I9LXP/ay+
RwUTsKZrr1ZoDjCN8FWSiQDD5wp0KSpF+gvVky7mDrE//obDceviar8dAlApQVJv
OC8WWY5FgVqKoyK8kHYGdakGdGW8ChTDUzdxcVMLvPNBSWnhcrHVnKF7YciyI3Dt
OXTX261PcPYiclWpr1xEenwpWPjctTb0nceF/M6zH0qdOj0+Md2rUG4ygJFqddnv
EFwAsLjEvd9xXAwFtu/ETllwejzyqrG0hwQRRTnJsKNlP3tjyLlqEkAm7gEnIQoB
901EsoXPavhs2GpxaKF0qK8cQcHhlYYHK92Vz9EtsLoRRnSaogkX7WC2YtVccApZ
pVEqAXTsj/ALBhC0gThhOZnrcftcL4Fo2nLNecBtgj8etZgYJN388fau7sA6OnXu
ey4HlpWybigr7MwRyVhjH9PJVzA5TxS0f60qxSA0vvFyV/BcLqOpr+sjSoFv6bB1
RR/dgxntHmv2BnpfZeAb6Zg4siLzHGguLLBIruG1x78viDZ0HKE1AByGMJwR4l6G
ka8XsJHK1NYOLnsNnAhUVOYUNuhOtWjqtJTjdwHtJSOpzoFQOO7OZqOCOergTWJG
BntSHJTrVyfRP0s6SdAsW7NIZrmPa+bSRMBHI7N65xCwfPklpgq6h5ouoohL8MaG
81CJgjXupszhAVyHQIrBUtS/lU82fHTDY10E9HZLtc91TOhZBT0jVlWRDjWWrwhA
5bDjZwO5iuGmJVa4QLj+04PoxiyhY9+wUiQRQL0YEx0ZQSwRFwYeBm0qgCNm9XWS
zrf5Jdsb3mbMquDij2yAesbOD8RFEx/lpj/XWEhFijxcD76/nFPqD8E6u4D/Z8M4
hjJy/Hx+7RZFSHMCPLdCY78bWycU1yfisBmGgETeEtO/8LgWMqKLmFHv7rCJfTSX
DzQFbwxzhKheICANGZV+0HjlIuAhYrYghWZiryuMIvoRByy+7k21TNkKtQ31Ww9V
QhhhKHw5QO1+00o0yBFnlpKTdXDUsYMGV+xElUPuiejsd0S5MD3ajWJBFsJbz47S
2SDDvEnpDkUGPBe4uFLmqdSajJv8WnhEY5f+vZCVs53BT4sq2m0LOCJkz7ffiNZa
4j5V4xvL9y9eGMw5PdAynuAw6ZRjKUVGxrznrDptishez2hLz0v7tFp3U2QgMiZf
5YS4sribeP2ZiSlSc2YQeJALPh1imoQ/qUlE++XK0DQHBNxXTLO0ovESm2KT+oG8
25lVN0GHJAaoLUaCz00lMiXxEZAuHm4P+o8Mj+N8XTuJw5FuASS6xtmQIiSDAZWN
E7Qz4BkoeMvfiqtJwpsXNTDFwdw7EYbOhvize0Oq+9kpGrqJNsqXqKXiNs9YZQrc
uUX8C+m8TuejJVcWiPDBIc7L8trPUx409XlhruR+XfQhvzmmbxCO6UgpuBDs8dvK
TTHQb7/iccJGcoitHRD8q2HJeVo1WUcvlgZq7Fbio2YSzrWBpezJ1UvN83dojSpl
Q1ZB1Kx+s+V2ncKRUMdgB6e/jCdsPsWEc58sFR0w4DEiy3+CB3izfJQo0cHAr4Xb
NjASyGUtGP6ZHNfPDACb4TgJy2bHytPXHjK9OXG6tdcWwZLz2YBeQBgeMJoZCkoq
OT3uXFM4f7uF/yLyVj303mCZ0Jhmx/SloJ+26Baws05HvtosGCju2oipfbVAWcvR
/3UYKUljxsP5rKPmxgRRjEhrS+nKYMRasyB0YNNOIhn6gNWMwYsMB00CmL0MLstM
5T6d36CIDop0QWu3K13fM3iitlXa57onM5yPgQt9SsJZ+KT5au9Nk+vBFlOZY3fc
ZDVgHJyNGkwUe+bzY6wYLdbJvQN/e7z7rVWMS/U42FcC8T2eiCtL6hZcTBmLtJpy
OPVCaq8TgChuWlb3kyjWQO0XXKRmKUq/1k6JNgw88/qY9UMC9o3jN/ynv+PaCglB
Tt1zOKb6oC/e9JEXIyu8nnY266I52NdKugJiN6DYb+PK5IlG7SZ8S8bG0fr6IiwZ
SoSfIMDokf90emoGeTRJ1IXQnCM/bFphqYyG9WpWHov6I0MkrYsqbgdhWBA3Nn1k
/Fa11lteRDVF9Ny0YGiowTdSurNxgJdz/918nS4ddQAXpXYZKUpM4X41vMN8kPVy
228EhrlQziDuPnFBXljhNiBYgjMKh78AVIiGb15p9CKl7xgsmORVwxtZC7NnDFPN
adr5eLg+qVNFX7S4YO2C34lgQOv65ERJ0rcYxEdvu6w9G2J6K701PGkFDUtsYgA4
ola2u/OQHIxqEDxDDBB1CZ8eTDRx4wiw3+oWbhD7rzuE8sLl3/VcBR58xxEGlJ7j
LQ5MrUBmcFPlvAR4mfSL7xVg8tFBXCJOstU1rcKpmlSv/1kyFeZhsGhE3Q5c6Gyx
KmtMdFwM81ZemdRMj8DzwVyT7cfsSd4BBkg4eVkamDxDqUZPbfEvNBRmP7tAtEDi
241Vy8FEoMfX8y2hPOYyEj4gPYH322JOEXhfJa1ZAlzc17tM8GEocZM0Jm+9MVxi
zoBbEZEy1sC+OsAPpWRc36t+hTD7Qiy6YqIGgwENNCsBL+k8Bv9pwrrYNHtpHafB
VQdp4xUAiV7jAELagdOcpPw7Q7FlRoi+Q8HXqneQS5DdeFSBMCb5Vq0R2ZUCsZQ2
k3Dii8/9bRfL7Z0lFCzBHmvrVDAtOgA/xF2EXZQK9bYS5DSJQ4I+PoIU1YipDUeQ
2eaoX2JKCOVoTkaDMD2lKmvl1s1p6wIrcAdilMbnl3KaJRZWb5Q2RMUjJtR4vZ47
lwraYq6zMvx6Y0ttgcynZb89Rgl9WBQ1nBHPmG5AQA/vCOmbEmZvlJTGHvTDHWMm
TkvRVn281CN99gK416oz0FM9oIC/X1w90C60cr2GwKWWYMaMrcCjm/588EIW38sz
fEbJD0lYl0Kb1F4sJF36/biS2/6wldrIT0x3hWMr0/0LsdNVn8ItUqiQqPaxyzWZ
i5RmdeZAE2v1/3la2xenLcbqbvjb1y2f0QFXJGLOTIqATujoQ6UUnxJRY6wN7uCL
ldL4KGiC9JSRmQmCVEQJ6TH5mUJmKfp3tPnQuaODCOOmVv6FY5a5AYJ9iE+lQ5uL
AnyYCZ/FncwX2Uj1tpQ1kbvMx1GdEE9hcejR9LMJyvH16axQdiFsLXQHVtgPgYwp
qwfxAA06D5UQ+bIlhJHyizqoM1io4yCCqWOsBqfHierkpFaPKYYW5J4q8/85xtR9
8HrnqeutRHZWSNJE6h3xN4XmQ/U/45m+LBhQK0605vj2UQd0neaLdLMxCf5C+WT4
TXvzb4hiSNAgvonZjkdePyyjubX8Wn/VOYQWaEQLI/7jN6dEpksF2Jsnc21tFGvv
8RCIXPA41tcuf81Ai7S58Cr1YTVEsO0FuCo4Am8frVNLxaxcBv43fxHlY43Bsz5B
iI3w2thR/RHks13K4fcqJS7v8HreaX5BoVgnWBDPurQacpY9VsO5SGH/X1srCvlK
buP+oMAZyNcOKiUyXpcg4YSQ89vgty5KBVlbr1xhEI7ALdXZm/3pbmQZWnt78IBx
3gspZcnAiNr5BFHSOireytUMK8ParGsSU/+MYmlkQY2+oGtHbNsKlC//+r1Hs5H6
4AqaJ485h0+9zHmPJNyQKZPrA8xzhxjbHnO3BjG1e1cJdKIaRMeZaj9j4+9q1NpZ
hbfcb5Rs57qxaabVRYvFMB7PGE8ZPAuNOy6sD8XIINN2cuuUvcPtiQzu8/qwkKFs
5vxjP/5/hFvowhu3u/tgcdb5Inaw1lJytyPXGANg5qYypsJjR/AZwgH8ObXR7j1G
mA7b8EKYlGn/k8GpvkjeFAFOaGTAHONY4aOgeEKM0SBJVY/58CYw9E7vf9ggXSbG
ArKbgHvuZtaDdfVTtPuw+Yken0+Wo10JY5j7LWheHWkRAF/BhKmjgY1OSC6Ypber
dYKN2mYclxHKKKee4ySZuB1D61RGoMpfHgoCSHPNfkSM+Va03RZxfzNNux038mfv
2svA+6qiMin9ljc498yw+2vAkNUxgSrXeCRYA3kirG/wTJOWG+mW+gL/I7spI1CN
8o2/wktEQzoan53HYBiKzoT6qonN+Yq7KDmGdeDMstU9J4k52oSPK/ziFjK0FJVw
Mww7LY6Md9kNrBcGPYKJSpJQOI1rX/Irmh79xswcVZK4H2RUTQzHyjg0wrWV4aDA
xmrUYji6VqNzeG9KH1aPBjqYTKanEHWlSRFdxPX2n1KwocVhAFlPG+69t4zVjxzK
4OugDVVBbcHUaz70JFcDlznwspbylmybhLnjA/asMruDqQpTyyFcdVyY0b5YqYfF
3f6DKGVaMr9NUXrX7FcpA4uj0dAIdPq9dYEr6G0ACKY6epkGpzEV/LWU6F1UVXme
BnHFDBolZgnos8L6Y7Bk7q0g4r4HMLwHLShPrHi/DubSl+LqnuIb8gSa03l7tJXe
ToYzUPJDKDKEYx9FS4jo0Dc/zH9QjZYjFmd14ZthesLIRDUToIyFTc/O30KmKqow
5KH3XMjfP3V0CYMIONw3zCafCPq/9DFxScfChAkeYO4z6GjNQ6WXgY2jZyVstDws
LKRNF/YBFWNb2fa4Enrv3gG14g4PiU6wRThGiglBx/Aeo7qXWJTQi3lcMS9dibcj
LjnESU6ekI4cKrSumU+NuJfuI0I/BcwmVisp34jzYceqKvK43L9KJNfrORoZR6gT
kJ/2iebGAWm8JNJq7UOj4JJt80nrG4xLpoOCqeeoqjADHXCBsqDY4DBULSr9OWID
xjUfElu1NfQkqvbcignMdsLHz5P6mdzdBy3reBwamSMZJ8ekQxRNY5W1lUon1Gtp
Mctn+4qD2Fx3F0xp1CqdlUemuWlBQRqhr3qrbKJnzeaE56N5GdmuFBYqovWimOO6
FGvajWVYfMn8NbnmMu8P6ji8OZn9y+5PwXKX5HLCB0S7qsZS0nIEsM7P20M3+cht
1Q2U6fx9BrbQRw7ANUZyrResPfZzADLeaTwAh1UY0PGmorSKdMUpu6jgAXsLm3tB
y5GeXxUufIGCXmRi/pd+gW8ak/OAC38qbyHCnk2rFKX7jNulGahKGbExrk/6ICra
Ea8RYYWTyuZQceoFamV6N342ajj2U8wBbGnOvh0GGOU6xPtL7u/xtGnt+Wc92ZA5
0MjXUXYFhjwyh3ybBl1BDY7SfSnKeqBHgo68blWvElZ0y41Q3SRsF9q8/QWV80+x
C+oPZDJmrj7i6Eo4+uXdNaMx3PHiioEh5SJ4WmJpo7GoJ+2k0cTPBWQiMVxvOQVw
0zEC2x/M/R+qvR5carg2qX5LuUxCdno+NU4cHo5ZGZeesqBMYYxcZz8FASFMjEc8
xccSEErnLcnCzpmxMw8FYizM7XjeyvHNbaUGzae/vMTu6kr+BuLqUFliCvjtAwZV
z2rfmzFwW62lP9I2lredWRVCb+JefUCe799LLBP/ONcF/v76/DSPD+4rmKyznz/Z
Xwa35P+RDxN+eXy2Oik30K1S38pj6tjHRAoUajzlSM24+IvHrDVdgWWmvzweEy4/
uGQ+Lqr9ETpyhZv97CtBntbYLhJN3L19ZbaR1+U+pHLKwEiiSNWhvHMxex/ut7WW
+UzYzwxc86/xiisS5jyj8PQgeN7MYqfz4GIi/8taKQqS+6rUQ1HskT9B8c03U2xa
xF1GTZVEXZHIw6uJ63KJle9crMyCE6fDvVOnJ/MgHlUeoRj3PYsJBBlijJfURTry
Q/6MMwzoK4hbJjrBN0S0mA==
`protect END_PROTECTED
