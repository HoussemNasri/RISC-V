`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J1pXtmFT+eiENzwhKL+jOtTdOXEvjjxvaLehMyiVaNBJ/46k98/i/qfmlkkxsyJ/
HI1nSzaLV7P2gr7bBrwbMy0PlO3/ZHUAqhcNnWRKTkZibFrWonDpMvkhBYO1kgrx
ZTkRbuSByDXkj1A+U0o4uV3GYHKqkyQ+sUXdDr7U5naWk5jL2n+5jgqAgr/qHVHn
7nHes9tCZNicsBowQ4fkAiU9mcDA6DbP93Cxu31/Ebgu5J0V0lcEhAxrwZVYXYGm
cN73WiDKzQ0+Wl9DKd2n733cGV8+php2IDXA2N8kNwnWjrtdkotQnzui45PvVwVU
P20TMkrRyLk1HmFrfuuN62KHSQsfO98F6BMU7hSMC+wphe4mQ1N6fLYSq2k/N3J8
Ndb9+TdE9ss4s8Q5pH0llQ==
`protect END_PROTECTED
