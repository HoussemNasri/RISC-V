`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8OgFkA/XDzgmnj2/a8bbLfrTBpsho06crFg0yjCwASHfaRZCYYDEDVsPn1g2fjFM
zLnLhgAZGL1IEDXXhYXh63azV3Ol2EU9cpcwx8OXdjJtiiIB9ggqaRjfttDQfffx
ZQ/byHQcE3fTTs5ELKXWyEOhi2x/7zLLgDMPzDsYgiKqNlZLVmUiFmvlQCGwetzj
/WzQih9+GV89TZ/RHvDad2G4ZAyHVYeUDPiC4Pwz6sNSp6zEXPXzZtA91ZdayxXR
XWF1/VG5SKVpJNOSTq0OkOQIVtxnSC/pWV7ThP1zTZknW2r0Dky3pAqfUryEdShx
a5cjcQoG0mPx5LzqjPmoKk/iG5snWugFbYHm6kU5GGcienwqDj1/cCOpu/45B0Aq
CzE5oRYroFZwx0OVvLn20UAm+pRFukli4uGXYsb+ZJk9TeChsjmK2UEp8y+FQgRw
KdyPNeQttXxSHIGn8WuL3zOUwsdlJwMlezpG2/oguRyxRMti8EfyU3RhiAXFBIkY
NmEIedEA4MvXGdwJiZOk/xfPNtGR12l3z5t+vRy40LEX7FZAY6XGUcFmWUrNjfFr
AT17bYxVphySFmLHXhmbzoKS4tMT9fyeQWl6TJjkX9zULzfktYJD7EO4i/L883LJ
3JB8OilJnCpRkHR2uIW6fPo+WAW2fuVBrBTDivWofWo81vYpUf6G31oiM+QhhC3n
83A2hIyoyEsbT41bnslQrNVrsim1vcrVkCU9Bs+LHXvvxEG0yaYzO8lMdITS1kQp
24Pc8ExgmJiWOlqHXiw42T3zUUZD1SSqLYWcmGPing2lFPys3ptceoa+a3/avpXR
Uvy8tDlKaG7VQ73n/d1FoTCtUYOPygC1IJ4vRoTJO2TnGmdbKBtUO0znNUxdwpS7
+RoKw8wN7JLZeE9RAcRckXgc34pTYWQtkHNbP4XxmQ6bIhKSg2Fl72ZONv+be7j0
NodYU0fUPmUl5LkfY17PD3dPun3Qz7twYVeKvqso+ke+mo0bQ2HdCkIMPyXp+xwt
rKBgkLZDJe7kCB6WkyqXs4cwZCyUmh0adouFbQmfY3SrtkjQskUh/kZSfD+jmIJV
zvt+anen0ahL2Ma4uOuLOfufVyGR0x4+h+dWCrWGnc1VRY6g798sqYxZVrUrvdMd
Iz4jg12r8+HAjNmtYtw+NCOz+2BCo58PklPgv/ucx9h3xlTPBb4Rtvd5kzmYpaWa
3qoLudybxRCfy2/Catx1UGHYHguP5SeXAUfvlxnzip62qmUPB8/3ELT/SeJ1888k
M5GmGMALG0Feb2i0bPCG3cmhec9xa7lJqDP/pInnnJEApJB50WXJqFwOWp0n+7MI
00og3pg9Z5fJKxPaoXL32lVza46lmWyva2oE1RNHUUFm6epT2gFv7uG5gf9mWnBn
zXD+TnOIBUrqtH10yuO+VKP0VtjUWRfR6MY3UxsG6rzSfWQ2CYFUaqGRCqX5gYQn
HWhlqnxcHUSjHxI6pD/dktnipTaUqf2BfdoQa32EqhwwqJ1XgzUCsxYvYbC1K2bH
9xaXkOaoEywHz8kKLV6Q2lbMSAYGnrE1T6iCDce0D3CTEeBD9NF1rhWH2pfN0IUU
MV0ZPQPtJubLuxXse3i6KIQI9vyOzvtyGpBJMTh/w3GJasWlziklkMkKqUk075ep
AOB0QwY59uKiwVZI8uhoyvuL4K8JVH2Ps1+RP79i5mn++5rSXjacybSPHMBLycgu
QnjWiL3cic4ewvusMia3bMyTScDs00jvaCOCn2u4vpz9ij9xgY5LrbXeEPNk1eBs
FW8raYmBNdG0ftzHZ/rdAcirMALsT9x47eqzVjsVEnahookuvWj1+udxCSu3oqK1
3aGqFdyQvjGq17xRAVhmOdeN1w9qi6SVjdRWmqjoGc06TcYKxnprVX9+dtYaujSf
9Vw3fsmcZJO7y2YfpdGvIJOhF+3PBw6zYS8zGSc4rmJTrrKIc7BVdaPudjn2T21S
/XLvU1QWKof6UH2bIonYabQhBvj1zwb2oGnpYG1KWKKaYI9FEvNnCVRZVsHBSbhf
Empi22c9OFjHuczex0X//ACA6mo9evQ+VO2RM58JzZRxA1p9R1IFdnzzlSqBNyZB
Aqb5tHEJmSdx9XU+eUaPg+ChPzEigykg8Gsed+WOihTW2T/FrfR2h2UpsFzOA+7A
sWnSr3A4HtIUErqF6tzMGXor516zPw7cjVWpSeASKc9+8hP2ct6IDEHlNXLusb6Q
GhrOcz6CwkCw3vCs/OqQhWYUcnO8bSlZOU5FouRJIADOPlkg2RoKtVzQ7FXnwdT9
BB4KeH06HneCh0avGDr2QLVZLieL3aQoLNj+Fu5uFG+pwcrglkopiBSMgd/VZq9A
m44PZBjkbB/3CFQep+PJlVvtrgoQK0IlMti6b2ZRiU65X5o5iIr+mWaqt+twet7H
Qj5PhOy9w7+D5VqY8PHoN+u27mPzQRN7wqZL+/xfRo/X05x6FIw5w0LAODPLxIdO
ADwiF/m5ygA9PC5dajBVJ/orbp8GWFi7247Un2UDyFNz0QpfXDbIS1bTpZxC2S3G
xwAv00dm7sAR8WnhQYS+4FvDMVDmIiU8PwxMF/LuO2y3DuQSd/OrwX+53Nvp3zyE
z1NRWuMTee0IT3IjKIYEROGZp4WolJ404fgMmLDamRhmn8iOO4osKMcFeTcaVu8A
1BxV4aFelex/Tl6om4Xk79xgS5uqLfaVFCti4KBXFLIwcZgyFecPvFFgWVJouoR1
C9u1qwBH0Ct4rSDfqSXUes+3AIA2Ml7rL8zsaKIkkOvrwz8z9dfE+XfGzIwjFce5
kXDqAYOPR4kdlC4bDplNZnyKmLi6vCtF5XA8gFMeesG212PcaY/d6OpkUJ+751ER
T+D4L8pdZCzmHPhGPBUT6C0SCWOcxhKbN1OAMoPZnr4oAba9mhKLXHNKt/1IXeAV
dfphGFjtFldpfcRlt+VwQBQkVYK853FnjmDynflvPyB4v1OKFFeZpQZNOxdeMsIO
VasQnBv3JIvMCu0cklFEUnTUn9UM0QXRKIXqMgVVr/ZCUYE/HR5E5ptR4j0pomV+
bANBJpbB59faSEwOcJs0OdAT/jchKfD7huHFCscWBGVh6cxAirPS0X6S3PhDE9Bo
aVq0MbMoFCj6cAv/stTX98hB5jVmBWm9NIRGtZbPyU5g/47PGb/ZW0zqs6/rjJDX
z82NHIocbcd9l413NotcTlJwKJbwZ64yuDy/NGOsLjHxKROgvd5+xU6c8mWIDgHk
WuuZzytzVe8ZNyW+KhuhtcIFsZXrPweSjbhfg6IJqZkhnkuSvSqQ7tgnvDK5W3U1
u9gf7lrggYNK7mvwG9OKxm4A7zluucGlmm9DXTmrgBo6J2ba/NyIkn6I4RXa15Nl
qTpOINTcK2RrAu2AWLpeK7CUvpv+nRrytmF3zyjenFs5R7+qedGg8lbDPioJaKCN
w6vpMXbdVYUPyD2nifDOqVWqemYr76FrTewD/k4iwEqMQBctxljM54CP1pgwvDRZ
xtaGe8BUdS3Px0H4kvWCUFUCYlyzrHz9T3aGHuXuvp/74lj7+i12QUVXiZoiQ46k
ruRankaUiRsIOkNXsl6uJh3bQ3swjmIBl6QgxV4jF5O/j6Q4ZDei6OMKxwOoG+rn
Cz16DYgenn943bWRzHesaQ==
`protect END_PROTECTED
