`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SjCpjPmvXEQjnsqSIIWWMqnVsDWXAL1YQUbBTvnc2YLQGnlsDt89pUx/dsW4rWmK
oFoCPchvIMIcnr5ExqxvmvII5OrnA3hoIdLroN8MXrnntBme49oPtDbwH8XqUyx5
TUecAKOL/ALM3sagRKcuUd4HavVtgqJu9yBfVq1oztNHI2Kfk+vh9PD1wy05264a
qu/gk0j5Kj65zbni2GNG+B6ua8U/ghifx5QKuqL+f0EuuygavrCHPqGpiWYd0zkB
wa+DOeFtfJkIbEzbTiTen38M2gL+jLPNrYe5J4oBObe3TyHTxRms5h4zSwsbSHCG
k38qgGd0w76EZWGQsMxWF08gCSwoXBPtdcRhnbMlEapetGB+0tuOF20Tpu41gCQu
bLWEmQN2GWbSIYhHOm03lGdD1kBHjxM72z1r/R8svEo=
`protect END_PROTECTED
