`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9AUl/EFmPZz6Suiz+tOQQpn07oBVdwNgpX+isXCvavWPXEAceLJUVJ8AOt2lszya
EmB7Rt3TbIx9lBtmV2ZXH5CvRJ1sKpKu2gmIjiiu12ZmtOMax/26xuG2eR71Yi7S
pUk51/icyeh3XL32xB+uOlI063oBQ7eMm7mb1w9E8l4Pa7nSYSQRdC3fk3rYVl+B
hKvhMaOmbELmG2a/YnZEhz1oPcqLocDePlR8jp1FFz9v1FNjCU6Le/9GIRG5PUi1
OZw1BwpOb+0Qgk1JcAjpZMKNWdXQp9J6IXBPh05ojJl0S4RMW3LEPbiyNAnakg2X
Lxa/gt2kUXRSKjha2JhDzINNGhfiOAyTVM2EMMyz/mZlQ4LOnd/h36OHI984VsK7
vv75HRqWIwrcob94eyI+jnK/zDjZUTy8qwS+ZCcR0gZ4pWt2iftuHhYAlCNgGhVR
I2Xpwr4W0pehGgzpP1W8kuVRAvEyHDhfnOwNVAWZ+98s3nQsDotFFmTO+VV1cOcu
5MlYH1px7S2p+X90V3qVXsryecy12QoS/+dZAC7XDa1CHlbbhVMyHSyDBkEicEhz
xqeiTpwu5k1/4EKpVyy/GHPuwNaLA2S3UJUouKZBwkRem/xsrsf0ySSU25RtmwpZ
P/QFM9OOKSYeYHetcxKMVN6gdQ1JkcKzq5bmAYQbwTXcvVk7f1d59WnUE9yRGei2
pBAEo36IORldJHTMBdISMjYY1wkn6H7QCac3acdOdBC1bt019K8cmeBnAq1S541Z
MV8CZ1ecYUibpnYX5Eek/ej9PUHpGY8ZiwLu/iBYpzfqmW05AUhFOeKTLE9by6bw
CY6rDk0pSL6HNOnLfTI7CbTwb9TK6toW6rxMbnlSoBF99S6ABUAwHAvFF8FqNSMU
nq4SsJRgGNQju2Ak1XrI3TvdcRF7V8B9uTE0qJiKAM+2XvvDvp//Njn9wZMAkQso
eD6UOg5NzFzy8Au2SJw+T0PwnUS+0YpspA/j181K84YRKj4+YydNka/gFGLLxJK0
i+Y2uwutxbrGAuAGiGhxosotIO8x3nedgtQbL1LOcJ1kk7jhWPouaV0JMnZH3BYE
Hz4kpJS8gQN9vLCYQpjw5oiWxMnVtNOk1j94dkOEnhAIIcoLoJ977tBNNRlzW6aX
1tpS/vt0XoRiO/96ikzcz302/IemcPsUACKZMsEilPuCx8h2+7pjlmBa3zYgF/Y4
Tp+P0PjurkN5r7jnZ0IABhs3lSiY5Rbs0eFyK2VA9Gqm6YdPbfxr2hcV2BA6Kypd
7TJ8dGAb99ybjiwt+JHOCHy+BTsuE+UlUHkXYFMJF77cKglJjkUB1tkuC73byCTF
1A6Wo/ZzPdQ3yLwsuTVb5MP67dAeyr3hxBfP6HmonIrctKUr0zagTJVqK2i7ymGg
/wmm0NGa796Bt2NOaVF3Kw9ssm1CKea+SU0tM2pqZi99eYxlwIPaXgPBw2tXLKBf
L58QDsxXGWfgtNhhyV5hpEdxbrHeJYYXg8SBrLrJuRIxTkUwjI+5cORXvJ0+INAC
QtIb7h7Ee1P3GfEpqvOs1H5GtuxRNKyLqmaE+BDySldweKpcLK9Fq77vzV62svqc
cp6USKGxXkbJNCdZWQKRAbGCrveNgbs/XUmFNHvqgXxTkaeiQGOWBg8iXchmHT65
1V6+I+7zKKXJChHrOE/bFzfa4hf3FBZVepkg6cmlp83Znnm+3V4YKvrN/BW5Cwmk
/HsXhImBktXIoNAhksOx6zLCR1I5tG8h2S7BI7ECfn5tzkCTLOgKxEqXy6kFmG4J
9dd0Ib+qaFHZqHBG2FAb8Vxz0Bj70lopQOIAqxO1TpMB2w2uwLbzVcSDXEfIWE3J
aASd99XQaamICdyBGI8KVyEQ7W/JTXGyK7n5dN8QTWE0GzlGqWLEcXarNfnzdIDZ
5T8nj8rEXCNLF9Bt0M4BjDZKWov5gZwRz9w3W97jFgDvGZS/7PkFzsDIhrLMz36+
gmOV8pJq4DoE0TeM6v3APdzbTg4EpDji624FWXR/2VBOXcDI3/sG3MwYfT2MGO4S
DSDsbx7zRQCyiG/YJepNQcKnix8sPGvw0AoHxZtI7NzOHd48NaYIrGBiJTXmQAw7
5gZi2KN46eR1UXjEZJNE//t8hnZI26g+1ZKNakMCA47T1j5aqNvB4RvVv3tlEncL
M2KYqHitllNwfRINaumiHjjbpOWklwbhyZgBjXeq3SbMGeyx3pSw7u7IY2oIflaG
ccOyexygDMgo5M6pWC+LuBkc4PBVzy0mB9ArThPVfQikJsr5d9A13i1i3PONA61V
l2DcynWBQckwqCDOHx+uP9ftVbJmiqVBBUvJzfWpS+iggonYU9oQW5e//vQ+6ra/
Nu2CzhZHXZPGwMKZZqSBBRoL0R/CNAWVirxkridDf0aj2G/XDOVzy7kRklwWhiX0
/l1u0OGn1DtdHFp55UzdWW+B8yKqkIyY6tdV3NrIMudSj6IBuhy+dFGMiZLjzM7G
BvraEC35VUzOLfVbFe8ozXanqiKyg++tATP4qcxtP3fNLCrjfNkI8R8W0XW6FSZ5
D8QFdmLWDVaOxakicFQ7WlwXZTa6k+OYU99HPYCtJLEWnXLx7xBmElJ5w/0ltCRE
5kLRhcmX08Aj5SPXIJLF+HVSUaB0ju9JUK+sSJt20Ddn3YM4k5DzcEZ5dWwfPp3B
aAkt2dIKjM9uMAEe/CcgeN2Wky2AklYifa646HChVT0FW5+SWlLrZO+ixQK7/CAZ
xsNbysvXPWx6U997wAPTraeScTk2OUY1apqNof3r6JsHb1Qj8KI00ZgS1RGbh7Uw
L5Oqat/DiiC+iTdl1RDmck3eHPuyATg2AvoNQRrZY2guWFx65M2KAnVGYY+CcexX
VMpfgkC0KDK/uFX/r2Ehj3o7aCsqzq0AOYZr1/tBEmVjzocs88sVIhZX8AKCFa9i
QATVtVsJIdJd/zcpod7skR4a4U/ekBhvZRM4IQv2nnscvRlRlSymB4ClX9eSN6nd
+EJe5myJrsiTRezdPXLsZURkjPtESWbPPeNhlbdWTVEgBvBk5SpiLAMnWls00eGY
LqgdfMRweHx9TNoxI600z1ekZnC5+EdAqar+1lkWdliVv8D/VF6/V54QjCKCkKdi
YE8wzAnZ1v8XYnTzFGVNxOvYw58e6cLo39+ASW45LnpwFBlL0EIoVBxwybDyCwF4
9k5uQl0PRv42clyfydpGGK8yGe25ld3ENi7l9nIIvOM6C3BguUtmsupAA/BkKWzB
VsHzbbxXBvQrlTxUfCxCP0L5YFsent0cJHfFROYZthuJ3M+2t4RRg2Ol6MR2PTSF
plqRViM0hAeOpDZCxKMV4quf76H4ZF0I+U2RuUwIkjSdCn/mAQLAOGcTbfUnoEMM
clog4WY+OJpt/8xQ6DM4F84SdS2jrtPYn9/KsZDl9L/YjlUkxpx4g1LyqU1ag8Dc
8Eg5yn2zTm3107LGAX8i+Sg5knXmNDmvBKo+TxtNnBLL6+orBGT/5snoUqfY65xv
sXrpEXDwnGJAkERcxI2HsjqrUhRHV/mi+i7zgskceGpGdUt42L1cWEh8OnGsrRGn
/UDrc+81EVFj9YKeI7hQZ96uBVfGZAMFSgVGa7mwSqRJZ6jbSQZSDVTBhirB7yOr
n8J9ohsATwm4wG7LEkGqs6CEmZvVDgKveA4pn4Uqg+VyIhJdMF8ktP5PzHTcZEYJ
v/XJK0qaQoukm1sAYWNVYUyCf9hCIsv3LH+L67c3bYoDDXpsNGB/IjDfTVTztddB
F77LBYw5PdDR6qBwW6g54Ud/+Ne3TQgDzndiY17w0ZypvIdvAXdXgm8336soENU4
pGJHCYsTt9IA7B1pp10JNeb52fVHTZDSjnHoglY/bCR5ksF5cPhMifh0DJIwDC0d
M+zi8QvlG8eBJOYItXvxTDv5o8nwUcrKwVELRbCgZhI9LYmS53gkhyHB1oexA3i4
mw9AG/eI37uWZewCVXg1hsHk/afpnKTM7dX4IYWCP7EZxl/M+4vbNsak7ZWH6Ftu
1rJp+Ydv7NfdcqiJLdQN9x7HL5iAqg75VrIQoXlzrUs+R+AkQlrXOK+MmmE+NPUA
8VjwRYduqJejrzMfAlRZYYbI1G0gNxPkXDud64bWynCEFAxhKWgLNe4CxShDspx4
C2IpX6Z/XDbzQqOf3om4gyAUk/RBq6ZGfiAHwlnrFDookXdf9cgAIJD6c+FkGHE2
ULcLI3SLl5UvnlLLEmkTniuQWyfRKONYrJbnXLNa7Nt5V2tgiUt6SALVmZLuTQKV
BhCowybgBA15c0T6IEw/in9vRaU2KBoeOC0Sl7evSY50BUAcMNNgpgXTdrIQoxYq
xA6Tyg50y65Rs53V9y+YU/xkDHgePDCU0qzkPaMzfDA+ucOdQlhHKkPDMjG4tge9
XytPxYQyVFrXy5P/Nk5hfaphgTqwmyKt8AwjwZ9LMDFqaNS8oS69YWv34rup1gIi
pbo0e9Lsd7aAXs0Wvxp/NVXUgZQfUYs07jbiTAsSR32m09Drs4DUwiNwTvaLlqOx
Pv/M75+d31g+IMdbMXb5LzY97MNJudv+xp2PmVEXoDBRBe3n/w4ZvgmzaPItlc2X
U+YEtGFYhArOW0wSD4HphlMhQL+FgAGX6i5eQKlBoPKMv47dEiac7WL8ulJfhZgz
fIp/kwtDhAuFkPcbsi5zdzwKljQw3VvF06kNJ5kUGasvtq14j6KkJLmn+oiyyA9M
2ktvISucAv9kKSjC6N0JwH6SdwoIpgZgQKzH85JGsGzjU6bQxy4z9Gp2SMIjKnkp
8O4sUp1bRoWBnonMElqMuvrU2oo6ySAW0zil9TL9L1AIsGPYTxNgQLaXuSHAJIvD
fh4OH9pZgMWdMpKBdhCHQjM7J2xGkZ1TPVLARvGLkkxbqCJvoBPXPe71u1mouCnt
yzu5NiBphqd5E2ETzexPdkvyz2Nsq8+UXdJdVOVgOqTpVeSVC/jhH9J37OZ/02O6
MyIPIiceRDl6XzJ/JQwwdKuG2GGYP3VEKxFAr1Te8tRXeGKptfrw847A1rwn5jOd
TvRsZo+yiw7xHoOloOSf2Dade+KcS/7jbP5DdAa4SmHqeOORj2IvoWN4LnC5cs4x
XxGGiJ7dEy6Ms4jjEFQSXnCrvwXQ52AlR8HGkNIUup+tboXdeTBQQFNR9w2KUqDy
uyPYGvMhVqGqIm9t/yzuxOAECZZZBNsMrWCHtPZqDpq23p50s0c03Cs2aXKh4v9V
+ZC8Dtyv/qwXzzvlcUTO+r/e6D79Dn3qXk6/USTFDP8altTquqgKtM+zYCDh6Unk
XbJQyRR1okMxzW9ueCQFl2/Vu+zCShSJwPGDeMUQRj0tGl11hE6GbqQLnkQPk9GZ
v3fVVgldiB1eymFKPPET7HZNITdN/PYSe13ON+PBO5L2Vqa9YlEaDIKCFffnXazC
fBRDNEo6NH/RVT45eL6jCoSqiNYMyB0TwH83NfDjsSUesVW73I60KHOTXgkpH2B3
uuLnQz1ohpNS3OHbBF5joEm8Z/ZJObEYc1+ny4g53Ym1jBEtKXelMIMQiacxdD55
ywHzn0wb9Uf3Lt27PBS4z/vjfX28Kb/TUpEJbRg9As8r3klszYyRgn8ONQRv2XRt
+asIImGPeQ8nJML5uAMHeQE5JO+6bB5WOlBUYIDtIr153QQvTsF85Mov+FeAyuFL
qkF8Gm12t+pz1HdjkTucR2cdqrZaydLd31F2/yhPPbxLBBUjMZFUcw061zkEWNlG
Uj+XyfpPB+EBAvbfFlUiRyieA24QowL4g3QsQ0wTe53vWbct+lw5hnlg2lmNPiep
rsts7Q4l1qTd/3OYx37TbCu8VntVLqV5K2xAv5TRk70I1AW7u22KK0iPwACcdk2B
TCV4yuUdX7S9JSLyBrTrrsbQNOTkHVJ5l5xqt9MDvqcwECOS0RG42CwIbxmik/xZ
6OufQ8Jkn2bWqMdPTwFFbDIfoYlRZO9GqfiNCvYgsZ+OyDX4onutSHSwXnsfbjne
ha8tWnNWVY/x/IqveO57UZ8b2Z74jbJbAMWS9YmhyBUd7cfTem5B++mzXHA56SSX
+AzLo22jxPUxszb5f4qZYxFopS6sMTMZJbgQlmovHdA1qa/fblMsZ/WX013vrbI8
L9M5DVkS7e7sJu0ENACXB3weWMa8r4rrFI0lqQZLdRzwct1NCSvfUS3OJuVScpUO
RPJYUwAVSZpXPLgZd7mIsEbpLYRAU5J6iEgyYo7812/oB9f8BJotDOqA1kCYnhp6
mTW7SWJjwNL4QwlRvy+Baqyz7aWVZytfpyJpjAFehTPwheETSkk5r0SVZptjV+Cd
8C2OiDWUNNdqyOxPU29ujzGskH/R67N/a2YXI+nB9/Ri0lhZkAU44bggf33VFNmM
XBy1uUh32y0I0Sk1bDk35gwU16R+7NEINNJZzUynYcEDFobuU2rr0h90GetcSCZW
nPxRW8secat0wh/3OC+RGodD9BgzNxrbT/jETxJcouq93DZl1arAKiN0FN2UOaUh
ByhjZCHcFDFGfRhCOhpkmz8Z9rsT5nN5SoJklYXxx6fovCkFuZcpS9JodAoDsLQz
xYQdTv6JD+ZZUdaubD2iVU85Dw+D97IA5xkASp7aNtaIzHyUpDPS4P5dSfaSQsSO
JTQXbZcBfS+sIwO8L7SbQ/vvqYugEmj/pQXjpcW54utbpgTDBggMYmHiRAW7vGHI
w7K5XoDvOHQwvwUvATDW426WU9+gvlTPp5tNg9cOeW8pFmjMfSHEOrxdLo+Cda14
0O02+DOcOhlT9sY9G/qHQ0prtezfbpJpskuapuN7/go7LRNa9mGDwivHfXCdGGYz
oXdhFhe87/JfUnX41Z7ALgg9RouhMjqX/hKT2U3A62eXkXtB1+ScKyRAvqJi7Vey
D/4cVCGpvkrOWPg424UUIHlgjF3+TtJ25gavWgGlmsRka2p/fmiX+y8AIT3ujjeE
pm6kqAZYNYrpRf0rdYdl79WoM92f6UgofMTQ4aWbm9vMDkYGeQPTtItxkvz04mNK
XGf9Cyu12jIBakmgwSzUl+iP9yA/r6hsqMx6F1n7oaZPZvsZN+zN0SmaB1Sd/UwH
9SZ1II/Q7zODx1MNURMoHQbVvWM8kPu013dNOsSRUJl+eLmAB/yswp+nQZdISqLy
4MVTeS293xeB2byItm4BiBlbgqYZmXMmj8oiKeOsF4pvYQ6gpx3+FK8QkcMddRJf
bYTwZu19Sf0X/zzE5DI6Nv7iFVisT2T4VcjQ8crtAbhBSYgcwofAmOeictOsKIdJ
lr9M/v2HYc7NFkmjTLRYxK0mbWwjpjINoGo+nNhV0+WOEw+HWXoJWqkMYTN+Zm/z
xbpGSwHbFLvbWthOu+seroIb6PJ7X1Wd96zIgDxcG17mCMHfQ1YcqQAic0QweNyy
D48TFSZ9gTEAbt0AUGwXWqm5otacfh/HV42VgZ/ue1LciOFqe4zga3tIG4T81X3l
jntyS5aPxl5up/l/khWAET1VLRKEe9pxhUuQSA1c9+lxJ4/mFg6ShunCVbfaacCL
jstdVcpX2E4ODvKYpWrh/kITQ984npwR8VXuwf9rTMwMW4PIkq1dS/spWQbEG+iJ
l2k1kxti6wJH4VejS6ypO6mh7j+nMJeSQnRyImOFxG473Ga+jk1jAnC/KXFIK95f
OA1LeBUdWBDxcPq8UoZaA1Qo1n29gYEQSTzRfTswHAC/IWZwXb0mzU7oNGd1b+L1
eLdV1VAa4iqI2crsmNuD9de+DS4iqG1Tz5o/dHCmaZWsLMgwgs5dexMFEvE3FR8W
2veRZZoTj/6dVHbAwKx/QcESxnao/0N7y51bYJ5fzn0LrrUw9lHEot8dN20BdJAz
KG8gBWd1Rocs+lFqUvPw/0UfJT7p2mhe3oq9DxzjLZ3Tc8qywD9NZOo2DcW1Khn7
TJm0+CPWkCJuDy8L/gAbdtTucx3ZmGYzaueHq1oVWbAqOubZUGUBBgz38HiWrYwY
JljzdnwtaADD7O9diEEyNiCBovUZfzXq3unUqMvcYxvoTdfdNoJPY3y5k7WYRANh
8pjj1oLpHmPn/Awm2OgiCHeivTpWXuXn1hIO0xrJ8mpALeyTd99W93SgDZTDk0Lo
pJG1c4ByzkQeCSmKkpDRffPZpTVoz2QtNRuOoijI8xsnPWo+jyzKVU2obfnrLQjk
NMIf8YM/Do22qKCa71YTWk7U00K8joZAJf/kvY+z6c4WqSdS28OfGcJwGd1Ufsfe
kKUEOaqCiiZW7v9gMSaniDH2IC5ud/CrkObvdSQifGDGo6qWWyYa7Os62Fy8sLAZ
x1Ix0dlgsHnzkGJAXl7Kbv0k39mtrZYOOt1pewcyGX/e8FlPJDNzij/xKQ33MhPn
RNLVmffjNiyjHcqzH9nN93vGy68HOGpTjs40CLXS7Zo4PpiZmfShzZB9KTXx9Z+a
bXoA9hb3hIk0QU9I+Gl7WV25cT+d732KH7A1FRvoMTanGRUbc3vydFXsJF4NY54A
Qdr14IJGd3HcqOWn+YzKTyU4TK5Bz3Vh8+EuNYB2N8TgLO6It2eX/WrJNMEqKAdL
pI63OXfCsQgQJfdIeuLB3gjaBB2VWA3u/q8Dtc1cx5k1+6eqI8XQt+l61H+weUXC
2my7hmE2wOCtaXa6Q2iGyvKaWL54kqzjuDXW62uHZUnLST/T4M0c8tDQB2SFthGC
VAkW9bNOZExP+x3LxGch8L3z7MOj0VpAX1dYSFswuCtmpgEWSnc0ApxbyXiUx5jJ
x4zijtjA07grOXj3OdxCZzBVZhC18sUtQ+nAOOnGg5LclJWdrauhAbn5b45FueYU
qHo/1VgHxJ9Z7FlH/I937FIkvz77zHikCJA6bNj6A2bi04xn+hA8bbgpK6nY9jDy
B2QdxI7iaJ5q8t4tp+4pwZEybKfOb1Ick9ZsDAj+CUPG6IjB6YuomtL7yrZm8J1t
LVQahhKv3CCB3zK3wUAvuQptibTEUKKBX0gTs1wia2dX9ZT+52mTeAQcN1AWqjrc
hXl3+DFLk6cvooy9VNIpUAM7qaDwJ5l6NWRDFA96iX70jSBLFZdKwmaW/DnzixuM
OQHw0KD2S9pNd+H83YUUUWUAAF8gYuP77m9T4kKy3+lh6IgihGxxvGyUU1br5GfH
PlGppOC2YXBO6dCxH6DPqQ7V1aN3Yspn1chBELCgS3fWiNw+Knvj2W3LtLEdiTvP
pTkpF0suvPCkhmnfby00FFbemO7lW/Vv+fLRGJa0y3/Zzhk99IULKj0hPOIxvbRX
iTpBAHn2oxRwsSshVOMMKqRH1JnoVev+WS1ohMOGU6/hFg2BmqzC5KJ3BHjjKJx6
AWBA0112T4dzq21rj1Zk9VKV45H2o2PItPfbJQSuhaYV7CS92wKi2zb7n6bnh8Pf
0Ji+QpQ9Q8RTqSTtft9vyBRCMKsMBL1VjJh4jlwB8Z9qyxdPBTagT9QB4BT7jzx4
l8VRC1FZeuYBw+S6lHVVQ26ECJPHjhlnBmiUfaSDvfy8Wd9rNVVc8XWEV8qO3oo+
zCJLmEUIOdNXD3bJ6tB9GPEP10S/b30gWnK486uwkVz6sPnSVLP4xSojMzZbpJQu
0yn1eVqvAyWxtqq32Avj9Fs+1ahYRQ/1gnmZwXslOf/SC1Bo1RBtHWjJdBgFKcTj
mvCiTLCokk+PAUOglTGcCEPxWqInwr6yTrzP8sUNoBSHW8SZ7eAYIQM00+Nog/Aq
01feWLNYDReg1wGZzwHwCEnI9rtxSlsP26sTAlm0p7lRLIUXAksfcZ6J916oCA2w
vtMeelT6KnaO1a9KAsOq1Fu374jGYL25YpRZQ/PyB+ofjLj3WVcybbze/S7dukc3
SHHK8viTuQFruWRLreFoiwwqNc7d8MVkMWE/rsgJI7U6zL2Un+QVGt4wB0pvNTM1
+XxhYFIY5bgNH/WVo8LwqDzfE9necfOqx7w0AgfnmhYLimJ7eTCXLLPQ4BymWBPM
GIhVOAf3BO+3RaXbmKVIcGly0chOIsm9hMkvJMUHV7Q7jcR62nPx1nDHM+FRInGN
z51gOeaW57MFNMSzQXhD72o/ek0PL8nkr+ZR9/nz09hN+m+hOrIkvDGrbU/zIgm/
Btd+9ZlklN6fnOjKO9kxSWC4Vayo/d8llYhUNykwUlBniv+nowt568C2d/n7ro9M
9VX7gx+mw+LZ/KbxQxIKskcFxLd5T9TyNdYTn6EHQjdFH0SXuobMcwaw8bTIcnvw
bl2NZ5WroEf3TDY8tzzuFvdZ+5eCFUyptWIcW77lt8upbH0kEGrh5ssmi33xzP5+
C6P//64RShQ3Qcui/eahbuFO6QDjEYe0MPAxktqn/l1A6OByA8Sh9tGGXBNuEvbP
nAPjdzGDM7+qFpdhPwZWz3r4aZp6Gy6TwkLNRZMmnhcJ3s+T12pjQWuVmDD5vSnJ
uyFrz+pYNi6FlObvHX6luj3Mnb/TbOG2fL3u27N7fxIC3PvsZ0F/KMceGSiHgdvZ
+BiG56qhHT4Qn+XCJTxILaHjBxqMTv8Sh7jj2xwExm+iJ5/r5rIl3mmwA/me7Bnz
q4bG71LOF83wryGIJPYX72AdwfG90oH47yUI3U4W2biPmxnRBaNseKIhiZVJU+ZJ
gNSWosJzrTAYSWHLwuuvesezlZX6wfgj0qbKYg+99xPpVomxdJA3Yi7IVHHVnw/2
JhcK4LtmqgVaffGL9FA9TuL45lHFSBZl9gHMk+gXDJZN1/VHzQT2xwcAAZaGy1TS
jo5M3+DZ1yeFdc+xLlQfluK2U+b2B5aUpWS1SATpzrAB+ag5f1dRZJnPw5sBbIHL
pgKXNmuZAXCC3qzr9KJSMtez9iwfgF3E2pWy5QP3xk7cFU1+DTtXjENZdLdL14+j
eBurJufmcM2w5T0967hQjdbN1jSaZ4qSuHR0+AHVULK6pcFQA4AaCtkPHhSooJIH
6Oo8WpfEn2saETdIzJPemORi/id7fSRh67xhDhu/6pBrQpjFzF8W0MlEhr8c7l1+
IluCrA4A22BETSSRJjAIuIXY+uQNHpcaGlifKFydbZEsVTjtEF0PR8UJfI6YaMNc
56+eOSUZthWdIQ+OZuhqxiwumRFb6TlMx50r5s748xp0VbddxwDepFyoaF3/UfZd
mWyXy0asHh7iBHmOZBztfWNc417JCDvV0fnREiSEnmtkD4zqtF5YZGLbXYprhMU8
l8eDPTe4ieX/n3ukNYnu92K+BLLnhdTCl+ZQFLC44x1jqtsWWSiWhntrQ/7q9GOe
+I1OxB4YPl1DlRC1HsELHzOA12WDYeTxR5feDIXLqh2C0+GFgWCZX/VNUGRosC8T
lGCpTJklMxcp31Ne+GLVHLsPVjo93qCILmgFgA81v7JMXsZSyUPMJutsBa0Ngxpu
KNBkYg0jV05V2m/bmm3K37plZPPO9rMUxfWEgmvmPSkVWR8zvi425ssa7ANoJKEk
OHy/NAVLIieTMISnS9/hElVTbQ47k6YkbiCbUAb7MPYp72DKiKUcniAPpQG000n8
UxHbC8ir7LP9/Emv1CDrYOv44PBHIQFUu2k++tmt32kTAwFCnXLDwRMvTm4Q7cTp
RmJTz/+edaYxokYhr70F0kQH9EPeVjjFzjixKhvF6hFPZe9BxQiI1ROMDNXgiZJ0
zMZmibuzp9biUk501sy4JO4/TYK9f76geIvbro0I9MDQmbki9vbn+DYbQznaE4ru
SnbBbJUXatNzAEbv8a+1TL12Q2JIRiqTaaLXvLTmLplaYffVtT3C3uFjbjXhrAz5
XFnf3b2jiFmuchxNuFmvRCYiNVlbBN+nsOh3zKR5lAsfR6ScTVUktjkPLZje+eKI
uRiVUt9iQlw4OiuvAdrvjl6GcXEYMqljNOBavl/P57a/2HHWr08y44L9Ne65pSKx
y1IB1IXQkZvlK+NQ5KRigGaYhdfaCG4eiHRcUk8NAdGDn0vGYF09IovuALnqSy6o
dUKMfSQx5tdqpjLmlintJu3IuVMB3Ce8el/jPiF6CD4xOy0k2erZUchioYr/tiIe
kW2g1KEaVMUV/PnD3CayZwOsGJfaUUzgl2RePoszvmkzwXuUtb/IhunLD/IlMPLz
/Cpw2nkf9SzI5O35F5OD52Y/4AbZr+Ih7/FQk5M/DNWHYLEEFJEiF/TpVJjCgLqZ
FEhPMvRKzYrwbKx5aSNa4aFZBhQwJ04uSf0VxhEkJuynTz2OyBZOTdOhLa0/es/d
+kl68uFKCoYO0xtUZY+ahDyqXIqWjQSlUqa3SfXIrF926JhIeGOnK1umFQxARWlH
Q7XtUP+RruDBSgATo4hlN7bysROi8r2xLQIDB1iXqJWwTDJp3Ee/F6Is7e4SrVbP
KEkWdrm5Mm5R5uxm24I7lGTcB+fKLBpVfqBbgqj34wQEe+LZAVtbe0W8XgVl1d2/
6njTdsgV9her7kY0h1Dv2B1X6odnwcND5swibdF8jjM/LdrFn7pUDsQp3ki2mjSt
BkP6KJnoo96yE4m87DfMxT+m7Sx/CcITAALDa0PnsQ3183kASs4Eh0oIK5VJdfmK
5EeMoVJj9onmvmiAoeQQ0HkC4Z6qmd2IKYWlYv3mmTGoQfBzuecwyRo5h3q7lgfU
AesV5MQxlSL30XXZOUHZU5+5pbr5dWLaylOq0aIW681d1wnYlDB/N0kM3d6XekU0
H9SaB4s0hzIvndbn2DB5LDheZwsNxURkDETZcGiqIbQP5OELxr2YZZfIzC60VzWU
wLBan+/H4Jz+SPZFTdpw/S7YML0iwZABN4iOqkfFuzthTv803Hk2LcVYam8d7Q3z
eeiT/IKqMBiD3qrNbClIIe7/8Qi3szNGCDtpj9hINB37P1WNQgr3pz6qrZ3ysWGM
2MDRTd4hMVhn8Ysr/tP+pDGPo7CyvUGpL4Lx5XZuRNDjkQrSM3HW+psdo83UUPLi
Y67V2VP4HplcqXzFEp9PTyWYicN60oXyu6cUPT3yMmEqdp+S1VjPLjZUFrIU6WCl
Fa5onB5sDL2LWeKDIJiLNB3aXXy2jrlxhbG7WEhTlOiGx6WE1uVOOV6vnmTy13We
p7lo26LiXkYY2mRtJvDL0Rk7AZ9fuv3Lc14DB37G/Quu9OACCIwwVBgfZwtOtlbo
sMnN12BocpDtFt5ZJ50r/hOEhMuXz547ZoBZXweb0UAobusNXZqC2Q92HyQyu1yF
ITyc8vVNV1stqyo3fAkQgFx8IQOP3/PWPYXcr431Rwk0CFEC8ZdlnhQHiR+zsk1e
SKFOg3iYanrqZ2MSacgPnw0Gp23VhFGuPxkWsaiLK6lWydq+ioyb3IJXbcmvsme9
j9Qdlm45NwCqkTwqHpU94+DlEvc2bLaqRqq70a28uCH+gEbfvIqrIgwa5CpRXSG2
/Y2ChFosLoOq+47hJUqFWVybOf8qNpEvdo2kTlNhaQAo3fVY8nO4jLMQ4EuLimND
+hGZyzXoUUdAFUrm/C6AMxL7KJ+yFq6HvfyV/ax+Sz1bB4Uw6qB1slYAM3/pNULM
z5hqPOQVQc0ckSlQ3hi/LBjy9k2ZUUt4GYDIc965QF36rrzVVWs/tzBw/wpA3E7G
aDkEZLVruH1CfIiLmsbSYfh6Jl4FLu1vt+Q233bkACAoIdiMrLEvPoq7o8ehuwdl
DSH8kqTkdrKl5JLzEgRerRjbKx91awOVH6AOaS63/AUnHvI8cab6Kw5uRJBAikQL
6Ue3Sm0E1abDzau1EiEZk3sj90165w4YMr8Tb4ES12vN4LQkLu9fSlsc9PCzjPys
ODQPIcx1SfuVTc05jaffsL++ikNfKLLy7srBfP8wdIvsSYsWTsHwlhH/Umwr1Q6H
pheFLBiHDcpMAX67TY3450qpckHMuOFMo8Y2CXDtmJzxDk+NHfvtATaS4DFUHFxH
tAjR98cB1KDXaAxNlLoBEeTsAD6mlKsYe7DnC5AqhDgw4sIwldJhxhVMBiB8JKXl
DOMTI43UXNi3M5ucSQIOUwoxhvTJ4PNIp+kvnY6YYAY8nDVoX/5LEOOU6Tjb8iqg
NwdZQc7JQ5WJcB5h5zeF0w0Bt2KJOm7Fe1F/c3ROV/uHFEaZPU4H8HjwHhy3QwBA
oIbCq9QZbEKZvkdFmWUDyNB+GdzRgYd3IbGdB0TeUwmGiOxZhT/wohF8P+izRPXZ
vvIDn7vRB/wYC/cvNWOTiICAIVTr4d7wYHavoq56Q3SBxPCndJ/6CFna8AaYSbFz
lHZqQpwRnL/ZkKLTzn37y4uZ7iMd7EQkc2QEAXMaOm3OuXI1UgTSePWlI2fHoy3J
0dbQus7TkwIDBEFe9YAURqS44hTjCMcZYTA7YH+cWXON4HVcU1V4RQaIu7mXJpjd
MJSzpfktL6dPCE4o000D0RtdMTDqbF6ugjnvPebyV8MPZ/JtQVreVqwNnbbLXMoC
KA2jzKTnbsowbqkPH3oJ3e8S9uF6q40Bo29PZydwLy2pwx7IVJsYMfNxmQ2g6X1a
QiuaXScq8NZCgLsIjChqfAsKGoiDAfg1hICi4tsF+O4spEnjia6eP2UQMI7XPLZS
Pm1z8GdGHpz5+RWQCHbFXd9bSeN9JJ354Cm0KtWuLm/LehZA1Bgw2bnNFBZmVhQs
Gg6HYJt0fWS2U6GCiXWgwLnORwOhkO6b5OhUvNGcFN9VYfbkMuZyYLii5GAW84HW
K1JYVQ+ZCyLljmM1jkuzEIIMVdwvdjkjAy8G/qTxpJjMXtmwfkInRHuQynCZW2+y
b/M4EFcXAEwbxY7ys6P/xtjwINcKr9PTKjKLqhKA9Z/jYgSQBXhD/4/G5Hvme7hk
NEoEyH43eUtsedOft7S1bveiusTm6f8ZoFP4wr0f/C4tMWGv2s/J/qhRjq4seAuV
n/3QmyEiN04jzJRHlMSer2j5glIIXOeLF5fdvmPfp14GuC0DYuT5m2XYCLLNEfiD
OYmDkeN3J6yaXVigpYwVB8Rul4pcppQQrkQpCq6UMalJnwO7keDTP3Oz3vNKtCMD
bmIWGekvppOlU1bS4LCKOkFQg6QS4DLe/AeNowwRvpVm9IIiTqYfLfB7YfrL6t7k
phPLLZmK5ZrTRkCOLQAqnpOY49EfDDQc5e505SZn6KrDXGu54y85wBfC1AqNc33I
Es4nas8xSUFmwEn+gBA+4RkILmyKy6SzcHrWtYAVUb+MVUGn92iS5L0vVdRKLDrM
6I/L8ahnxTKpABm7RNhmOA2zinqE9MzFoPUu/eVhfenex8RdEYb1bWd6tGL0xxq4
W6XpOOksWFMKlAJUzmMeNqlAz+83GDsFvjUmtcHpFBDg1N5txYNUnooe2D01M9L7
gR2t6R4EymGwHWE312BBQcHRR92F3wPALPYkm8JTBmLPLh4UFQ7SQn0PyXzveGlx
zd5NQKvcDHwIgYtHI0yBqRhqAo1pwKQXyYSy+WkbJUAKDk1MLBA6brIWQhK0R3aL
vPyd+iC4u4kBibWL5Zkhz7eB1Ib9gph6KYHQ+VEF1WlT4Np9TSHeGK+2HmRa6PU7
Z1PldttC3O540oGbDfc4EGan7hfeQ+PlmBImkyvZIUn5oc+JPIwyvwJeHg4CriUe
Xe/9/94A7k7jz/LCn0Z6mPmIjTK8gXNhZHgYbCah3lx22dwYaWD/+vYpseLLS+HZ
/BIDLaF4jS56eOWybMQUYHaX0KNaYbNHbMBHvB4ojUIuxPTiVahHYe5EDDgyd/JS
mKiOWzExVBJTOPLbx2zdWLhI4rxDeVu+KysWDrWHurczWSL/t112UTAvp6esKGLz
ou6c605jimA6UA7+FAFjh21ieJUL85aMRxVOLHxi/yLp7SDS2UCnSbah55y2pmDa
afCvA/VAbA3jeasTpdNRmyhK9FaJXJr0YmFwmpz1bKXLuAvPfEqeoJsDd5O8JBgx
kAJkxnLbFSPKBCgjeKd6o1vYFdJsP1yu/q6oApVhFy39gzH6lRtRVKbNNoKatMIV
LiYuGjpn8IEPpuSKMZQcVmfcHg78hl6FqfO4xb2GXGg9ysjseHiKyvZgHspV2qKF
ZiEnSbM2qnok80ivjBUFpjW7njTQwyqaRVrcZOYtbfr678g3h8lnnPgq0wgB3Z6O
7VXlFUDzglG9F+Rrt7wSxAzhEox8cU/uRqWLLWwrzlwzkCBh9Eeh2gJSi1MQEGwF
/YElWoXhYiTyWSkHMt8gCkdTL8nmibQIWjEVSOlGktIGhNa6+ksbsSSxiqAiS4kx
a2T74PiSEhBkCgSlkdljIV7TdBVbVH1frG2d2OqaWIOl5bCm5noVGv2ktrU9mlXR
QBIoNBYLfDby6/a3kPjs2vgL9pSikB+J0iItnPZh5zy5tvf8LcMzcSskNLenVQ56
MY7+awKQgjiqzsMZu/1SO1ZiGX7jz+ns1oQoX+11jCg+hXEMeJF+ITIeG6NoTsMQ
5Hofv8cORydEqg+NuzkHcTquGf9jLd3iWw2MaagnLK9jvd3B26Vzmd+va3a/ME8y
puGIqD4z0NC2FHdH9yfCUYhsTkhlbA+yTqOD28Wu/sqc+XkMWMdbkVClYd+Qn9TT
u6d1p114Y2GVK3IS3x3KRD4EMj4XF4bdwdoQgLvw1AEk2kOLPkLXYYyEtmEvhNh8
z433XGSeb9MvvMfw5kFf0yCGB5KJgn86MFlgWnov5iBvSrP8I2Bx9FLZ+T9zY/ZD
MUi37IY4kVJN+XQ+fQ7339o+ZvayAbgT6eiLp3xnAs8fpYxcw9Ck/nSgwJkDxxKz
JN8iREH1HS2c3Gsc3pWhMJFsv+tS8uz64415D8V0OB736u32kF1UEoHRVzO7I/VB
tkTxyOWZ8HmaVD79fhqwVNQgpr90O9rDSRFU0vtZzaCsZol048BmAi32T2SiBpMA
5OmtJ7IL2privHcJuKt8eWa6NAcLlaCzXwxoaITDv2N/6YtUSObtsXdnPu6Qxodu
hkza+v2hZNM6b2T+f1OltoQcU1Te8+QoHAbCF6XO+v9zrxPhjLFaRy/p0LUQDpdO
zYcCUFtkCudELZv7lzhNJQVwWhxF5numplgpFLAu6gY8qzfp+CUh6NrkE1wBQgMx
KCMnrAZvICQzyCpDEsI629lumFIxMLXDVmzOBAbWFh8WOg3KXECkiglqfWYEgqOF
alK9Ejq1Rd98BvCMV2WccrBFVttDi7YUxd2NX2zbL8fSRx9tZ5f8HAkutU7lmUOe
3rBxpalE12hvXWtJBxsw4hkn2AEl/DAEQWOzb9EWD/VX8XLFdptT/Wr5BQvzbsCc
EDPZ4jZDSsf8RMGDXT7PhRAjMYfMFY5LzqwZkYSzgfagFrCHUmWmHGVjYmYJi72z
UF1zF3bUEuYXKSkR+Yze4EmsoFaI/68wsfpUiRZe6o2otfRgm1H0dafHab9cGB+M
xvDEZ9sOSOb0k506b1I9h416fLHQFREj/2aj+G0MZ98fr45DPPfAYQVE4Ab6LhrN
np80kbUvQ2IWRM0wtnigBfIKwPaVVcpazkQGiikzjkrvsYiTEvDrPt2VZG5bAHwV
92ONxOx72zJ9gEpeVPmusWebYlSZx0WwJPkD0aBAsXukAIpnhrEr0bNDWX0CF4vB
BES/ZL7ufSNFZh8bGCj7LYrVP4qGQAeJs5PvFKCjhLcao13SjjWf3noPLfcNoGqS
WvI6EBEpvsDvlZAEXr6hKeNNVZK+FVxddcReNIYK98RbG2sHQKKO1gLLNOjVtPYq
dNUV5LLu/MbTXepiUdS3RC3ZWRnhlRJr2e9xOP0HjVJvl8fR6T7D3Gahm5d3rCDs
KM1P4PsnUjfkfylAvX2/T2p5IACgGon96hlqjmeOEXraDql9QSI46edcBM1wnPBA
4XkKw57YAtUjHCa+BaIZJUqElvf30pQ7eZ79ZuBpHX2qsficE3r8rMipW1ck39jC
lOW7eEeM1xs+w9/tydBdTSIf9QjH21KGZKFp4Fbc+8GsnthSCCggv/AFqv2Khc4m
hZA/NbcrglZ5dxxaPibVayRrGMqyB9vfinRWHO0JLVYhsMUtXJYL1rJ118WFQrTL
Ep5W2Wj7sJQKkZTApS+BKUxKmuPq9GkryAWXHoqy9HyNBcyA/adc+kS40wWhP1tD
DB6LvnhEbGY/hlkclPlReujoXuyo/4N0kM0mcAan25HkkkvsZy7fvdGEmGMehwNH
v/w3nUVfdzQSspRlxcEAKqzTaaSLBhFpQjenJd1je5mXGd+LNBmjrAEAenGPCahD
IL6OXjdz+995mWDNDMo5ZGByMmzBYifk8OadHxg4/YzpnxdMYsFnU1L+VcJ8NDci
k6KuKA2/meVPlG51zm/wlste+MUHaonlrdusuSzbdudg2SWisuSn1LDP10qjYxjC
eRG7jywkkCnsAIvot15qNQwkoJsD5oX5xxF3wsvec5ZyjZRnBumT57ksDc4nGOYT
FN62OBwjdfjJ8AVa9yV25OyZbi6ogKxv086vAdNItfs+b5IIFGqsBavEmawwwZLY
yXLlIEAEfY+KZJDTrsX4V2YJi2I29zcXoiKxhZV7qnh3iZnwW4ytxlgwY+818lrT
k+6PqA0NrtwbixCwb0+uwOjlC2Oa8ETIu8aZWbn9ljw2uIih0wK10hIT27Gmjwh+
RNNbJ4nwbymurxzo8iISESBC5MVWJg0ZKb2EmNkWGS/Rdd6XCfX6S7FCKnbVAppv
ABqV2J7WYPK1wvQ5M8Mj6P8CgX2EhIUk7+s5VT/OYk3RdnNbfZ6GazorXd1QQ91R
4A6MVl2fyj/bdiEEDAv+EHuxuxSX3lZ1gE3gO4wFE9zzDmGEUxc+aGuYtouWJ+I5
9lMXLAEjtxEVQAKB6j+V/EaFXPkajS+SAs1oq/2KSttxjaAcbsY0a0pcJE3X5tVG
PLaVnVwnIUFwt5bxqc0ej4OAcbCerM1VB7ZluQfj9P51OrN7UampJs7TKKRgvDwf
UZKJthbI9tW6qkUMVkvrpgbSuCTiRGT4nCmq8pMpLYJkBPR4WoXRX42/ftZFtPto
WRh/RviXgHkEGeegu5jHNxukvxZ/RAoFTqZZquYHwdEuEAGJceO9MmMZFYEublSJ
0vMQ9mCVvGBkikRqRS1pAdlqFp0uoGTD0jmGgGYsy3UOMhFLqNkRxzfVfCKS7UMa
UeJHL2UfsOEtEtKCXeTyNkm0TJtZwt+aU8B1QSo/HzvyUsKAUpydv1X+BoJQEnaX
HH+ddwL2LYagWWEXu63Vlyxip3FoFFT52O6q4TArmv7sJspHEBRxOF/J80Gq8vQ9
MGqvhxcV1Y/W4XmGKWakVnDNiFPe0CFan4TpMdHPbmfFrjp/yZ62cVCGhW7Tzq+N
Tt9Lj/yDAgaw1pe8TTphUK1Tgk+NpPAnDPR1c8SsNfxsQFlP/G/1TAytRIkRjyIg
ijKOKPmjT3rO3XWBxFzlYRx5ow8eXiMmMgu4vl1Inbb4pnQcBGXCJAgLJGB1njOY
wa0+H3cd+GNxglj15LHsixrnxabknM3oUO7b1kZYI7QTzAUJUP9sAWDKb4lp0TGL
IfJFBJFquf0and/3vE00qaT0K8NfA99NdyB8jM3BHBDdU01Y1jxYETB4MwHeeqgt
C4YnmRAvaIlJdTraOOypS35F4fUEITt4TVcTePEna0vW9HoCYiuasPhdKtP/l0As
fDyxyOwohd2+oFH0TTTfPPV7Zhxfdp9bxgn9UpOQX3wYyu+thWSVYzNPoosDZmrU
emEVkAsPjL4YBvMa0yUqd//f3VHQi9zf54sdI46OOmuNq1dH3QxLUK86ks99COl9
zY72Rnik9eS2sCEAIzW+dFOpGvO2e9ECv5wsc2Po3PBHY1EEGAKyWMTGK2elmhl2
1nRNpbZBfpXeFpDTem6WZgeuGTkggflUd3c3otiKqdlA/HHPrJMgQj8LGStVoiqi
dyox30OPK9ZDurw++R1kq7Ws8WfyPlVoejgLfuOdTgmHIITG/d/zGj9urdENz3J3
miHlTKkDQvNbSZgpfmUv4mnl1zT1hEaB9i7Ur6Uq6cKnDJWPf8LCroQIe3DSjhO1
/TuAMZo6zOrl2J1XTJJXGsrZp6znnC+zP2mCsyBA7NgqN7AHb+MeZHHak/rtIlCh
21IUqnPZvQv4ZoxC/nmKfD1GZbwzXhI6BS3/6k0H9X9R5BFhZRHRI5sPJQVNh3Ki
n9NRINDPcfMbEADXSC8k3kjU8/EpEJjSo87lbPdX4y6yP9SCp13CkhFU0TmQJoJ4
LqrZqa9t8TSQQIJba/sw68gYhEdT0tfAirXq5yzMTF2yQ0JLyvwK2hTkrw8+YuMW
/vQlQbyLBS5T7FJJRvMgEKF+6SR9JQcfq0Mem2qnzRZIGsufO0nU2152LndPQ96l
cepHWMx4Nq0Kw8sO/453F1TVGMJlZwGewk7CWu1oMQ1QOljN6mm5zfF6Qn5q4/uI
AYE08/tH1GhgvZvhmg9CqoB2YBft+EFDYDM6meGZqny/ZcornMRLVclx+TsB2dzc
0HUo+xv+jgvscF7SCI0JtLaHJrjR+3ZVGF5dVTa2b8xbd5iZGE0ajDHH6s67bsQs
HGVEyLcnlG0mjxEmjBeTd/0uIF5IDseaLPbGsfNUa8GSvE7OnVeoOM9sHQ5kRJvJ
A1EVRh/1pWLYdyRz/bldRf+Ns4Mk+b45dkCppmOw+g/iIqT1jQm9iObiFGhxBKtp
OpMtAwdMEJWPj2lz+qbk22OJi0OAfQuUS4z2d4u+AyckwkF4JnaNQfyJPyyllr7w
O279F58U1PMC895P7Tj/72snkAbLW/mVrEXuOW7+53AZmciMHAvMfUKX0L1lPisP
vZ5sFnunKAdRmTcWahvg9hPmSy7vADcWSPx5AHl+twTtnB+Shog1naZibvVT25hf
ez7POl1KU/YWmFN8oMWSLpOyXitEcST6c+zZMEZPyDxvabDlCjCbrKXsEo9yPylQ
aj34X7Em5QyS+hcVd4lsxbuBsvTHOXVaXvVXEfAlNmO/wn1sBjB/FPgwdsJteq1t
4to/neKSj9L4BrVF8yrHSrISpIKT4EnGfPBQmpRpgeFfu4d3zRv0/sYhcWFKHv+Y
UwRxykFFuqM4vC8BWfVP1eECK8wzPMBzsl5ryvOsAzfyIrZ+lMkpRHH70hKVMWtT
yLmb39bC+UHek5uBqUSvO8lLjQbgLOYlZrL1NXBfY0w9LjbndxibkO0lZ+xNX7l8
s/DOJfjfnV9UR8LoiZ3NhM8BnT3r+I3A2QkNaagwTciriMjTqZV1vq7s3OfLjAad
Hlex5bDfvna3+66Qv8PhjFUcNu1jZHrlyrX9wktfYW25giRR0SVNk4NxL5BunKVr
93o7Uxs8XSmIvyn480RN0dLJPGSXnhgUc59zEgAL3y20+b+0x53Fk+BA7YgAktKL
6uqc/aX9PIimcN5rKk2US2Q8NTK5dM9UkSktW1tzj4gR9v2i4XLH/2JbTuU/HN9U
asGUDf/e9za0LE8FhbvY9jcu29zeTWDBBSnaITmnC1I3XCUZU5ZjS7cg2iMRZTyt
5v2OQATkG99lh3Cq4QtRMFmuE2G/3HH1mWhvJ84WZ9qp2Yj7Xky33RJqNjubewr+
WOmUBMCEZtJF4s3fOTERcIC6+dr2Gd8MZc8WCNDy28z/dPbeZgDllNB+lrJfRmdt
HPvI5snqn7BKOUqw+ZQWzxNDA6Sz3VqOifuImmIoppCYU84RmoHOwkVYm0lNHt9T
qid2IQ6ypdtJxGC6pm6tI+qXYSvifgMC2WbIbw/V77j7HiQ6Cm1A9ffVQWTACC0n
9/leJU1EP6ylPrGMH6yaoC39lK9b1Q56ahiawwV2coOVCWg3+WcmN5qJAbGic/HI
r0v8YM60VuhxaZcgoWCGWWzDpUWgXn2bzh4nYMaoOx/MRu4UluvJd50qKKRYvh8j
Znn62ht3jXZY9scOSNVN3bclTWbfOz8trB17qbIzLdO45qqj9SRfRrnRZbqxIAyz
3kXCNcgTezQ845VPK8mu/oRo2MAE4XeJpZFuVeEp/7o+NUlnVdTqIVBB2rHJfzm4
ByjQ5UcqgGtHoFyDv1pf3j4PxOzwKusUYyxwB4zWlBiF/t12/Q9Lpv/5WxxUhr06
L9lmLNNln3z4hkfw1OP/tV5LoR1dGcCQ1XuXmjCkk0Ylx0YlekBAEhr1s+f/J/aS
VVP1dXiR7GG4TNoZOBBormcfCoPeTo6UTRC2gDkJMVhVxPIzkExRHOyPR1OiMhkU
PjwOwQgcYrVtUjt4mcD2P270NZJcq23KeUhPs/nKpn/iFmkymhi5PMKWzaPmrYss
WtQerUMu+49XqwAT3gFcilU1H718i2anEs5AuBRnGgOKTpzJbU8eAWw3RPU7ZB3O
mXYtutbYZQic2W3QPejhj8NKnFq7PU0M5AOtcAhIqwNAQvVQljfkw/Z3YfI0CxVd
4smn5p5I+Fy9l7JWrGoF1StEoErlTeONwZKyMcv9C2pQAOqm2L1QyYt8nBb0wJKk
9kSjSlwfnhUbNYXUivelPlq80zMcgVYfHLtzXTPMFXdcC2wUFblZJAAaroIb2Bex
4Nb/XYM82RnTbBzq/M8wpaFq8kSs/7hP4Fx/4StQjSu+SCe5mihom8l2SkiVXhlX
mtbGj/OgqWlAcJeISYX2aWEmPzPNG/m2VPMBWQPRlXjebawYpB2mH4g2m0Ecsd6s
cVMIo/GQ9w9L4qR9K84hkrfGi9zs/NTcAI+1VhCa9BaMnj5NcNp8fgw6e8+LZ6qc
Ghw60Z0cPmhNRwel1UuBw7ne+C3m1X3tkS5p1FRCHt/ABrjt/br+JB/BUHuGDcUC
fTqAK4HM/d5hAO0RFyc5COS9raSRpaI11MJcKlSb68IeBz0pUGYhS2u/vq1hiL51
p9kEimHmsAIcMhRcwxOZTykiyJDY8Jic7b64RsiKo9rA0Mx1bdgp7PvX8OgR0Pb4
7oqQF2vAyuD3sOyLJnEM8Eq+7y4VQZpUk8op71hXfsjQYt2z9EaafQlQrlv6Ke4e
ITKh45lVC5tecTFjWAcPvtpVSA4GqLSH05XQJNz0vnPKHpDX8fJHxJOJsJ33fzUI
bw7D4BSUMSHdW8hwdLMW+TspOlSkeUmyjr3hQxStEUBF3ZPT5HYFkYHLEcnTixXi
KkWXQUBnbwILGgCkt6g4Qsp8yp8LcXmsMogSKkmycGPy3iNekeXO555RvPq4rv/P
puyjYfQp5kBLkC7o2mRWSfutLqoUlP3tZmDf4ylLIsBSl+86WUmNsIYsGwMQkwaK
0dLjcwVvr/cY2BUBpDQlKAFVaLt8oRN9kprsUbL5WTlBolpEPEaLWrzffmyEH6xn
qWaKoYA+U1R9Za3uwUWxNtv1HrOUUsrwz2OYuJedxIP7dz3LLXfzRruunfoTR1pj
o32C1LRus/EeWtq7r6PfVlMdoH+AfA2prJJMBIbVfXsyX4mtQHdyBGgkv3VMrVw6
/OZihaGHv0AMiiul5fzSZPtEc3v9YOXiyPcHnnfChWQuZOG2A0MXO2rXGPt08F80
ZfqI/1fWOUbtWRmszMZgJosjYOYIz5qDZ3AymLyomVCygF+FyNq53x4qk6lwEv0F
QE8K/iZWcKFG4F7Mfoen6q9V1jRhqGPDntfoi6XinHlRtcXHoU7LXTyJ3vai3QJf
KwXntudywVxvCfb74gspEuJy4BNkJtK0UTKU43PxSFCjwbs+A8MgIajO/beDcU1l
4f5DXl2ZCmF3gTw9w8JjDkuSfXQbEcr0j9IGiuBcCo1xkQM2bnS3+7TzfGZakQh7
BrXUiKmmy4+Ow38L4avif6EXOtzr1t5tZoV/mFGgSZmrwVn8iyC89xRr4qLb128O
N4i+WpOUdmrnIzOJFShCH05QQfHkL0AWUHTQ5xWllcNYLg/VnPB8WTyQhQ5aQ4ov
I9B4rAsGv+CykCknroq5ldOCjXNC9QTvvxHs1I07tVGbLp+guCnMCTDA2qz2h/Xm
E/NudmbBlIgUo4aB8HT60z7NmUQ6SYvmWLWlFz/rXe6Ky7gNfWrrIatQCYxrwGHc
b9DWH2TVWZKEXspSjgNZsmB8ujAFSo3pTyqaC63NPDbhzafRQZ/KAP7xXrsob8cq
C2HSoTpxyGD6F3onEotV32djXxlsD+SPkTUI+JyUYc0R7ItrkYbvhnYUtzTbxlef
vjH0HNuB1ptf6V+v7qBKp+lH9dO7FFvazF5Zb9/kRXk91rbKIWLBiGv2KrqhG+yz
i11tvKbGCL2KLIBHBB3cmCi0F2pxWN8xKbJKG5SCfolk2WEte9509iRcKxFJZMXJ
gEQPa8Pfb0PbFwFFy/VauVMgOX5+kyzcDs4Rdua6ITAkmjtVh/au09WZ5EjLnrbd
5a14CWq9wnmpPesHYk0ak2SCxeTcPDnHwnX4nQmvrpR80EkrkxT7YpRbZrqx2dpl
hKms+PHe7CBOLrneYa3lpG5k2ijz3/HTOebCWoUR7o7nRSQBsyk+yt289Itcnbmg
NKE5WlL8vPrG41MQ2rBPAaI69ZLcPB/emj0kP9/WZ4spbZHDUc3t2uuD+mwMTHIt
wJxBj4Foggr3bljrlNx2RleNx3SJpikcvlteuml9nmbzeqpRKm43RLpCQOpmOMvZ
zqLI6MflAGdB5yB5mGSJWMdPJCAt28lekJy1+JeIL/A=
`protect END_PROTECTED
