`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FB8YncpFRCr5ism5wiXOeVQttxMj+8s74jjYxSlw+ex38KP1MpgvMM+HYfjA/lk4
UtmSPp2jQ9b3xxhYtjgORyPUHsKrEd21/3iLfPzxO+ixPCGUvpn1WQ3x2ZAxJyHO
xzlLCJbTwogL4yatZdYddQvnjvzj3u+Q5gCB0PTpMXe+2vCJY0OadI1QoiKFIPa0
oCMt7HImo/RBzesoJHD3Mq0S/ZdAQiLA/PavisVMETZ4trNV2uQA2cjALQKRGB/6
TMJ/X3Xju6WNvHI8I+AZdtlBSXXNZBco4SJ8hphRKDFOiw1Kl4HuOZzDWXPgzegp
79iLLRkx1IHmees0rxqzc6rrqQa3BJ4NyGZK/ojtger7BfRfOfYEj5n9wk4044Er
Fij+8Rl3dVn9b9lVSGErOdjgj1RV8P2D7viK3KFDVUZVru9mxxvXMqozbYmpuvEe
HHw4ZNfHYsUAtDo3U9CWtq0o11TeWAem7g4pGtVtz0z7/tJ4N5Uztg1fGaUo0xW5
Ba2g4IvB/4hVsCSJt6+czzZ3hQj2BxqjbfICaAEG3L5gWiTu50KGuN9aKLRCoyni
zT0vyvy51vuO3okJl9M4is1pvlizLADBfZ5w3DJGKahHkfOHjx0y9bxsfCpuRJQP
y6raUaPv3cI/Wl7W6df5h9zJxqmNcjHRrgyH5Kmj+jyjJxDfMoSesEEJXp7Cs1Oj
`protect END_PROTECTED
