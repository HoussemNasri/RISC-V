`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+hwPqN6m06YgvhXdHLVn7pkIzPJlNO+RVm/YZ9cBuceLmoEplnIMRPcYzTlvBhik
RuI5PokO7/3i2QXKJxcm2uapNn2EQeLkVvsrpL9gEHnX1Qxw1JXad3CvCQXOC8Qf
3FQXzfJbmTka1wPaqkRr+tuBKL5ABCRhlSkxYGTzcVAVo1BzSz2Qz0gLNC83CUz8
caO/kFB66r0ETqgyfcl2ilFx1EM1b5hi/wueqe7R5pDIkw41xeNkHtrhosrW7aUm
1XQrIYi93YS13iVe8a0JiOcp4XswBWpRzfoUqgrSAofQgeCEvWF82XMZCsOFH+7a
IPu/tgHNykGsTSJXAjIMw4xVLYaazYnq6qU/JcZZ0BhPBHfRra+56nxIc+ZDZLUa
5rdnNZustHOOJfBMUI1jxA2kLPW+z404LIEJ8rvdZHJ72RvmlziNuQLtcbgWTLgQ
AElqcFHhBtvdIriV+zm1DL+G+D3RuMx+l3SgxM1J+Wk/2j/hVSKnBsC4qzBOpwNJ
v2MNSLfKT2WWOMbUYBfagKOZVHQbtdVYINJSj1zkGk0xOccB7Jf538van/ERv/Sa
8i4Ph8tq7/TiweNTqNlM/SimgT4qNFb8dOd1x2yg0gPqfrfX5GjODF/n6oQYYqdO
z/vSm1aVwUFyl5ctHhyUB1553+zWQdn7GJaY8Dkvw680pZ+hrHLvdRMrjN4fPc6V
Djo2m1Ixx3Pph8+M7SE/oR2XUdCqDrQORcP40u7X9Wwl4HBFgQLVLoEZFIZMmuw9
1yP930YXbLjFU7V4hi1LFZ5Vfa4LxW7rjTIiEpZU6BkaYAVqSPAQM7jJB4WABz2y
PT3kmob9O7hK8qJZAFbO5W2vHyI+qwFspVddJl/htM2N4KS/ayJXLkaDYNrIOXvz
AthJi0koeiole3shgjRV9D7cCEtg82nKApHjKdzsJbDNcdK+8ZLCuVSn9zT9o128
OeGoEcX5jV6URIgqt1oVMtsOZ/NX0tqbKO2F+c9b/vqsH0oaIxp0voM6DyiJtMVF
H9jHvOSjVuP1sjvwAUNEYU+6nKqUe8OzSs36ET488FWj44nq1wuSZua6zQJG1b55
HYHPYaawrLtHbrToBZASK+t63LmTFEWFuNgLEaO8T8HmEdAwn740PCFuwsFk7Y/r
MbXyaKatP+5+nku/OirYUsaJb09U0GuOwj7R+6GVx0s31aT+mwizebfo7fFnM8d8
MfhiP02OVPLwBlaV+Vr6fThwl2g6VtCgSRBkY4D2Ef0K3er0qH67nCjxUPDYmqLS
PbG+PzUCn5paCON22QY53nBkWwgoqDDuoOiCeIU6Avfpb6cyg25BoPQzmPJ8uSzr
5vBukV2k/SMNcPcCY5LKOwN0vuc7WvvqNMKCjxDoGWt2St8pL2nbsATdEMNpk6y6
N1Q2SyCn/Y8+XHIFh80hvc5FTgeTMtjoKMIpHsA0T5C2plcqaKIfgSY1+PeQEEpo
9tRZ6rwpwqMG32zdNnQEuqROOBwajkNL3qW17MYDdmCAX1J/u8VLRuUR+3hjMQ9h
0DYMgiUFrDpCmlXvwV/bIg==
`protect END_PROTECTED
