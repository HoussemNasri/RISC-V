`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NzRDyHZrMDQR64EXJOzMx3grkr0WRC7Xw4uUMKxbUpekn6OtPEuECj6zqRZkkog0
MkIZdCZMMrmZsWdJdyY4/lhsCtILpgX97NOAzGCQXweA6SZWQ8MTCsj5A1rtptVh
6HdGyjaw0o7t7dyKzF68d9f1sVLMv6do6aDSyvQ1ss1TVX7rDQk1a4VLUfeekh7L
WDu8w25hS13hWjiwaX9SaquYx1oavULoFxIK6LPMm8RdzviEdHFKMk3stxRmYYFN
smIjzF3ffWXy+4FN8mAZBF/e/Yu2CUvtOeL74QL0gxXOKM/wogBGRjxT2tTyUtEq
dVPTHoPAZNezqIpTmFKmLkmmNUG66V3ZfKYtpuDa8ABfLFhSBIQlmSjSxF3tEQJw
MVRNrzR8ypx3wsHOhZXjfuhgGHbbP6cLDUxdX/9aJ59A8wkKUiOjC+4w24b/nddi
4KGjwxu11SmtywHm/zNIVcIrR1QE7FfJg2e4ohX3vdLrdeRUJskflIw14WRU7S+9
E6uckFARy38b19gecQeolkV+g2Ow9AGkvhY5MUIbl3iYrszIeXjxyK6NZmk35jw5
CxczmPS8fzRXAUuctuopESns2eMqT4eBmu7/tTW8j/luhaLqjjYVbW5xOT4ZqQHZ
lXrIWv2NwZnm+YOKD1tsXvRiMmliRWYbb/HiI+wreFVIirQy9piRlqK1MgTrKf/c
fsOnGuQcEKn9mMuVggdANd5cZM//8ad5HoyImf06B+JBi5oktMH8Qb0tNCmsAdm4
jDjXQAE/XZMw4ygFZk/r733/+y8CJ6QRHZJrFoyWv3Q1AtJ74zLgH9Ueys6UmTli
3Mclccl34nL2frE5gGx3ypY77o4MrNqGgP7TPPvv/MFaUjdlnp1Ud3jEhYn1EX1K
XvyC2YboMHA777Y2QiVk/ZcI0G1dZYbczYA2p0YEV+XlzLEkYf7Y3JkysZSDbGt7
UCOotbAutP2xx4pLYIOXch5K4Q+La0XHDzNPd9K5T4ugQaTfgeaNBadGkspI0q8W
GBg8aH88MpHtoMCexPC++6Xxta/4Rput3NPKA0wTdvlsY14BnUr6Uqc0zJKupYw6
YpB7OqqsJ7Ayw2mHuAw507tbY6mlNt+SFgY5ksdOPJWMqtVqqkN0trwb9avUPIQt
CRq3Y868SPE9SEcjoXD+6NzZetDAke27PG4iiBNtslQXd7DIl2jQkNI+c1WUgdTB
XwRx12QFt+MraEZS8su610zen8La6mPVn7DIJw8udGY+tlqxtJSBTtrTIzQkzOjM
jSGgx+QoiQN2G90O8Wis1tmBmOtCsNVRgQoBETzGGK9z0+AZGVi56crD3RcxQcfl
Z8vxXG/w1IbBWg8VY8hDJthdHncfzMcSYyrXtiJgjZ5NRJUBgVzYmy2IH8MfO/zP
IHi+6RIQCeQAEDOWpfX8r/Lu0cffPlPbhLLDKt+gIrUF/4s7A/1txlEdtIBLSVOo
Zdd3BXjmEDMUwzE/THJdRxQruP8zfcwvUeeiFHWCC2twalZ4Yu/Nwp34c4qhhJpd
9khL7cbaS2W8hJ6tmRTd+o/lv2h5JeY7YWesAM6qM35UD4+nJbLKTmM7qAKyDn7m
BA482x7Z/ZcoihdaXlsuPefi6uMJOdOJg3JEPysqR+6Ho/M/NLrRpl8COiq/gHN5
OQllToxS/hJJjM4wbQNlgWOBypShvi1BuskD948GCni6Z5jWYp8Qq8fH3H3XN9hk
hxwIYu+XC9tlN5RhGgVDHGZj5WIbZGlYzVouowpNTQt23aERn+CNx2cERzWybm83
N0p0XgNaJ2MvJrz/b7mt/dI2MTXXBqoAVmEX88AG/htwxSI3qXeuPXxUap5hAdmL
N4mEU4e0vUH0Hyvqgbu/FmBDoFjjj5daYLajWJIPV5YYjhzgeoBLD4SkmJKAQMtS
5NOxC2dQntjNcoxVbz/mp3vNxDD3szb2RZdMUhNZwLsNb+epfv0jmYxkKqv1cKJg
CeH8g6k5ldGllRixXyU4EC/MtvAt9Bv+G4NdNK9Fk/L4M3eGSxdH8X3lmWsNAu0e
rMCt9jnJ5d1aAFc0rGjun8PiyENjztIJx+G+tZ4bZjFrEmWz90sqE1v+aOep1NCo
F2EAXxOui1+Qbn0+oIVV/eIKRhg+OjrAxbZReg04TMl4qMY/qgJSUpahwhUhd2DU
t5c51bSEIgGEjO3OOSD7Ya/jEWwXVJAGXchorm0kBhDa5hJHKqFze9d/xalPcyHM
652lDUs57lkPsHNLW1yd+FDeBdOAcSyARWYedHyWz4BJf0MbGyZv5LPy9a17mf+6
8GuH7faZUeccmmU5OX9VYxpxEWVduriNF8Yhf2mfbfjXqLfJnHfFFkPyHXagL+ro
lI035ol8Q9IEsybviaX4Og==
`protect END_PROTECTED
