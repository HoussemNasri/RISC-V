`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2eqtVIKxP4DXHEz/NQYDMkoAArk6HcchoGxvwVhranNm9eVZPSNzrWnRkTiQ/z2
7ZtnGYY76bsU9zgSDhcgQ/HCNymdIOJcLdYhMJ+rma2yQe4JNj/P0uBHKAfeNopW
c/L+1c0LdrShgqD9stOb59Av4L73HQcyerpnxKNud8UZWVr9/kglhLYzKR+lV+wn
z93ytRMkkoDslBLX5tm2dDWoVNQmTVsFu2db/o9l85VLkM3F5CAo35q6YfDjhBbA
TaqizT8M5SXZ5T3woXaXfHg6Cyt2Y7Kk6uGRcGVnVWMt/GxVv5s+Y6dihCrPICCe
alD/oG1Oay+zmiMB9yCS0wpm7Jhh0zxb/o0DJ03qZTTXi0pfARLiY6lBT3T4RFF4
GZ0eXuEBOFz1SBRlR5fGGP4LtxKHovf3e9bGUghkyimakV0taC/YpP4KHIgUESMv
lY8B3tpmSp70sp19YULyV1Jvga/40K+XhLqip1L7f2hyfIn3d1mokrfWS1GMtgWI
1cPmFmj5nhnMJgHvAr3pnLeumJPgCzT/yligQF2xFNaJR8ZBSDypPb21iYnwWBJe
o1qVkmrH/QYHt6r1slOU2PPuJRSyBh9cCJbLxylK/bxt78QqCrNAijY1igjfQ0Jh
z3W6tgU1LVK6MXXrbMgOdZDo1eOtg3qg675fpor3QKm6WSSG3QKuoP4NRIftwh05
Ydc/fHpF+uuZS5E9IG+V3nyRKrLtb5lIiFa/3Jokx5fA3cVr1hnRF0o2k8VvXNEn
plOFE9AzdeCgmLedhSG6Hz5QiS8FFvBDykymR7DXrBtSA8Rrep/eGCmLqM9VMXkz
dqUexPtM2OIyvUcyzd8zYvKIlWxJww3CrubG5h/4t1PxaOvfnZDLuPZPZporBQQX
ME0wVHh20H2ygXk9U6U2jwtmvp+habVaQCUJI0uAH5J5ToA1gYI0QUGnrTc0N2jA
elT95l0B8FQxm13tXClzWvyKoI9xE4DnwjpfvPRFf6F2N2x5s5wF2hU9sxwKKiQt
CsQkCsDMparUW1a92OTW20TVV5Xlv8zaNHpOkvrdFQYbVoFUvYxoQAfbMmRPDtEF
kOlxG3qB9kfCBeuZHFd57aOnCZDXLd0dezJAwlULHl+A46hhVrDlbPyp8jEGPQhx
ggAJ7lcB4+NzJV7WYpbGW7JsF6UbgkMI4/OHdTrK8kml0BN0MpLAaW3iDvF80ZvK
3KCILNwyfSOECUOSH4JI3XBLEsfTT9QMYYYt/dNILHmwMSAYPjeT7AnA7UlYtbPQ
xnDNlO8B1BAt398Uw2gWJa0/FEQlTSSmCN+TWSm6gKP8GXCOXbSlf1z0EQ4agKw/
VMwok/NYGCFihlW3R2cwR+pW7uSA1GQco5sCmD2wn00HE9cv5CdOXNODJKySTatK
z2uNn8ZZX5MfPbszjwzassyFvhAyvs68gkN/iGragPCTW6VPODo13lpzPpYTFB94
HVb3yDYFbzSPM1dDUL8/hpdli1isUL3ZKVFO7Bv4srRhGy+s1QoqkJL8SVmxmla4
d7VFjCc2c05+8fdw2/K6FOPVjZaIHDWCspS051e5TYUQ7NCcZY2vUnAn4jkYNuoN
Wsr8xFcWdFKMGLpR9ViSgnrzjqivBAI6f+AG2CyutKdGCoM9Vs4R2IkCCgSYfYUo
0xTT8pljcSuVxws+4AnlTwoexjSOwbgzwjb6DMimVS7OdiQIq55m7Q0gr5yhhh2y
Tf5DxmXjBRGTl/hqc/fOukTFuFfCSnqW95UohBJKBGo6intSE6/4/4xfTO8yP0i4
vYMpC7XXCVJRD+rqQI7cnWyHvT2RD16BZ5BJL8FWL76Zh/7xzatJtu0XXzQfOgry
qiD0jestTNdRIIjs5vezyteNu6S6hBqUEjYimc6TumUs2WGATf2TFEuNMC0YX0Z4
PR8oPSMD2ngwnvl6u3Q0hOHfm7JXcYumQP26riqTvwoM3hdMoMf9MvOjPTxP1Qyf
b2KQoXSMAOkSJCNN0yJt0ZS8YUlu8ijL6Ofy8wmzuarDbKLo7dXFmxmKfE72mvhQ
4cNcNt50ByA2vjUgdWp5TDC6O5+ZtV+pQVVlFlMLko7HYWdzJdr8JXJSUB1nDyxy
H8RMecO9ae5IBCHOqxc2tbbMG96S3TZK5ew7bhuwzWQyhdluK89WW3xzgYS3j9WR
zEIAkjb4lji6G2lgmJk+sy7UUBWttfZDWawqBwJPq/CispjnWFFTY5O2Au7W+cju
rN/U5sFKlf6qUIH5MULktsRvsxsy7MYqUrF1JViAoo6hSs+eJMOtmo9bGNwGuaId
oSNq6K8YM4bTgt/8caI07INXtoH9OHhmA0hem+dDxvC7YpUFlmvkSmI0szV1XP13
FcFhyFPz0O0uLMpQn06BS6omx0Yx72uvCfQkvUJOiyoygy/KgcxBJsNCfUZ1O2Ac
qBrM3hSyUtbwGkVCL57zlgHd3yZoerSmm0WeMh2rCwtzvJWh3GrgZK5bcmqs662u
+F89z8SAEwKRaMXzHSKD/gHOWHUJXcVBpPAcbTMo6ang5kdYZ01oLomwzTA3TDl4
/t/RQEuvw2q62zICm8s636GkakCC5eWKEJfXqpNL4JPRDK1yJCkz9Xo4H4nxyxKl
83jMvTBofKzhMa/9M/+FAEQ58hYng0HXFgy0xE0Rb9AFgwt76qK+CtHB7tJkScvw
x9igsElUHF4XfS5YGxKs9dqz1IvLfZ+XjBeMnAYWl8QE9pmZJ+/NJHu776vdjN+c
Iw/4G8Qyey7ndPQ1OEjubOr9oGvMCKj7mtB31XTdygP8LGE/O5dOh2bgnc+e1NgE
4tQIic8D6G3idkOa9YCG07LtxriV2nqpHbhsvRCTiN+q+Ab3Vj0GcZJE52YT/EZl
VyoVQWMsO0kBsLAikaKvisaBYTEylcWLqEH9Nuj75BIKSCiNLC8IG0BZaECVNs0E
DwrOpUqEXyzc8M5yRWzQg66mlBRdI3NMLvh2bDz0vP2bwBerO2JutMFotBxd78VB
kigvGj9BMSYvKmDJA7F4Us5knkh8iJzwvt+WQoPVf7Nsl2gEz0l0LKXwDtW1RCzi
A9EJ22Bk7vNFX069vDTD+YyGGvOE/todFm5ErlA8h0PtJUo0n5LeQ+lKJUCdbIyh
QuZ4yqhsJesWGmaFSssCO6ixmxcEbxI/nPJr0yS5oi1lI1cUfYQRwukigF916+ZU
f8sDz197y4MMjS5TFKkA3Qun9CMfd9nK0pbjptdwbHBqD6PpkEZESovwd43p1cxY
2hB9WBzBFH0NGJm36Vjl7cqJeDASalCJiro06jxKai+RASQ3omHHtNJk0GdspoTW
yVfSG+C+9b2faOuJAB2H7S4sPQEbpJzj3ViA5tAx6a134i7CnS+iUt9Sa/+YLasg
68oxyn36CZCOFW3UaoBoPu2QclIlBXCD6DXRWiq42OeYw0gnxfAqyADaX1lallP5
rDTU7zCiVUAmYVFb6r3OKVhcHlLxk3tlE4/LsHDOmbd7P0JKU+p1JSjFVfpt9DaH
99/+tjDMxsN+gZYk/wnSAFIth1hUWyGh/wMHKfHx7n8HUDsN8JBCUw/G5A2zzHTK
GD2ufXgvC6BlFXUmmOCaBmxqyVyO1xgC/AnZ52/QWG6ptoLtPAB7Vxu0KLouCsmU
4garmzhZqpiV6ILKUj3ZhbM0EJDcpuES6NVQgr2xVPpElfGFyeCcgfSlODeppb80
VVetCWTDlSY2+tOc6pWLOnpG9pxltSzMEKNfVoGhg8z8inIY8LknvkRcsf8bU8sB
lzwVEKieXdLTz2mCNjFwojHtwQEkV2bd5rEB8DpjOD3oCL6hBErZ+DQtobNkqQZi
m+txO2NTTZQGyFEgam4OUqocgKAWh0J6gNWggTzXql4U2pd/jP4VzncoyG4cgkeX
jp7Mh7wfaePQ0V4nMmKOYV7RfRd+onNYn5finS9T8Xcin7vyL9pj5o8Qg2fXfAK0
drOGfFnf8RRMTgsYaUl9lyxC0bIBvMz+V0mjl9rAzN3F8lRhh9ghV12oPAi/aAnn
fT54oJoJ7037LoXTbQT588KXyAkbx+RJ+Aji8usf1w2i6Bmd3kF/ynNWJCQpjaPR
5HYzhMf+rzyl+Yqgzn76Ofblu6QGR2LoQ4p7AW7YRK0BKxNQA0/LjI0jnCUBaP1w
F8XYsICpF5o8ziK02+LJ5cP1uf3MuEe4dGIeVA5V8DGT+4VAkQ1CYJvVT5snNy1X
4nxAjeGgOSO2KF5zVIFl9tZzUBE3SeksPOA/ydAZ1nWxmBhUyYgPmYCr8T88o5Zm
koO9LfG4nn7/0P4j8Bi3ySO8FogekGUOZE6CCpaV2Fhhnh+rgZWviDSw0tLQ+8gS
qpbVtsdAZdqpnfjmqheCNBc3vLQvLt063XMyzsZ7MXB16VHWbXi35sghQPuw4wWS
k0pSUH0bWNN1JEXVBhs9sCnhq5XlCE4duCac4Mxlk5Msfmf8nAU9ac/q+idk+0Dl
aCXvWtiRoCzaCW7Se7lxzaz2fbIW0NHms5BFrBI3frzTgSB2KphbdeAJF9xW9vBk
PibZAywTKWnlXtuVGIUf9De+fgn9wNeozhbqugKtk4MLsDAJ3+Tl3OFp8Vfs+GwH
Ete9r5t87QIG7ruEDQH6mVaNy1nbm4X+pGT6tqVpktr7hK15k0A+mjt5v8zSmKJY
b6cNyu+frJ0z04Mr3Mkj+K7eH8qTBFBaFJeOCTP/X/75KSlOZWuQGGnShCkphDNa
l2sJLIJbXbDbLg0U7vc2JiLynZ6AM73nUplSdxTOX8t4lMvNIF8/iZ+kt2Laz4/I
4eA3AHRUw40/blkftSzNRameNv19b8BDVpb4P6aYrTMk+XJ5el8J6SktUv/nLzKh
PRVVOOaBroEINJVB0Wix78OEStTn1CQlozQ7uueUA/XgYJuyTfQ8HYstExtJ2+sG
6z/RBw3sFzMvyiTqVbPFsw/OSWJ4oLTqR2YRUsyalGXv8CvKBzjOBqlHXLdEGeAm
FfQKu9oVHdz+m5CkRj4KLt+T7V48/Zz1EnoxD8ZzJuoqjKrbW67URQQ3P9+zxPJ8
6pSUXzr8LgAPbsVS9hNbtienFCcnFQGO+FKTjtUj8DSp3OY/g4+wCfg2oaiOHzEu
NSmkBHYP4m5HSLm5pN4531QIaaeL4C1HzYk7igrR8H1bXDMWJMCTU/2wkTjoBDJ5
JoG/SaWBSbYVlcK7V4yBBx1FqibFB5X3OY/P614ZKPdl3mN4zM5pMtQJD81AOMYt
aYXunBuInO52jX/ZaiqLwsarGtMWDGFobKuyxAkXvPqZnfJayU3n4sq1rGVTtGT3
RteutPdbRYr5dP3QehOBTzASLGsPm5NqZ0GyQ1jK2FwGi88vMngBqShHIAe0S9rZ
tvj4flFPi1rBusd0PZO53IWzMrHsN29ti5MZbSSzbWgQ4Tmiu8abmapuCnXPr+Za
/2TLoDX02nsyY2oAVuixUCheGU14ztH31cT2L2yxMvVfday6sHK3wVjVn61TxGXu
8VERCjEOXJ3Zj5016yn4vWtbgnXqirvnZPMxTi5aquymqNjTAktlTMMLE4ORwHYz
rvIAEMYw2vgoXDUD8JZuXCqDRtZGaHyAr5/AYRK6UEobhW+BcvNMzst9mwF+LCSi
s8sIERLvTY6+yKBvot+UfPhleyG9/ORBXGKz7Oq8TNos+wd5umC3wkCN8HZ4Z2bC
OpRztN/+klkDFlgl7++PKA4/Vdx1XgQUwmfCjZr49sLVFeTNUFyPkCY+l09ZLjxY
hhXK7ug2E/DmbqhtbuXiM68Rc0OEuKl3yayyYtU3jII1mURTRfGATMmTRjTgm5aw
cvhQVITOYHf5eEwpiFv5T69OKxPHbwl8sj4X3yF2G4z0ssRW7p61/DAo9OoMTJ0c
Z88iD/2RG0nJi41F1fS+bhn7teS0f26JnYKyEdvei4uJGgAgOSSmh2kOTTYjcqNz
/+QgylbK/ebpORWwFakHIBg5LUNWwfXVpOZ5jZE+EPxhsPjkOWBMH2X6A2n4NhQl
/CDtx4crSQqNyKvRL+tmQge7BqlS5+N7LXiINeXRR5npf3cerA3/yjqQUaOEss/R
7w7p6SlAzI2dUz+GD7gxzHnklWn5HHCbnBs+Wud6NO6FYPCeaikHiWblQthc3n4f
ncTQOFWAcGfmKYsVqZBu2Oq33//0a6cEW+a0rkgXPaftcuKd8LBfXGrKQt5TShFv
rWOmHKO9CvG4KNRwZ2SlzIOacufpjGbhrk55f2uxSj2DLHSTahuQvVAxKe+6Iesz
VEX1OchPUduIwwXPCN3p8dtUUnMGThArO1ho9uQwGwDcb5dJ7zx6XgZQ75OTjZMM
e1YT221zGEHOrkza51dLaBq0WQiY9Y9BMTIc6d42FY9PpMSuJXDXKRnH188ewlrP
ewgh+x9jHA7+mMK141SFGAwQyPCJjTa2rcmCo6GA1og1OWujbg/yBclmEN9wAe+2
b15wTWPVTDm63jK4f2cz3EEeSTWlpdBlmbhmTmQcyS8HyswxlW9hOIfEml9YuRvw
SAL/Xr9+6IN1359s0aUqCY8iv5ONjPXwd2M0Ul9Yo5AWUs6hbz0kbqNDgghvJNdx
B9v6KpZHek/TfE/asqgsBOEnrZQe52oIDMO8ClHyELqz6MCjW5t9pd3apw4z5mKl
1x9y+uk3/o1ZyiWQ8LIXraHFAh48tt+1ua3AooV1z5vZ34trKq9NPXLwA4nUDSS/
DtcZ/pqu2r21PGngBoWiJRJvqcGnWqB56ZuucZJYvgXr00FJtc1ycbvKMAm79+vP
e1ysOMtIBZ7qmlerg9kcl+41UyXm5+1fyxPWc4I9Ej8W8l7HRSxYOL6ZYmo9226u
`protect END_PROTECTED
