`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5hpsrIT5bWqkQ4yq9xlXQGnofL4fi3x6K8g/mPBATu4o21dHUBOjn0HyX9FWB/Z5
byaaFb9CFLcPaWgvQwU/wMX7ARuKsPcIlN8w/nGRqDKj2C/TPL5H5Ho2Qef0q3p1
HbEs1VMIT58Y7mfICj5TenVCpdOR6J78d+9bqbdlQguDsDvH18M4ypuFTGZnc1Jj
xelH7QasmwvVrUmBn46rWTbLL9t4nasl8sIjNY3Cf+1v8c32O4hHfaOcvheK6UHq
Da7CAhZcoi/f0mJQg+i7YLLh6fwF11E72HrP0lm3rapu9yHJZQaCYyWZdKd0jXnc
0r6KGtMNwOcfKlCxCdtEqEEmI+G+28pmroNh3auh4NjVKVTU4ZQ/dLzkmqMCYfd1
Vo53q50W4mSC9cF8mQlI6IwF20U4J36aInTpQ4YzJlJLv47+duKIiSWCflP+XWjq
9bYUjDiAqdHhx0kTToSp7rCMbWx/1KuuahPI4tW9XKw8H69TSSooSOkv1WoPu2PS
am8PL7Y/cxJoorBTeJO+kInZ5mU4/HtbCC7jQi27ezdSbmFnKSgW8wMxBrPeJJ0+
Mxq9BrO30vDxwkNsw3XiMkUnG4zHPuOaRgGFlhg4Fq6lwRTEeK3UYPy2GmogKod3
W/+JEpb23Alrg5XAz3gUXJno1iqqg4a3QQZejQa0oCPf13E2yD5GBQk2JTBbEjfP
rT1hJ+QYPUkR2ssttPbBmof6x49ChjKPgLXAbM6MqUFJT61jCsC8As6lFiNFDoP6
xfC6NLx1aNWQxjmhjoLMSvHyPeluxEROqc/UEoNyq63r4WV83xrjbdTPaPR8JRhj
cHXWuEhTnx7EVpt00ehq7JytoJFj+HLbCLEGGujz3Jg1XvpTvWonSq5PbnyAC4Pi
3DfrZO3LA5qacQ6T1s2nttTaJWACmU5hF0/sln+maHkSjcwGYgEZ55lp44SkEnXI
5obutqFpjZkiingXKxQQ9jluafnoCkWvm9woLQdgHt3EWU63bXkYekeCUB8+EqIC
lULibn6QrWcZCoClNB35qjelix/fX9j5MXfIfhqOCrJEFHfGkv5E2mdlwp1M+Y3s
LJpLP3hPUx3kjHvoH4a3nE+AqI737t0pziufqmK4QHHjhu5U8tSvX5afWXbOOALw
iYjEdvQ+y70RK3m4rLJmUP5bgf3uFF3eK90weyja57J5lAaVCLiyS5Kngw2t8Koh
qnoUv/tijMJM40Q3+J+rN3KPou1NYLDYs9yh3NfY56QduzjvvowzyJCtiXuT0Tmf
0Y7mjQdpXBj6wciuASsKoZ2QpGm5w+xub8UkLFvJxfAli/JojWr3XPx6DCG95S2a
xyQqejEnrec6hLsGzWVwK+ESmVFXWBqcwpSwfMPGl0CU77fRVFJ9fNNo+jPdLQpL
hu0Poo1AXmqLB3VnE5UoEjpxps1jICw4Zzbjua9/E783+0cyd3NI4VpesYQm4QT7
1wG8M6H/tVQryzwwVa72m5mScp2UdnEvbdBjCvt1JQHy6cqszVw02i90Mp23liXh
K3YasjzDvqJCmaZxJvSh4/EZPPqG1nZKZD7Pb3wZ0zoYKyCVdgnEkpCllNi/I/kj
8iErM+6i6f8BA+MpEcDETasOl8oohIRwZSxdIqbpd1xJvoNcHzJIceJkVjHqpp+9
46bzFl3lwMoT6PcJX7DSx+Ftu/cJ1ACDjYuqGvCmNge6CML3UkpPrOIxoPLZvBKN
queAHsRx43+W+nGLWGeCHn0F+USCUbtQKaT6KDmKixkbtxzwqHR3p8TEZCOGFN88
F+joHtec7ZaGNZhghat6GJl1yGlVlut0lApvRf570D9FCMpsFoX/NlOZ6niKazKY
XNdNSDHkuXZD3G1K0dMY8osfdHroCwV8LwOcDXAmQbYYvTypNlRz7mPeE3WmhOZy
2jiuYTI+JrgFMqSBzuglO3QWfQXuAkjA8G88VUByZn/FPvKJH9seRPrTE7Yd7VnK
gZ7OG6Kilhvi+YW2cqRjLCKie9MFKuAkT4kTU1yb/zpI9XfMa0ByEs1Z4M5D0un0
UarWyzgtzPVyOV3qGCuHGmvZ5U3XQEBJML8c93AebUaz2nZnh8JYT461MhB7puqy
M0o614K194hm4spsjGEou9YVZedeuNzLmLDFBPzZ4mEkgsNBp/mTEqNwm7W8etyB
xJQF/ehjYtjHhIATE4hz509Jj/LiIqT+RrLmQ0bs+3haq/VmSz+LcC3Q67s9Pn7P
F0+I4GH6mjL/i3wO/aUqiCIstL/ualj30zRUBWRJk0xBnhM1cqm9sbK9yRoyOtGs
Ox32iazM3lcJlXwftCRVF+CYZ1/yAR21KS2DOkJpNgU/6h5KPlkzQqKHnuZP1SfQ
QXkwXJgoLlPIV8/GijBLQyIE3KVbkGUlpVDFxuRJlH7yDMxPk3xNocx0Xm0DKT+U
ZRSdLguPbwenKEFj7nkORjUiZeqZU1bGpZ+6AR2fID48A2f83a/D1A887mp4clQj
rC6UqiJrL8xUeYMXY4QV8RpJcNim771d5AvkjBkyBABXumNzMd2GZy3EO1GXEOpn
i/eU/SZk3jYBGQjvzlEJu9OAkJ2dW3hR6xGEfbIeWRmn7tmnIK3DybmCXjRCFZ0Z
H01Ws38Se9FfuEzcbPqW43OskDPC2YJjHnhULIr0NgDLDSvWKXd+esOE4Xp+WDeh
SCMdCb08g4kO7wxQQdPae9RGG3n43P70z8ra4bR5LA1v9Rom9XTaBdNGlh7U3cMf
OCmKNV2ukKQmYSizBujJcOmzLqbylRGAi2pLCWRNcB/MRMSXLifdFmf/xzxF9GuO
i2l5344JTYznRhsz3eWCmckoW/ul2kecatEk3OKvG+m4Lmbf+Sq+m17h2CtOT0aU
bGfwRX3WeRvQBol4hoo3/KPDwKp/g0KZkdp2RGKtkERSDX1gbXZ8BYj04BNAQtUp
07t6mjfuTD57Xo/OUIOrUX1L86aIVhKP6jyPXhQS/t+5PHg96uoZpgL5ICbRybni
wDUdqTG5xXKlytKFSa162u1uUKc8b2QefjfdzZqmQTlQQlBoJkv1CM3QNwr0hbBT
jHDLAWAYtvFVAyrg/d53tg6c4zOfaOlq4SzFr2PAo4OQ06cu2svieFxDt3y/1eQC
VxJ+wdhEL3udUVqptnk9nA+MyDGgTdynXBte5unDK6NtgQm23fKmPOullXXNJ2oV
/eSd6wnGZMJYtI/HpMDDCxv48Y6bvnURyCu2jaXAGQDxQu+qrjRDBUJVWrLW0TCX
izGCYT8W9S/lxPhUiP4u92Lw+6pXHt4d2DzJMRruJnJOi/4vA5q+rgYFrlUduFKH
4oB17stDluoV3QlMPSjKufglviWb7tvowgumDT13Kf/NCzsjuoI8qUgx2wQGVeKr
0973H8KvT1WWQJAjWJF1z37wS8LaejWdzBQ9DBUUgrX9GjY+VfKMQF56+mMK7Jnq
C+O/xPkSpbE2vx1JFFCx356hUgX0lN0D2dCWdM/O526QFzKTNmjXmoTb1OZkfy7r
V20S0VZHJnOgZ1QQfMY5/bkXwrwPaKZUymnLXAezoKhzJG0dSxEKcqwbiCG1E+Mm
X19V4WxFD80tF+pCOjz+xaPvI476h6MU6qpp/y8C052ZIH7hxM+1bK5DguNaSB6j
ZUD1C3MF3enFILDGVoHloc6HUiO9aO1JdgUN5MgxZ/7OaJpywWreNqRdZsC5E1Z8
OY48AXQNZVMnOvELQF3J9Crtb79C8+D2X9b33nVR63BNnUIq/kq+fJSe9LDz1kmx
xChfdYFct9FZX+TvearRGdjC78x6TVIsChikZgFl4EoDBzumCTbN0MZf+1Dv+DDz
F4oXIz05Pf1uPN8O/vIRvTDn2vQzPHuH3Sats39+0LYr2cR/6r82pqj0mpHO61T2
QBBGgMqR45fbGFxv5Fnf1NS1j4NqtxJZvqCZV3+SC9KUKiormOfSaqg9SH/m7jZK
SNMqKl9954/sM39OVInrOVqKUNpcLbKMcsk+d7ad082FeBQhk5sNxKDeWDqFySuh
5GnhnEjLsUDD8y2mHXQVFwN17hhJnIQGsQPGd7za7cWZFEDw4ByZtRCOtCgX0DTw
QlL7w+WuL+Ee+1uKHSIXAIAWBtv1MJOgQvkx+lU9jal/qsmYPjiHfQi6RHXDAOGQ
WgxLGK7cIzsStdeUXdzEhkDjWC/RWcOnUiLG+BwiKtNTQJhuScc8WE4+zlRbhQXb
5fkSOH4dr5QiQfmTgygIPpXfDx8C9kTYmZctDlb4Xnrv1fKB7J9PF8sUS+u1PgGB
GzfhNp5m6gQjf/ajDUztuTaAIHm5M524YUv32tvNJ6mVLqipyK09Ybrb1ddmw1Qw
1XbKV94jfSlOtRjUhtKqfcOwOiBZWGNNMNe6Ve8if0w0cUilxFJatCYp7n3VdpDA
YTzJygWda15MmcS08WW/+oOj3LXtWVVOwFiX3Pvqyo/N0zZzvWrpIRrBqo7Y5Lnz
abcdZVGSdWq4Sf9jnkCs4p9ait5j+ZAKMQ5GfHcPLhuRNKvVB4qYPJWpeV7iC31P
yPfHyCTPLnb7c8AVXCIJ+ZvS5oKWw/clxRDfU4Sn09of4JPiYS4siYmNsLghWH3T
+wvYLJDInvddtyHF+w0DEFiAtG6VttyM1yAQMCilcR715MaQJo/7TgXsrbOBx9GX
NdKclFxgaUutCgf4x8mBep9dUNUWgOi7jgbalhuQHH0KB5mZLaAENiwL5THk6q+y
B9c2EmZ7mt9VrDAsmlxC9RuRP0EZE7oaTj2MD0EvlDh6movFi+Pcxy5Ea3LUWBNM
g6SpOKEueiv0CTS6nVvi1POV/lUf0t0LznqaAYvg1C7yPpHWVMv4gSurMtrE7jhQ
qQ8cDxUDZ1unsLJ3u1BzqIKT1M6z8+YytsmxL2dXTkhX/yvpbTyjPe5Py6nLOUN8
rAEZzgqYOi/7OIC1zN7jsvXAfC29bk0ObfPrPqKWqEIyK4UFeE7aI03adBwgxbek
f70oAIJIQhzxAbz/4/mkm/2BI0odpHPRSuhKoWleMF8IY+5eVjdhaDL54xt43slp
MmyKl0ncPdamEprPzkr1ksGSahQPHXy9laxuwRtR8SOtipvhSgHv5uvkMw6e+Dmn
YvKVpa+DcRvKK1hTvTuoVeh3/BKua6bcvmRx8TOECXowMap56tNmb4mzgt2LCQtX
MAVSoIyi6f2qujpHWbSTdL8qk/rFBLrr7tRanugZ4wl7E4M6Pg8qyNJaSPT5sh/T
L2z7B35DGVYFbpbebYqu3GZ5xBjkDoeiVgBLuBT5OBiAgSekZlt3MZPIVNYBsgGu
+g38E1d3uN9SskZEJYDdg16a7u4+qGa85TkgSozjf/phuvrEXR0mz0MP/krXIn8n
CrEi9xKSslGVCD/1bQtFTSmUoJs60tp1Rzh1C6kTw4p87wRYNz7izvr3upLtomJQ
LBuow80htTH+MdIuGRwhCrV9CnQ/uRYNS433cHwXzqwV9VErvqg6B1RQVmMwxeit
W00Fpt9MAqfQIIChyXE4ZF8WF3Ri6k6+a/xQsjIPJii2tefxVTSEjOz8apFcxv3I
SK1+ziFg2BtrPgKgFH4uRXVtgU5NIbiAYlBOAQGjdWteEzQ/kQKdHQhmGvoQmnbW
qMba+IewRT8g0E3gRhUQ0hggPcQwDUG2FyVSwXNzJJXAAxBMJVIguuSjYhJQdyqm
0DwIQIO2BYLtH83m/2XoXOSttGs/tG9DCQh0jlPsKANXEAcqLTbhkL9Ax5/HIboi
U0n0U4eZjN8Y6Ff40R/Q5iTzWMG5xNVUqRwi+CtSPJMEe4og7f5YJxFCn7EiFvn4
5HL/3zoyE0BZYbi8qniUkA3JnWLqqcWzIZU5L8ebCQVnVRDL9BcUOlomwcpHV9Hx
kjxZqWpPbayzNcbYogRdpo2xjLQZZ1uWKGMvpXb5hCBhuATiQSUGd3RXBYC15bw2
K4hHb4O7TSwYmcl4JlIjsYAvA4nFsKi6gD+bdbREnCd8EU4XyU7KTAaeJpM8a3Hv
k+wJhPh5gMHA4ux2TXdoxKd0nvXG7mQx61zNd0hp8OAnlBHwuvyMvcCALiI+7IKF
hu7ScoDx5SdIYKMhPxdY/SVlLA5t1Wy99uTkvKfHCjc6sZn2Q0C5aCpKBG+HwSAP
5/DgUly1wrz7nXym5meAWwlUpcw7cuZjGUxUG/P+8d0q1eN0XgXXEPU/CAqOD0wn
RoT623YQCENOFtWSxLFoubpUNSrDZwZ0aZXJZrhLDZ2FmY8H4h/4fveIULVF6WYv
NXDDVlosY8WUgPMmkWfbo/iz1off0A5BiULNIA5MYkUGKk/XSlloEtax67U10/ss
PktX2j8qtWSqxuSrQpjFVh5akDEC2WjgUTQJiEeM298mX0YZtUh4g2xV9IN1c9z/
aVIG10tyEid8tHlnHqsmJ7kI3jJNUmJM7etlRYNo/wUlLz88mgW/BHrE+hU3mUXP
s+PMC07Jg1HXlyLECY1i2ouVqm6sZ/7bu1vEyT7bRqbj1LYRX2L6FccUc9dYJIsS
cVMdjhj16svm/mOlwZmEEyqP2+h+BEheOO+ybNiANoApm0wVcYqCei+pgd69nayj
ZAfbxMR7juIvkM9wRoclqmpmhgPq5imSFnP0Tm95mtDi/rTMyKD8NcMXLlP4rEMz
7JrXc5t/YYHrinNZdZ/SUYvNODtMzqvC0I9cgvBp2AGXhuqVb7I2f82pVQw1zhkm
P7/16TRQVuye4t0vQE4uzuY2ZFWYcUTWSH2/vpN5V3NHHdN4ZUrS9DK3HGMOjDjE
YafZq83C07tJxrfBWDHKxMJLc1cSAxsb/+SHDZVnJhpzm5YbXbnbHLER5Jn2c5OU
EoOKYup0ntRn6j3zA08ZR1liGRTtq1lZUUDQvv2Jjxq46dmHR/GocuGSDIZe8Veg
vJBulh5g56vFmRRlMZ3dJ7HbS2YFGIKa9dMlFYaFjHssIY1s+LQlkoTu8lwpD7Co
w6zTzP1z74/tFNnhAbdTYotxfmiPJF6psSfRqwlIAICj88LEys0RETreG5oUOqLK
qQRJlOuhDdynbaGpNcD1k5mQobvlD4JSrQkrI+IQdZpXPgMybO/DtdZThRYZgXDs
2H9BFhDnNIBGWZh34n4Wc9pm9RFy28xzR1P9C0zDIsSly/H2QGiZoXEJG4eifb3h
7uHQEH2gio5cMrSuqSzVmajBkeZ+YgJ6GzUJJVm8XFZie61ejTnTXn3FylUj/mLL
j9bdqlboAiqHvzcP0XgyUwsvynCQy643FQFDDZ1V8hRNDcHZAoBHzAH5KE/MBpFN
iXhKrvniGOgPeAXzTs7NELRssGCVPuU6cD84/Sq2P16xtBNTPgLrbkfN2yPBpM+E
Gq+0RXOJ+WlDoeGrL+n7swwPBtE4rvvSgmgkYbpS1ajfOV+Ub/Cu4BAck/4wwy/A
Ae+wETvjN3d+3p3b4dR5o80QjHLI+Tnk1zelqoHe64+6MgwDBzGm7P6jLvrV0amn
3Z943c0Ohgtqms+oh9tloLQUWDk2v0nqeJTfPcwHHdAJIF+TMqo8U8lFwZbwYUO7
EfxvbDzx/krCRmIwue0k4RuG0RuNif1zza/K4Vus4KVqaS6GKZS/OKl9UXV6nthm
nMV25k9SjyJPnpvGOzFzF6BOWdlINK0TsSzy2Spz2wCCL/fdQh3VDvQkQOdMCrGa
lE7rjgr17LZBGYuBRyyPR2Y0waSkaVjw3Er/vj6mYcPqx1/KoUjODccp2F8QKjUp
JUtuB199L/zKgkBt2R45bL+iAvjNe/M26YjRhH8XJrlV6DBurqc7Fs9vcrbBS6W8
Vip5onHY0Jpf/6KcE8HTsCxK1JOxiM/iPjPLthWEX635J0Np7BF4Vgxk/hOns6fp
PCoPQO8nqsTyNNwuJNFL3esNlOn++a9H5UL6hSuvt64dQ2hoh95Nhpe+a0QkZJYv
/UdqHg5f5jGtsO4YoOOTlMvwpKpOwPtnpA3cwvEHupG2LsKEicy35weuNhLRJdOw
af3y0XOiqW9A+irvZd9kRvqYu7qaxcFSSNO0vLw/VnPTwyXHXkul8ncjTeZOTUa5
tnZS0bgTBUWEjQGjwPQzuZoLOxqCrPi7vTo+SJtJWM17X/tcotVKjRTy7olAFswM
hf80znxpgRoMYo0O5619yZRdIo2t70o9YYpJb32uoOog+0RLaYZHYcQCuL+cDjMn
VuOZbbGlN/7IocIFIwrx3WqNXQPRtJjh6e4mpWm5hYg0mb/3d6LkWFa4TSmhXQ7F
8ZDzEsDlJ8z9ypxgdASotsqExVwzdW/iUb4fSlS1AmaFpzHUhBYkrAJL9/l/73Ge
Mq+L8LTHEjJPdJQ1/ME1IMTwdf8nMEGldWHlQBfsnTuAufhW0E3WFcnc5H3CVaEb
p+toBNe35dYUUrzLturXhEIFWZlrdXysHx1P4YS4+yicPfP3OK1ShvkOOyNQ97tF
wPPq5kvpaxoWC54y+F2pqsb9gxs/VllUudZmlMu+Mp7B7zjDkh3kIW3crGPOacM1
fS97jjWXrYJooY0PSyKtF29VI8e9HuBXcRDFfRHtqjskAHjUXgxH3HFoguBxt/Vw
vEbIHLXOmIOO7OwqszqgczPS/eMfq09jhBcI5NU5dcCsS1/iz9GTC1Ubr8fXf15r
jPjjv7VBGUiShUXXwqcqSOXA1R9s7Msj7XGwQLjVbffRIP/tF6GbTqnZ9w4z0DyB
/TVLuECOz9Nux1aDVeqqp7MOqjq5IjlWeLMII/k+Agrmjz8PhejNmEAANB61DOky
+QlPsKP1PsuQv/DkMPHx1CpvbqNPpgjjtgv7MApAEJcTJQ5wyyEsNF8ELUAUSdzc
JR+rwM1x9kUD+mMTbSnMeAc8W1gbhVrzxOyi4PSU26ttVk76/CxRZjpKbXs0U6/h
e0+wD1tbsJKVE+3isbsz2ItKBFn7DAqtkwB6DIoJouiDx5BkkCd3ggX9tjf57qI9
qugrLuY64v0kLcvtsc9XngfZ5CPqgw/CUjkOvDnSzOLJoKcln0MMGaEAO13d129T
lb6g7FKOPnNiZ3l42xb8yaFh5ra2qLEeXfYV0gSP/oO09a05LmJTVPf4fpujTy3P
RaCVg3IKbJAwm+Gmu0lu5YBHIOvREAmQF07NtX3zG7I1Z8wZlmUpd1RQNK9RjomA
H8w7Qt5rt9FOGxmQ+p+1JlCLETzjqIqtPCgKc2sb5Vu/voU+H2cBUEbBZeMEoOrN
KBZqVap1URBfXNHlRiXYPARMLP34I8dacff4GcKAVVY4sGRmzMbLUUjFsc6wb4dJ
Rpr8VLXkA7/bGKTQgn0u1DEXqViD6eSGPaszXeFCccVoAzXz4oKslG7A09pq8ghx
5rn9W+E75tyT9WsCr1GYxSQe6iXi4cbAAF79HWMbG4PUPyiPysYcadyHfxkB5fO9
O9OlnoKbhv7nSd3AZboWidl1yn70gIqq00k53ZKHfTejHwc/fan/IPs+wchCf7Gd
2bFILkQoySY2wK5KhbqTxVpwHWEN3sDhDnz4UUC/kOAkNcyAXcvnvSo4hYuPzll4
5JXtHmiF5k67lwrbdkJKi4WC/efKhup937Bi6b7PEWkk4g+PTW/ZxfARvO4WU+z6
+3DqPBydjwsB2aGSLPLgEG6RnaxjvmfwCe9b3+s/jO9RQjfVf3Nfu2Z6PDyPgu2x
JBdVvirZOqmYv0pHdhUh13eyKAgsEb5vhWIYajLL65+uT7onXrFo0TzWTO/GHbOt
m4ba83HAr1g5SZcMi34wQl/HcUuEjEpsPPvkv+mF4TILUJeh0Ll2yN5Nwa5gFZCg
DtzNjHlJI06ZYlnlc39tjf1KrJy1iAwOb+mUZxvUD6lOBEyb63+CrqR+AKz0/yu/
gO1Dk1XO7WePap+gW5dTt5U5iThNBXnTwXQhaIYqqg1buRgsOtVLeTIPgVPO0uWT
Mz8deaiPhl2dVzPnU2A72AjRmDk6LYo5x5Jy7BBpFeuU0rrnyTC2RN2dkapAQQyF
fUZZmeIAqpf8Qq38M+06BjuLv/jvn95n3GPwvqXHbYMa7t+UlwlESA5Q4t0ZhheN
OWEcT8ur3zsqyEEnIn/YMX04OSkAHaTU/rFOkBZZjHHGjau8RylMDeo8J8oj8zkL
DJxJqcnInzlwNWGg9EPw3Ah8pGp+2aZWre8X6+CoZIwkjAVlw9qbfEgkUwJz5tJM
d3qqs7l23T0MeGioat0hTVF5cXU40aGgJ+/pUHARnENs8gQ5uFRod9hlm2UWXK7X
Ohvko8S+KfjYp3jqLxOKd4FSmLZwhXBT55/4+Jukuy3rA5oVhbvJxSnLscZrrjWu
ABL1BEFIOzZ2gVPXlFTWUCLwX0w0rdfyiBqZQbaF8ZMW4GnmtT0Gjuq9YS8M4KVw
kFOuEQnUaWG/+opIN+jb+oHh7eZU8yKUg7zmscEo9dn7SK9GWM1mWiGIrcGd4mrR
QilxKv7h0RM352JIJ6ix4B+Xu6bl0Jx28Exn0+wXWUOvlFwiKoEDVP/Euy0SPSHM
D6aG3You5PAGCeXByl8LuZDHygHNPz5KUAcftoKbskpJXtC18WyymhE5Q6YJ/0p9
3peWuJQ9u0k3Or3E+Y7OPU2p9xvn9iVfHonW+22Nt/9KUTAZfxyurq/ZrA6iWXQ9
5qeFLNlPiFAeomwwRZoycGRk2vBUZrrA3RKfkuYVYtwErntGnWsO0DPP1fKdKdJV
e4Kxn4eUoVh8m2nOSkHMRPYbf83pcVVNZCQ9gHg1QqU7pOC++V7kbHxh6nz5fsqX
V9DORUBB3E4/HUJpyepOX3N75s4sHDEPEhlgnIe/uoZXvMDgTQXbPALs0VHLclBi
hRC71o9o4qX1zGCsG2ghblL1L1R4pt0XP192eI0FT7E=
`protect END_PROTECTED
