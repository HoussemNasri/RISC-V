`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
La3UxdypfWJeFCepJcMxxU+XhDLHU7k40QH5IyIDv/FmS7mzumyPrETopZi+r1HZ
BeTIqiCsh0s4SZzDNvHYY6L4r3z5IXCfvHNCO4LQp3QJjFnDqjd/AgK/DEX833il
tSsKMkRIc+owFqzae35SEXmx6ZxhV1E+aOHVbGSlT55Lmj+PK6geeaxMl2yGd44m
O6G4aDrQNymhb49E+JpaMpVTVCxvry0L4NSjoC+aAnpqrtNPzle8dP4n4q54y0ce
TrnmyLmQVsDQ7uAIDtAqiH0qfQJ+hPXneI+/AKf3NwBVbwVQ4bmR+6Aqb+5yOYIm
+mP69RlsxRP8n8sp3nmavzs76chg4N94yfCWL71J+QiRZp3G8D8/yOeIomuQ76Bn
K0iXFkySNSERvNWBXpK4cI1bTaZ2NWreUp/3VzJJ5dPeILfhsTbZ70nJCPsH/i5Q
zAtZagkN8tuMuSJ0kJUyVmedidn0J+u14Oyp6Nej9OE/fjTL7svB4GHe/68zWKAa
fW0GP81qQOkTjALTDIwj42U5+CwGowYSYEvJn7HHzBDFt2vQabMx+tOTnQYmpefj
SzjzBpDchkKbrsnoVdDa+N/Fib6DbXqnqwGX2EUCmx+R6FBB/HGvuyqvUH/gk2h4
M+R9lTQhqsy8YBjKOa0sdFIUylpDxY/Yns1p/4Boxoaz55g1lnkLINARls1M16C3
8o2nguLDAY7ucSEXVcnCL01nUVj4ny0cq1M/NhHOYe89Krgfwe25bts3Ss1CYC6T
BA4dqoi4I3SrnfD3Y0TGzJ39z5cNglHwy/0NBuIRF1LzHLW52LyxIWvv0JFqJVKr
2WpkjLGvve3v6bfqCtBiEkja2E7Cce5QS/4QBM9FeTwXexZ6KYDCPgOWsn6ilmiT
whznY7cU/PwbGJoeYWg3BUfkzYvCRSxmh6Cyx7th1pTzye3bPSlb3QKBuxN7lUPV
92BywmQ4NpfoZA+UW6DepOPH5I2bxWfVdpi4X6F5Zp4BPmv1GjS5rY4/qE8Fq0Cg
BwRs+804fEwGQVov0l75mgPoUF6+PhSCwaNh/KVxiYGViCOywbFfduoRYkr84wye
Ojqi931NkvxLR1p2aUETuJum6Y7bOzAq1W9D267oJGI/s6wGwOmqMQRMXWKnmV10
vEEaA8kN+UZWfwJuKtCRwmMUx164b5TJlWLA9JK9dbOgKkDnG5ltdHkBuXbi/Cv1
0+S1CzC21d+X1ko6zIKR59lkynfo2iYKp6zdenSph20fKSdHNO/dacKAxGE5mLL7
mpCrV/Lciwt1w8cToweuiiv+GxrFQIInD0t2eowIWpN150YYDTwfW8JdEV5rKDNL
FxbQ/wG6cSfj+5v9p871ETRvGOM48ud6EMXp47zmrxyD2EsDkoOv5Y4/SZcsyvdV
w/uA8e+z0Kek/rjnQGMLbIQcaBv2g4Th8eitxvJtxWe+Fhf+KZdw3ECVEKoJggwo
KtTipJg1VIU/XtjptFpXFauJGZkSwhMwFlO4/jAuAZc=
`protect END_PROTECTED
