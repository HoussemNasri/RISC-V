library IEEE;
use IEEE.std_logic_1164.all;

entity EntryPoint is 
	port (
		A: in std_logic
	);
end;


architecture Behaviour of EntryPoint is 
begin

end;