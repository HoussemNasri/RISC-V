`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVjZl68Vt42x84Sz041r5M4zJ7XMnW6/5YxpZRgAS+hy5aM8/Z7bIr68lvh9LTjg
HMho0ftYzItGV/vWFWhKbR+TT+ZD6bHYEQI0Ghx2/rDstyGO+khlyYN5u5CiM3ME
OCmUVhNSfopxkxzcy+CRM1yRnpz2zvx5imynNxJg4fODZYy3OrWn6JaAFGT76hQf
pumW+b60b8CzDHHsntzwkuRzZSXCAkIFwnoRNxH53LA1RAyWQ0fVRYak4ufBaega
t35OH6x+MhU3tqLezlMWNIUABqZlgHDFgJy3jPVENbowqMBxWv8YUxrB3E0r/11p
jd+WJPShNAS9N3mIqijOn3uCtEwHz1lSYymLuPxDjzGX6fvsqO5yZseHJsHzFCw4
RtQfCB8UNlBjlbhDP6JlLKxM3fJ6cPtntFv9WtIIIZFbdyI48JimFJEjK1W6IluF
Us4pZ5TDrYzAN/OMhA+ZifJ+en/Jf13kKvkgYqOzB3LRSscdppxcVvnoWz/8Zrar
s0Lo7XnCoDUspVQU4uIPEMV0TYNImn7g4/37/9CUPZ4QOjoHHYq/fcEBW/ewGFwO
Y9R9HowFithxXL0OUqe+IrT4iIG595rbAN9aIzNygd18QWm2D1kzxTj70l4MxkW9
TW/nQYLg02Vorcop02vcVr8hB8Jv7jh/moGMjZVK+oh6r3ab06XtfJ0AD6ZakB5m
ZtjuGT5EadFeFCtoNHeHvu/w0nji1Am1O3hchGj05wEfsGi/XyBSo7zJsfogE5KH
ZKmc824UP2CSPODGYcPJzTlgTvpzARzxnjaP95PoO7X40sjqWHYaidpCuJyk+EDE
TLp6xIkuUh/DPerRp1rSjiuXXUVJDnvqTqqhkBQznZugSULVFCqg3VywGO5xDSD+
HD8ZSHkyvM8o3prI8vmtQrdiHpRtat008YDuh0fuqeH7dYRGnRsJXxfFe7E4JJSj
DouKUf9PNasgLFjnVdlt5RXdNX0XmBkfC/cvKCC90yUzkUcIXzrfHfQzTWJNaPJd
SgsM46nxgdxhyqJ/V2mZLVt3nMAgd3l/e0dCNrvt5KWtrlKxOgYkClIffWzu05PN
6vhpX/w5KTKuz1dcral9NUZENasCfi/ovHTQ7HU6dgF2B4Pz8EG7IaE67ALnjMYs
5GDPm1li515VKxdIo9YS2uFOC3S02xfibNtXX6aigsxoEocHm2FOpi1VjUDyFyKb
8gi/ecx3Bl2o5eRpGLRkGxtMscAbkFaUh7fwqEy/Y7G9KrR6UqfrgTr/ywQZdePn
`protect END_PROTECTED
