`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kdgovTE5bQ7rd6FEAa+G+ElwyV0k0acKVv3fwU7gRC0dkmrJA3PwPEGS/6rvdIb
jT3siaPbDjKOomdD3tSw5LszjcemjDFpIK1jNMmKqk80tOswaHcZN+LwVP+QmvJ7
G3Fm6MA3te84FmE2DxbqcLWjpMisgoGsmCUE54i28ZJphc2S7Afhj1rQjUtasTCn
SHsIC0fMugCW2nyp1mMTsMHkLgMi0+T6MStDzBL8JgJBs9fGZFmZz6aQvHpdpsae
o3grZm3I45BZeJ9JCXO9yRH/vYrqSA/rz8S1VDqMOmbX0Qzo1wglhhZzZ26uOEQ9
+4qWnAOZTXc3XX0/pfbSBIBQvtQDujyRlRklyP6A3JVqDKk1tkZB+Snddj6/fx2S
blz/S7Sz/dZ3igW6CdZp/xAl7332SwGj/eENQol0vpR2bUrpIj1gudQzdmx+F3FG
MMPMi+yPpOVas2JgnzjCjc/Nu7Oq9vR4dHdixqJKV1aOrhREk8+bHUY6rV74cV+C
F9xiPHpitOEDygR4U5oAbOWvYfkvC+Quw2uEgZ+uP0tHdrnNGHevi0VHPak015ZT
kQ1FEnnbad+r0Oh7fI7dHq+OZJsyxNyfjkq0TttXOQTyLB7LYkxLliER8z3RsUoJ
+CycRO+ZcSE8BPtAafpwpsEL8iacumeCfMrtyoqzmEsefI7LMpJB+hPRiAfKsA4c
CJsYhL7hRP1voj+UxhZBquS4YpNIBvUZyoCnNBhW01SZj9ozYMLqFYDq1953hxMn
Y0uyAO3MgX8PNcj1QmJCw6ZO+Yg0xiXoywsmMJ7AQXQWCUCh6MQggf67WH1na5MH
86zsFXWtEIeuwI6JBZEwVcsaWhosFYI34iMAAEQOFipEvE0nWjRJaQlkeExStYRC
HjtWpfda9lnoaqxG7OlnAar7x3TqlgiENWt3eDGxnLEmGDZBG8peAVxcRWX1rQBL
+NC6uAU6Ez8gvxA9x210O91+5xA8n+qoiw0ol/jHrc8XeIJr5dYF0FWvOGxT9tln
XHGqMwLZbv9uCLCf1M7Xm0F00622yDrCPC6xdunM2G2TML6/PQhUVP1L805ZrT/6
i8uDrCiACEaqaKYXrxutozF+To1c97zjF5TVv8DmTZQNj2ilveI1cK79GSJHEMVT
Mz/URUF4XnYjL1zmwS+8RpAR4TWGqwqMbgdcj/7/pMoodrtf5XBkmaz/a8E6CMsy
rJCyWEizTAHhnjbPyQLvx1rqK7jPoYn5jSTmXPK5wjosjz0iSHfGlVvyog0EiVM5
sSTqgTItiqKzNL6AwmEIlfVykTfnwOvMUC9qxrNeBxsSw0GfmnAOQsV7uiCiSou4
oZ0B1sgYpOR18TACZqFxjXoPmWyYNAUDXeaqP5Jyeg5EbT87zDaCv4Ei3gVHdNC2
a5TknNjTPyjPkSs+uHpdoB4JfP1jHx8sLQL1K1zi9cKyPfc3NHiQethCMfT2Lztc
aDqcCR2XE8K5uXaqAn/KmMX1XcYdGbosdTohGgNP6XhHlicn7xmIFeDeSTFH4noL
OhUEjpa8Js2vhJL1DBeEotaBHVRjjBbQcoyg5cpdxccn1aRY2h2VcQrFcyEmxFBz
6fFoPG+KzfTBJ1glXzPsJ09KkzbgKTgixWL5cdKvCto0d3huU7seQeojXjIq5V5k
f7TgJu7nezwOcQgIHZz5FBvY+eMNELVvYUiI6+TLwXZMKZ78mZE8nvDYeFwPLmW0
Up/jkZgCFnpdJtSyZNxIXcwDzzGF9RGNZHuo4mHU7eadfbyF5/97GTWBAEy1BfrA
b1sMBRj9dJuBo30qV2HSog21469nozmwrvihG5ThqAXKpBKhHMwZxhBk5uXEFOjk
IasE5Fhg4/iB8Q3pol4hONXmCgF2JCCBYb8lYxRJluaaWyt2MHeeOYrLSrXM5Fzo
EDwkIQi6RBpfFKJgu5Vp9tznFn+T9Ru+b7xOMDthyBkyMN1TCu1bhxz64dFFDPKV
nEEFp1uXyPK7og+cEnMD+3DaBxE5eKHK7nJyr1ajQkjljhCu3SnX+SUZ8BFAUfqF
m9NkQDr3KHqBZpN3g6nAPjKS83u9sz11ElQRLGpq+rFWMOmMw2PT4eWn+3JmvJ2z
OOeXqqgoBxv+X+hvZ7MQ7uLne9xjQnKh4eLdGsuEqP9gscoHdHQlPl6nuExXA23U
TQCho1vqEwXve9pnnmoj/4n5/GpCjwsDKjCaqgUpXAi6z0y2IOkNZ4UCt8Fd6Xdk
cxEQu6pJD7NjLgAh8TsfIn4C1m6H65D6+ZqiOI6/lyRAh/Y5ozUnuQE/tYUxXMWf
Rxrrm6Fw2nCVI9OZNQqm7XvyM0Kk8FvB8TbLxOn3FCF6LD3lI/1jc7QMXnpKwtTG
rxrUHeL+LyJZ3nUNWtPrkIARxEAqQDwW+/E8P2nixpV3SjGgoEPuM/9jom1Wk8ZJ
3WKZ75mTcFrdB9L9zDQHb0sBhAbx/b4+HkcJ6CocAoD+ixs6J0XSFngev5cik0aD
d+Xthr5M7tuajmmEE3Z6att/udP1t0r8tfnxc/uF3H/DpLv9MgRdLZ2cTuKtbNjA
2XBQaZLL0M0FoM064X9Nzcm58ZAbQmBLoZYZHJ4+8/ybwZaGIJPs9eNKcxqawwml
5FObMcjRAHjQgIb8vsSTavP+B8Fe5nuEOAcXyzXGauuGBDJSBnWo2n6Q2JVKSMkr
2vmtRcl2zABJEdpY5AXvpkXBBQpQOsm+vZxEp2DztF/0o9RtOfQEvn2uHSsCRp3z
4BipLhUxQq593GEOUApT+2sR98/KbiQpcJ4Vvap8xLEhQEhxj65hfNhBJKA6no7Z
5G9hklS58pQsdd5F+sY+kFgstWUprrVOouWmxF9tYiSLdfP4arWd/+IHELgXZgmE
kmGdnviR5LG4mYVOjsolAmi+DxUEgqKFWUFM7UdDlaE0RVBFg+JnKXDxG4xn5eSi
8QtFsWT3OTBt9jrDbgaYtZyQwDZekyuGJ4Qfg1KYQ/1FUDpoNbEutdmMa7Oy0TLu
ddwuflUxhQ9blh0YTRJnRROFmkjdLnn2mPXfPiSLYFD7jMgR/5kwf1YeWU7drOkm
e+kBG/42iqYpPpXbbHsu8eV16cUElCHiS5ZBJu5CmI3rmev9DSEuz3ehNkiyO/Do
ILrv3y9YQx0TwAjgvhgVgviuXz/1IBk7UFzKRR9SHicKNQegKQQm63e/C/ABW1R6
6B7N352B+Quhmh0l+dZ4jAIVpdAXXmKNRnP452ixjjg5wwE3/sbVTMRNHDBXjveE
AvLDUhGf8QhDoGF87msOHROD2CqokSNcUcEp3mSnSbbRTkRjcY7i5L8d+Wq055y1
NecA4f0U+Tf3zctSEMwiE6qJiIo/yJKWFGl0fYe3EhmWF7xeKRXDETpX+nj+Us21
xGZZ9ffL4TrGJN1L1niWfmRl7S3dVsPfn7e7AyNCYCgYZS/K4c5mND0euqWCQkwg
F2CnI6I6mu9YsU7tEy4HMmw1RGvw4SmKTBnGlU/i3BrZuk0XKnLG41FXQ1kEjouI
6qtas5qSsBvI/FDeKv8WGPO/uzIoB/XhJUPcYhuAkdgeTJT3fQOd9xs0d/Ojkg5Q
/p437a69yCSzGE92TGtLb4x/nzVAT8nWVYgGdm5eFAhyQdWMdSo5rXyDwGyhyTTA
tIiC8jJ1zPGgkkU8TvtBU0xvwpfydcgN/q8v3MpbVCqzSl9Fsp7CcpAnUjBh2Oiq
aJ74CoaEGk6Gk1OyxEliAAXbejJfdD21kRNNyMhnhf4oqImDPEJRffwGXmfBb7Ch
1kW39ZeTFIHhKdhbpoYpZmZlRfA1++yek5uckdUmlESZxUA+sHbjnNBIOlLPN4TY
TeSyxGTx3CmgIkApRExegmVtZR9aF0fHN7sWOR0ga997p8NmhxPuFHS+xz37SRE9
v1Od4H4/s3wfxPvdUX1xzsKnC0ULTO15JugSzzBbFyCRMS/oTdDIHxTu5TR1J7j6
9a/uEhAW0WRAxHEli5yIEk7q5zIxpBEwBpqDf5Uv4NcR0D4XPSeiMnXX3ttUcQ4i
u73XNRCKlldtR9f2yL7tuanM1F9YewL4wj8fFnrrjw/U0G3GNcbEpZvCrGy82DDW
/rdISW0VJsSvxdW3tcYzZHYntAk5PSqnhV/ELfHcAH5DUrYhv/+QlWmZYxLMaDC6
Y76e/kNx8Dx2nGcdTrWNx+7+6Aepm/ihV4IpMUAHPnDasAagqR5CxpI8Qr4Uuzlf
/wbBp9JcnjbiH+w8yKZ/EWpDKRY7DKUePOkkc28o13G8invb8wjESbB5eZKd12yz
nWHzmlK//UHCnnJiDqYR42gWnPFAxYuBwRg6Pvmog7M97hbTZYHH3VYAbstjJyFE
Ur5BtQO1FeBdMXHThB6dh3eyVTGsjDJfV/XBA/N8ucu8Us/xeBZA6LTR5EDhEksz
ovOomZSPNSOz9UUTG3mNzgdacIAfCCvn0AS24Ox+XfqiWWW3Y8S+mNsFh+jcO7QK
O6pd9mvrAOIMYFW0hzd/Zm7EhxRsEb+iLTFkLcCVM8XTf3I/2cNb9Un+puo2qCc4
MfKoiydDI6i0c2YKNnen1YXJevIBWmhPBlZKQhNmY1cG7a/J4ci6C/lc+G1ulLG+
mvHm31NeewefzSWHOYHDySK2NI2sx+dnbDzaCfBdnv3QNNBdZdQAmOMbswyL2Q1F
6kTVJwtYbljpz/TnMql5FJyijisNf0pihDCEj5XuQtckrC8c1HaarenR6EYA4xp6
y7hDILCx4kd8NpDjImKCiOh5AMDI7usSOPb7NTXHuMnG3LAyO4ENs459hwI/tk+d
81cI9U7kCmVR9YuRwbog669zfMldDndpSrXhQXqma4tSPO7rgWlJFrPUvgXJfKY6
q6dB30xPs8Mpsq63AXIS3qmuK+XCJWqZHBY6kIN3ZpaQUSQw43C+asbNpm+nIUSK
RXKahPEKXotMnPF8M8Lkv0xcyF4I+CUMQKREqVr+62jfnjcEmtGnrj/0YnQwoSrR
nsXv6Q0WIFQQsdOmu2dbK5bDiL1eGKB/yRxJv9urbufCcasxJBb+P5xt7N1xpMWb
rSrjsadMr9zmvThlueaZVTRWbrxDW5rQJNrai+4eVXKL6Tq0TfQZXniOj/G/NZ1A
R1O2UHbFDcWNemPIpBjVBTwVwxF1YnKXg7Nm4ndaOCISH4FaK9eL8ilU7WRbONqP
tu4E1XOzna0CogdbM38CS5oNip1S8Xl5KZwfCeOH42m8oHkGmj8pTL1hTDjeeWne
9kmAiYMbrDifn3/FrMHykyk73bJYV7XikhgqlI+7C4SqE6a4/h33kK7KsUTERnu0
kthg7Tf4tomo5bxWqMBidHrV/QFFy1SHzM4vxl1xyRRrEk3i7qukDwJlvM8n7kC2
y312lEP7fNFnEX8e6OkW1hsO3xCV9Fi0qlBzD5FcEmNH3rSXKb8O8D0mDOfxhyTL
4KlolSXh2e9fWHAb+uUpxkLaUW0kKALw5LvmDz1K/vDYDFtriPuCA2HRAEzmLMTi
4Qk1TzK9Zx6C23sBJF8P+xM6KLtPi1nQ/Oo4yrA2A6fsBMXR6FhShbEuyzbY9l8G
1L57YHfnZ4D8tZ1OqiU0+ME7/KEH2bVhwmf22DV1OyEX9d24SDBAffYGsfsMFaRS
EAPVYz42d+Q/4COsloxljp8vu4KYDgljhIm/CVzj8vhmFoN8/3muXs5ZTCvLleNg
WepOcs+xN04nGhvtcN0PSRh7L9xV3thAvj7birCW7448FvB9nW69KATYuFf97vUC
SYfTk/32wy5gKgLXam48EavQ6sxVoegL8KcjDOsv/OBPtPYEw5Sz4JGY7mRcsEMz
94Z8TjHg5fhaZEhxb8PExo+Bu5+xjHIdP6LJWjKAIqoqzeviUD71CI4PchwbbtJX
gKCULaK/3uPThoZWnodm6dPIFm3aasLEO6GOfL16JNO1kzdefJ1gcn4BvTRtBzTR
u57/+7lB/H8tkjpzeeE5XQLW9v8N1N3O8snRVzhtAa52lK7TixF0BBNDbnqYgX1o
R2pZ1fCrxDX5lzxVhF/VYs1QMUL6AOIlfXYEpX7G46w8c0+eVaW2luLeFp2NYe3d
xb+XXYOh6hPCCTOVbi1E3lNUjxOv1CBdreXZHuOEHJgVGQoCCsgalx0vEBdgVfSE
74Wqqi2nnzKj0lEflFXZX4sRhihctXTX5wFfwRowOkw3i3LsMPuWFUkW5lq30q3j
xPuUzkIXMJxFCt1rwLlnUEr406DBPZ8eRwPrFtyBR+m1jdZN4yK0aR8urKabRA54
oRQBcZVGTf1gXj3ONjEpP9AFEGheu6Jl7m9hZ/A5IhWgmibNoimxvwHl64UCsl2/
eou9d4V7Niv3sUAdqSRl9+sFPU8NYvnSLEfHYpyA2mAPR9ZNnRvdiK+SBAMp9ZE/
Vl/Iy/t9utDTZ8vE2cTnHBs8kUCeHYfVtjf0IiRXzNmMs+Jxn+5+evjPzBVvWJb6
abhSiRQRZwP8BkpGC2T1uZURH+kN2unucvHqcIpXs7qASaTCgCEwpGqFVYQu4Ocm
TU7FH1Sh4kV4LCPw+WvbRv1UiJDIGk2iKY/GvJG7wxk0WKvCVf6Cgd3b6M79Qtap
bCDjwm45rmOf6SjZ3/WWgwIA+X7pTwHsa9r4ttNV5ohQhaMOiPKm1ZJS+9HTchqZ
+WfmQg8yyA6zF9YCROvDosFjJjhPHeR4L8MST+go5Ema1THhDd4lZ+jYPwzmEV2U
ZE5MyB7jebvlOGtTtgqb/Wk6KXu2WZCO8k2gwltvF3d+DdR1K5sZqWR1+Hv9TM1f
/mbiF8MM193NhBvlGX3KsMko1CFriEbsS7hrSf1ade2XFci8wKT0kNahcMNTBw+i
KRsDNgoEYFW6PSePre3QBBaQK/MJfXzmCP/PgurJI4A8gYfpegT+mlAUFARG4TXm
LAw9XgReMYUfPfGtcpe72hLtq2H+DGGO40k0aPS1rn6gI8q4b3LKP/msagb475ID
oO7eqHk4aQVjYG5CaeIjoRYT0+7KMTQ+bWvhSTwt4F2XAs4U4m2hMhskm2ZJTWXK
+/asHFVg1lj7IimAslktgOHDn21tD06PE/4bfqt9nJs8P30kT0gxkuhro/gyFklW
BKRYTGJ2pUYY8GkNizLxOVxM0BNwGVpQvRIKGaoPpp7VzcS85nr6h/fOBp1xkCL5
TSYSNHvN5y3aFj/cEWUUcqKWn2TTNsM4zZeA5DMru/WMa5i10rr6hUzdZnkdhTUt
cOI/I4Ij/Z720w7MoxABiX7WNEHe5b2aU0GYYIHauFPuo5C1BcgAilPhsqNAOOB0
yWwY/ywol1NjSIz/bYatii5KHju1WrsUKm/skiB2v1sMibClQK8WCtvfjqbIo/qc
ghJKIRllJsQBEywo5zllK23dGLFqY0fwVArx98sZvvr0QsFETn+6NsL/HD3cBUde
HYNaHfw2xxU3f9IRb+Ex0ShBa05ak2mttADS/MZW3F8HiH8+Fyzka2cTor9UEEiZ
xpq4+YalNkDqr7Pqk1v9j2meGv2VEFJoOWLrJGmyXF5Dgpp32EtxSN1IQL4XgqUB
dmYKhJOMnwOeQ18LvKLYcpZsNfjx13i6u0cGJcB/5TMoOXyw6paY6s4un1CAZVB6
0RPmy4DESgdAItFo7zo+5kGQJjJzUeth85PDYdB0+O5HElfNP74QWWb5/hw0lbef
HDbEoPYeM+DHQcmXIfSXyFNv4cwvmYHTFvimk3COzSsTulsGPHWmc1qV3H2GsO6Q
ApWCHGIjqPih4K+sMm5PcDXo9jghTvMuC5yE6nDmAfYh4lEeDVQjEKvDYLHUmFDw
jCnfmAbqdAmX28dgv62KlBB5jfLHLCp+xttI+MqDbCbmuMI3sclDoqPaYgmLLt4K
wC9KMLa9zymJ4Exz8zuv3f8eIfmIvbh1ExNzyrh/5oaJf3EQ6fNSzVdJlvWBHGzU
CBQlqL4IAuh+tXb7H9H/4R9f/5YwVj8QYkdGVQ2CpAKgOQ3dFUHg8Br6E73YmZEh
0XCQPHuQBGAmRvJf0BgP4RZy8855hL6viaVHC2gQaYZALfGoeUBKFQ9WljxYnHGM
FyGHTmuW9nClfAQcMiQ+oa4OBsEhhtkH2D/4Vln5AFsdVD/FRIIOZsiHGgCPR1+K
uj9yUvx15kdHZzK7rsTHv0/yhl5TEurqG203lxtocOaopY/yBKNFN+wYYhN6xwmX
EJFVRoikakzIzSyATttQk7wZ6ruCEP0cQJ0QNKDRCQuDqx/L7IuqIxs+rUW22zMu
9yNjQqz9NxiMED51kGQrjyW2ygPYpAr+r9ZBqZ/uo9tq/X1wad663X7tiAoqHGCF
cLCGg75CcbDYHYTKlnRMkjTO4F47AwAgTTi4426pl0DKZ22lAxAy5aV7VDeJOYq/
UFwNo5nF+kjWrbOXh0Qk+NAMKyuczyhheyYO0xBWCww+ET9aVCsDi/M8dth3cKah
Iin8Q6v44Xt42P7hmRAHe/RAugr7KvX1XGydt2JOq5Ilk61RGJY4dtAbjdiZqcW5
KmTfr7oEbv9bvF3al15eiHWye302yAQqlOUq8CwaVVvWsqwCVje8gZaoO3sC8hDi
M1+VGTTjQcLCYUUgnRc5aq7JcYaeBA0RUkp2OcXabn17TiSj0QR/tzPeyF7gDnv3
6FNAnNWcIjIeWQR5+WZ83iwxSFchh/zn6yrPIBf5jdbKWi8Uivq1QL93G2qQaiAz
401KLRPkkRSPpnhNoa9i5qSKwl4RpMfrSnZes329+n3lMWREdLi6bGF9aQ8Og2kb
NQXprxstBEuQUpUwgUU5pmC/Bq1rFGsxXcRBnFLvquIL19aHYlSAtRQee5yXZI4V
7A8d2vqWxRAqkSjeVAAw5Ria2nBxfXLPrP4IrpzIxm1hJstIwauf10dXQ1XgPCob
hbrfqgZISjqzUdq6219z2pmVtp0GSbC9KR95BvlVVraBu595rw5a2HmbjX7RCNyX
KnrkxJ59rBi3OtKCeOUP1dolzuBQ6iHX18ZjJMqoSQl1y5nEbGbkrBvyl6UwYAJw
Byb3OiSdBWCpiBDacp+Go3zPCjsOfCY0nWl2puSg7ckg7UGAXkIM24txuhpFJZLm
YCyNbfAcYQaKzw93JsUTsjVkUe3Fp0e0+qEYcX+DsTPBGky/oBlCHar0RMOdFVpA
JkdfoJAvy9TSZaiGTvYvdJfp+doACk66hnrMtLU9J/b2MUOO4l6RQ8dSVWzapyrl
zNTQ++7/G9BwtkN/0CaE1dUm4nsD4tcRLskuqhFP88ngMD75lFdFOai7/SFg0m8j
e49SnjCzlPOIdZV3MZBNZLID/sys8GncjskqIJiOiqSOEObLOnAgtw4eCZbJ7DLV
cLPX9bwakCY9RuAhHteGHYnCSzoL0kJ6rXkhOHZ57te4H0vurshnrPfcMm9pPihn
O7AhpJMg+ahrZh/Gnsur7D4bMHeVgdDOFJq607b2Dcuwgt7eal1p9dhNNdx1xbz9
PXZdFbmnc4M+mO2LGCcDKM3TC24heDFDQWcPfRU5U445shzGdo9EomhRdjpviQPi
JS5qHZ1hNhdOH8oSelw0YxYMBSuyhtDbT1/dxtm6DCN4iFHm3ubICAfp3yEBZQ37
YlkSVl5+mX+OPmQPxvqHlIQ9eLzb1Br4e4PPh+93P/8o+3SwgyhJeP4W8UHT69h/
GFsZpW8fkWy6XECeXrB4jGcPzYxzQlSjnDyg1Nw/ZnYN7lXSfqOiA4xiX/vZEmtM
lMg9Mle7RG9ptc61MDmouAeSBSuLmjhJL5bRkbZborRPz15V8E3c6kk9MFhn5tsK
MB/3LM9K+W1hzhhfFBzqyL6OZFAB/tulgG+/6nTCHLGAMD+IC2i66NAqGf0uDccb
OLIvnT+IClKIhCJB1SHknK4XhC6CdIC7yKprTyPVXn3OMXd8wZ3Rvyr0bLQiuzuw
sR2ErswSo5hUc4K5Xr1YERrJCgd3kHwlAp0158v3QGBEb/3zqpz/8/ILd3+bsipm
aT+RF9lOaE3NyHQEuSpiFazml2jjAErq2HkyhcHXHmZbw+RURmtLGrV//1P8Kzq+
VXIA60pBm2LzjWeyNUjvJ/cwcqWrzSaGDPd8g/mWhfgfbV+EMe/E1qM5RiYqNYaK
lE2vNG2w42UD6oh0FL6Xt+qCKuqOZ+voyN0OWXHI5fL6jytwxvwbhKIvtCz43dQZ
VyW9j2cRDd9hKTMYd69zArYnI+udLvdp2/lQYF8f+zDEpK4DD264GvqUjUXBlL1J
PhlsID28OiOmT4dqXnZJWj5u9TDXEZ+h5VJ7XBKbMgOjehUFaj6zkjzwIE2vB1Fm
ISep9rzbrTAShXfF4QrOocqv+gkcSwCmWqfLwVNm22FkvI8tSaLYMRGY29VKfLS9
zCrD58vdFMlqkZcxq8MU850HY4u4GJhGbTJi4lVDNDDUK+L5H5DKHUkAOcwTEkaq
S0LTTf3Vs24mkYVtkBVgOV6FgcB/rziy53p4LWomBKQgTs5Cs2Tgpxoj4r7l8xCW
xJFiUeuny61qF41U2+9OPHnbFK8k0x9JmQIeBjhgvlbxffTCsefrcaX1RJd7NDZq
kNInRxK9MrKb2bBuJChC8hCynCfeueB2pjEjFzTZxHr1H1Bk8DZAgYaYgtsedLhr
n8N3eqG/naBYccPaSshvfd2trxaLyPJjwZErxtf8+xhsSK0e1YZkH7najNswnVTr
9QszU1J4FziDy01zfJ96QoN2VJYYjmCPdWojZrThJWshP1ebJVUErVy7ynszck/Z
UAY7lI+oDORmpf5Kd+0xgCYIQ1FblNgC83RoNGBZSSmDpmy/1xxpa4RV+H7eaYrR
HteiGFsiQlz1OKTwrs8JH7ZyABPrOqWPbbqJMGEEggGnJJOq42Ku1VqaVBBOUnDW
ZHZHGEkD50UWWm6Efa8vyF9vEtvQr/weg4WkfktCnM4=
`protect END_PROTECTED
