`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLZlZs+Ln7m6QDPYJJbsBktwoab3LQI/K1BvofRmWuk9eLKsr3x8rqxvPmz/hiAv
s7Yz2l/0oIiarq6lKrOwVh9bDSFNi4U/Y+DRjgq7VzfmPDEozgzp26BP9lIu8hgs
L9ET9JSp0fwpQE6QRlQ4LxXGPzdChPESA403jvYTOn+4Pv2EN9l85AtjTDRXUSo5
AY0KJJ8HI6WZISTwZO3QyfM6QBJMCzOEO1T/KyGnNPt3Bmh+FIBbmASbhJ6EsFKh
hB1xROAvUr9JAKvs67SD06GBvASShFYhp+u6npZ1fYa0H5+ITHFVNzySN7/aA5UW
kId6saxPNHwc8ycQiRiGRF11rgJdqYGbhTuGc31MKiGBaiJaWeuXhEmbfG8Q1ZGk
b97aVo9F5eiHRlc224GcMHIyTKOBXgJjqJXqgkVIoe5PfF7rXNEDU/LTYXfDtH47
QZiP5Ibd0mv6XLSFuveHQGpHGhEvyJ1QeSLTfXq8vCcRTWv+qtfxU5yrje3VQKtu
MPlaGVdSLdJWhkQ38Npe+mGibv3Va6FabvFJE/BUz1a0qE0TE60QhnXEnhIVgAiW
ydrITJtwp1B4AAMgo0jGGerQ8PctkxLDi1yDIVTtqoPEHLhdNQYZbDQbxJSIBB3N
VIkp84qQqGwI+sabRWiNQlxoqwGv/HciGC/DAs3eGAevvdPW1VlGqV1gqT4NcESf
sreP3y48tOqZ6/zJarot+QY5GaahCQ9cz97dyuM9DjxLsQzsJK+JOK8/n/V3P4Cw
YBS4y0sOwV7n5EcOgLzfVeqqcR9x44visayC9LJa02lEwpCGxewth9Sn88j/mWLq
pH9UkSgTKX7Ckif0X2yCYA==
`protect END_PROTECTED
