`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nq0DouqLAq55nAPqQZ2q3Aj4B0/dSCxZeWrHI+FYyUf2h1H2DjxVCXIfNXyQVgJK
5tdWonXSWkeyOhzUt039Y/rec3kSs4w6OhxH74axA3ujRc+8Jv37y3jqtMwZJ5TP
fqStrbUEdsB2UQCTl10e2LTwXGKbsmA2MAg3Uct8STcPPBXh2++ZGjrlN5v1rC96
tPoBAt+yc3hMe+xM2sgUTFyLh/MUY5by7jkZ/n6J+yBYQKnivOq4XoTkj9GMVGgP
yRkrySjOePIhI3IJZxL3V13qcwqPWBe7SHV2EiA3goHE/0HUCQ48O+CDcoQz9cda
+Kh7D+Y08tq+U3R6trmL6AlFisDn1etFEnSRtu02e3VWHXP/37a8gVkd2gBYoCMD
KAc8/a2wHDO3lQwff0Xp1vfVPp8rEQjhZuaYew6ml7Rm3R+CGN6/MooKC3aTWldp
lnlhXX1xI9U5zfqRXEfJGc1xs9nKXjQPXIHUE9fKcrBNbfKC9OoqmnUcFvQUkQtO
ld3YljgkVFDvXkSbLOws9s9lf+NPvvtBN0+uorWyI+leLKYwtviFL1MLPY1l8XaV
mKTRSpac8YrIm/GHk6DIAswMm/heqMtGSQl/bsMHfYduje3ZeD31HqlchwrgGDDO
Sj9vSDUUkATOV8LYEt1XFjlQmiqVVhQFPp12ZhwrVQjY4QhNJ9KCx/1Lg1UIAbmy
JucbP+u97ZbNTbS+LzU5nL93EoYeS4PKo6RI2NDaumFbB34pa9eiOr2pxRf9Hxjw
4/oiwv5ww90/IaOTUa98hx3afErl1z09CYTCMQo6xCGABdr/PAidMhhaxnYxwwAc
iTK3lLIrKLXh18CuM8t1MAM1D0x5TMPD01LiD61JBPKJszsKkiv3KM+0Ysackwc9
wIusA174UWeqUr8dPOhL+DO0XTH/usRzWXofmX9udwcecS8jTFVqU4HtlRNX89Ee
ZU/tcH3LS4sOxha/MF+farH+XVFXtKtejjyllel+UxGiydzsASYrlO1EeR0GVfED
KL3emkcW77xGruut4zJhO2IFcWgLYsUm3u5vdMZth1J4hHQ4Tw0WD8Y5a7WuMHXS
1fF8uDc7hT4J+MWD7G1flGSiy6Ikr4ZJUvRymN6jflKAzmI7dAJI4VdUWixGWvdQ
JKiju6IgIoniZejEpaIPz9hZi3I1M0NQjCsnez/CCOINONYEWTSaQpyWeA+oVQ/M
Pdl7n1P39GW/QyRKOE8oWAjMwBpLL9KbuVoHojUx7BkiN5Ev05qijdm+Uz9uPJA9
`protect END_PROTECTED
