`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/q8FlK8/fi2OyLuOpdzirJxwADR+XqX2/3dAPmmD/ZYlaQ6KOxYgJQtwK78tPuC
AxZDcrcIPlVBlTKwzMGSSypJuU/yyJ/STOXpE9J0HDqgj3Pdcekb5EHUWlwOfnaU
cx3f7FwE4PBftooFD4i5J2VYw+AQIzwKBOc/zrCkQ+KmvJrViro9QNsYxS2bf5pd
+I8Z4/aL/atqAk/7GWluDVj2bDQnuO/6VeaRtC4WLHpKlSRy0VbqRnuN5JsQJfBs
D7OxSZpSPqZDuEg/O+tBp6IaxIChEiTs840P2WLsseaLwAsfHt53TJJRYqebti3t
K/qfAPg+oYhPj1iMu4Ws74nAT4azevuRi3Jxb8EywlPs0TwNlDNJxfYNYtynovgR
FiA3fZFtdpubCjjMWxMq0pd8sK8cL1D7RIsKmhtB8GsxBHIXNuG4V6p6M5UNw430
RjG0lPw8FcC7xWKDVgxaxdyaODpL/GvfiC7Rig7Ppxs51Y8iXjUtqNXczX25L9HN
Jy+tFGohw5EJw/bwF9EqSADCqeBQEK81psueUX8jetygg2mxqINFESMPZDZsZ7+H
w6hmmx4uLyi82i0NuwrhykMT5Tn/VS2Uf0OGPDtc09oblkxsrnLx41ec5iq4sp/9
+4elQWF1Vo+/CF4szDfGDbVE4D3EMiO+sIZ/SDNvU37gzcrkC0JV0UsY72WmU/5/
P/2PLvrZtCykPhYHArjsBKzTB4yTzzlEOVrBbCoQRuq3eXffA4Bbe+VKHgp7sr+Z
+4LtOF1k9TKCznb41tG05KLFcGQXZUjyVCubCxvUXQGQd3zhiR1a09rBPDuxWSht
JiyCwNIN878ffvg6p1CiMn3weN63/OQOXj4vHcNvKXFZGmRhF2n5Tf3GbOyXNenE
hTM0JdRro+glICaeljD80eBro2Jq8uZ4SB6KY+Dl70o17DWBErMqMrX0PcLTz+Gu
7jihDyVxb5VGZVfUqzuT35Uva+bDVg6T3bAJ3qoOf39NFwGkF/WQ3z1ZSKRgQ6qt
H5P0nj5ukGU3sThB4K76Bwx7JYZGfCUZ/uQSr/Q/OliiGax0kYBYperxVWf7UOSL
OtXjO6kM3BMYhZCHq5cTul73boEhUJYEIhBRbhLN7qPjx6Srd5dBaDRAt8gPT5rk
f7OdSdvQNL5DDPi015z9Ml5GZW8eYiWsHsJG+gReW/aqp/rzpgDVdGeUwkUnWhWD
52iqYzUifT64IHjtaXrp31Bsaqlh1Bjw6C4tHfTkbfOJ+v85vTx5S7AYpqv7IoLn
marux5SRkqdzaWZOIsCjbAlrzmhW1MUs6h6mbUcpxvNMzeY7evOv0wRbnoFN4y78
jczsgNAxKlUTjMVzGL4B5K6tYKQDm6/gueTgZEVLP5DYG8wtNb/KAxnvQJMPZkwe
vU58uZ2d1hd9wj/6eLuaNYWorY0mCrk9eADQBrji8vfhDxQKkSxabr5FKmQFBdcW
JufdV1Y8kOoUZZx2443AF0bWQNc8TWTA9dhYOGksgf+52xiydUqBgadX/Oj3/zDc
0AfDUSZuwBSnz8395h9kBYio2f3FM0nY6sqvso8w/BGXnr7O6q984UqOqtgY+aM6
HHaAEjEDX6oHmtHADCjP0kyX+cf7+LZqWLqS0j/O009atw/dFwakGwCq5fTKg/KW
fL3jPHr0f8ZvCXLGdDl8q5u6+1064w5jLiq0gbVnCiFmD0Lcol7NEdgCrGz6sP1x
CdkGNuRdlbPvk2XlBKSzR+3tlhZs5ySa6O4d5StHTjsiunYCTgTo7l3mL+cOayiP
WJOKq+xSojgERkSV/p7G7LYFNTvQVZeBlSMi/GgZZu8FpqJ+6T6CKyj0RzkcBGbR
UA7cxVYNvCbg8/RcWV8GgFD1WbLPLKzpUu/ZXPVKkinE/3RHEm87Wqtkt0l0Fqmg
+fRbBr2ek4uHAnybPnPogjGS+iQpYDfN08JQLoG4K3Ds2B3kBfvmBOExRy9a1OFj
rPwgUDktf3CMwuj8rvxPeKbSxTzWWSeXPqfqG/PxyyVNlh9sv1q8HVlPkFoSScBd
hZWsls1oaVKc3pcv7r2FLyCn0kVuUogKnAsdfLJxx31Tnj5IqXWIrmIojA9JnsAn
v2GGY44BEuoTQufMaFZzTCjHDanhuKRrwA2prZiMFgupKHtYLdVitsThZXUsBQIk
uRfkNY6pamvDpuKIuEHa732lqwhN/b9EmQ2PyEdyA1uLFgUmNAnd2ntNrDVRmrxH
ZidDDOkH7EHsUZeg6vEmttALRQKeV35CUMsc2RH3c+Hr9eMqEJOJ0pHWXBASvNEB
jW7YOGu32TF/NOc46MtaqDKcAv4TgtC9Y+xUQm/ZHUYGRMZ7hav6Jv265Uaxus60
NGnWJR/UGZ8QumUZQeY8e/V4lqGYfNT3dPIHOWCzbu+FM8rQVopQOvEb9VB6AKwq
590t51fybM71AuCM2q0XGXES4HICTx0LMxfgkSYGf9dXY4hsuK5mbLqaZXmY+6xP
EUqj9ntrMqFutedwZ3cD9pt5tHq7GxDLpJECYCyi/JJ7HTCd53xAkG6v1MrI9P/V
HSFYXQxOXTldOTLl/+9T1Ufmvk8RD38/nXYPKB4Z58LiWha1Ifc12xboibZ3QslK
as113HoaQcGy/DqNXMtK1semiRajfMoQQ/s8nznsxFmahZXWLL3xV8sDOpfs8QYa
lRp9R0D9566TP/TAM92IwCmsa2ungfIv/KYgFLxAgF/1wDrpZnW1EfIUZ1fdAQ6j
aNSCF7vI2M/Cr7aW0dLwiSWvjSF+T4Nm9qOEOyKWt+N13xlhXNvEicUUTVf8dIeT
PA9L5AzJPZuCRYK5xqebMvKmvS5SMEprZ4XHFh/nNXSYWOovNmsvIzQYLi/1MfmM
ih/t4SSe5grN+NklPSIALK8KptD+Ef8R+ezQnkMyrr4cfs+LJ38tLyV0wXH2btRd
9uicOx96KfiRyTbe/Z8+ce7/EtuMiKPtukeCH4gYN74wLnEJMMz01RfW8mEvYprD
mB61jToLi3xjo4HWPPV88Y5DYl/MHZo/Bdnw3W1UD6+iOcEhAr4DdGa8J535CpJe
ukoP4TU3SsQpt7Egy1yDFrmN4H8D3f5VtR2VOKKvOA/W4PwbCiyUDCtC6SXdRrm2
AIs+EmKXXXT3+1Zn2FbaE5lJbvObxgeqIlO4Jh0e77XRDlbLBkoPGX0RBI2ZIQ9F
ZmJWZ216NlUjUmTZQTSeaxapDJ5q7D9m1703l030BSqpBGUobruJYCcTNfIiKDAy
fkI7ESvzBij2iw3JZWSNBeSvGH/X6lalJjmg2nXqotKZnE4UGtbPCynCyIVkASYa
AHj7s+b4qqO+X1ZAHE4//QgVMcA70+9IQDomJ2qqN1+TCTQM4kwZPBYUkwOGdxah
5bRkUv0iX+tytpBoWMBA1ZHwPv7c012hYfP0v7abyXZzhYUsmvUID4gTBOjOSnoG
x9NS4EOo8npRBSgSnLezBqAuWn02GHKjqVp8rBzs5B048rwT9Gh2ueWZqAg9ET77
IuVGqtZ2FCJhNNPOeS01BhYTrirXf6mhmGLVH0uppGbtjZpQz2TocCke2SNw/FCG
RiY47wfLlwf15kh0ZqTtvCHX02lTvBt1G7vi7iQxfKh8IpTQCzRoZNyaMgjSH2Hd
EO6lCBGV0xY7i62YjQFPWjS0hqipy0uxrLr4wsy99LjS0HRBFfuoUXOuKWHW/BFY
p9N1NVLAJP5jN+c+uT+deGAJ1FQZsyQbt6QHzrLjGc7DJaU137C6jeAQ9o6wF988
8e06Ra3Yf+fQs7HzmT9UfM8ZWQY0pK00AejNNy9kA2ZAOijRVFCY/VMg05ZugGlr
GugPn3RwEacqyqLRviS4nxTrJznLdMxmPU8cQoUfp/j7wqqCKv0Z3XE+Fazqppwk
H7gEKqx33VKagXOgMvEd7EqWiRQey/FhAFiOrjurJqVb4R4ZbaxxKTrzERz99w3u
aqoDvSbXadpApFbVx2/whWbFdQnB8jNG34KoabiDBA2wpxQ1Sv0iiSv/CTo9nqXb
1V91pgW28IBYDSJ79vYwlvc1LRKHJQyOTVKoWZEaQjtsJ9AsJ48DDG+IwrmTkCyV
jIj7muFSMKzr0WoAYTazZEUz/uDHuryejBVZ+QDQ3OWqexJrQGwZDddWeUnSIKw3
VZodDTqnJGwf9lad7L++i9hhpBYeDv5QCk3nRIOCl8f5vDL/gqka3sDDBe8ZKGtA
KGQbv7syOv8vZkiQFK2GWsq4BHCyJ6mC718AAW5gSPTKofclW3ShN2bDmuVIrVs/
CHqNOliAaclRG3OnOBSy2JwoNCXUP5gRIiFB8L6/YTiMYCjVjmaEe1PBF6ub7o9F
6NyCkoy0uNbGQEy+j/dm7iueT/8+SUPFPwO2y/CuTyf7L7VZifJsjL8EZ76O6iUe
DyY33mVALoahcts+dqvhnFlcwkb19OxLMopXM9FgGGMuTa7fdB+SwA+Vss8gbjHb
GngYMn9jXfqgh7H+ya5r6lGQ3Lk4WckSmNp1u0/Vamv3JjJRB/fdPA9+WY1TYpAa
jknFOBoimWp9u67Y4VZpy0nBK61LKj3vOGCdpoOifsQGKdQb2DFtxXvttJV/jS7V
WHCuwADoMpSO4CscYGgfU99p7z/67TtSWrc46bY4cYnFrqTiJ3BXeB5/+7bG5dCO
O0f5vzZz7xKnMunfZIgM49y9PPQNPOiR3Vh6rGR3Q0FJJqB0M6LZqaLnqHAcMcMD
/Jbu3O66MV9nyI2jL8Ebn3IR2OnZ1BJJJQiTc39CrAaq511nns1+oA655X4fkrcX
FW6AC3QYriZff1ac1QiJRMAv3xIV64FM23fjDflz7MjGlxoOlVwEt6Ogw71qRgBY
/5BmuC9RsPRbtPcJyWBnKK2cy2l+KnvcTn2856gfhXC5IkmYg/dQveyBykr8viBQ
+Eie5cWk69uBn+LXkop+zSmvwYfuHfpMHKkx2LZgPBdiVUbuqyxuLhKTE/RvIBx/
l+F6qxUTYHjNWybCCwCG5D+tpZGwniyMPnexG53mBXgdUj8r4hOH0+8PmR5T5wlE
SrLuRJ769YNc8jd9S6tqOO0nKMn5nsGN3AqsFfp6vQEsXrH4Co3Q0ujwiB5LK/tB
yRehwlyGZuu3KdVPkICUpdOiVF4XZt4NDh1CYdiKkElMMJCBaCmGq16xoPbnjExW
wI2vcI8AfUSKBCu9IMrhYReyBk9W1l8POCnSoIgUcpFejyZYUHIZXZDLbFpXJ1Fi
Meeg43oIXt9BABzizdmT6DiCuDghON47tC9LwCdBTCuDzVxkIQnnV3XAMJtHUmvm
36VF8eJMcRKfRwxhOFZJD3L0kVYIPa0hvnacCFqfBweVTV7SSXXVLEqxq+MpdOjo
p0JNGQ3CynGQQuzvzyo0Nuv/iFoJzBYDRwIHg0o6q9WFY2bOGn5acQQ2D8VRA8rA
SjYTmFMut+cVS29nKPl5F4qz8lFcCkysvg1Z5BosBmc8q1z9IGriMVyr3unA/BWl
YRiP3/IlkRsyQXpv/ngxAfVprLkrmvI+K/0afcWGUBU/MZ2yJu58ckwS14aJKNvn
vFVAl/sHCtGkBiOfjPyrmAAOcpU228w0hKGASk6j6CK7DQFbIBU+SjZTqjYDNXv6
gWQTPwMMBSfWKOHktqx8SsbAPJ23Wl9x8qrQC5IumpE/meK8SE5HBnkwVXgW6A+/
qbZ+psWjyu664GRE1TWDplztm+w+wIjBV0N0GJzhgC4qlfwvZWTY/hJM1vWpLEmQ
RiItc86cLmeoBntC4U/3GlQ1CGdrpOcV+SX3ltnALtA4AlZ3GcEnhjGcgVmHw/xc
1LKIdknULgbaOooj0rwxF8zKXc0Iic+SxForXuZhK5cbGgBGksxO534bdU3/DcoP
58hR1L6ya0JlQw693nLr/e23Y5O4M+jIgoSSyCf8ss1xAw3FwmEKi1GCQijEhhPX
FxGCG6/qEQOmlZnyToaOTYkUaai11iQVzOVFo5Z55BjvjOwWrxovlfh34MgJP9ej
W4y9Hm4+CF/LynE9y5xFAPHIkeW+/yvoD0LWgfVPcPEGfMPaQgEAOr7m87jbiGFB
A6aeVQsabAyLvl03CgN5LSlKMRVPAmk/6a48+5scAw8JiVb9zxzEJTL93vC0Xqok
4u+Jz6zWVeKeMdez/+uXZdVB47VDqqSwbNFnyZW14adL4VeDzJFdPKJhIFlXWE+M
3/VUKMoLxaRlOVPlcZGxtTn1Rv86aBoawWe4K2d3V9vkfKqqbpn4LETiID43nWC6
d2H5jYCNJ4QqoBPrBPL9CHKsX55rqh63d2oYDwegzZvXga3VikXazOYf7c4q4iv1
lk4j5s0VY8uqArVPwZ/1qepPhXcz2UZhbBlf86AhFFYrdh31oVBr4dNuxdK+s6MO
lx6FSfCH8XF52S+kx4r/iIhM7iKXMZCuVShC7wlRrACucTinES6DOdd1wBiCvuPI
Jv8l50vvsENL2QxYeOcsM4YE/DN27Z7HiVnJIxKCSwtiIyNzFd026LAww0M8qbMB
91UkGQrtRAJBpqrlfOQwzHG7OcISeRfIbpzLXMW0o5PhLf803N7Hm7iK2I/ywLgl
WG+1tFAbmU6Qzcb+X0kpZPNFOJEW5Y4uMhn5IhqRjoQNIrxHEQV4R1pfTT9h8Rn/
Lc6vPmZCC1nTwECzs+T+ajcO3nz4SayjS1sU2z7FlfBTwMHLza/tRBZR1iJ89K4B
6K1ttSsI9DV1pMjQr0TwL5TnpfiixGJYnjNyEegZAhza7Fk4on0pk/AeaOaoR+1D
PC0AGQQOob0csDwImrgkZ/5Lx5UvLRe+QU/7oiCdwYpz/3uVH9gWm4rffgGc3NaD
kkM7OKnpU1poDTSswGl31yQxKna02JtjwXIhcGq/0s9C/V24RvJJwUivwuznzuOs
z4drVOyErM+gdMJN3SZ9XRZgk+C42i8icTUd206BZw5lkz3kjGu3C2ZtqsQKfsQD
AVgqhYFwqh2JiiF4EORs4XcJSDX6ZZSFkAl6Acq541rDBXXD1ProJnoQjoOqenXM
i2tNgM5GrIel+0IVV98NVN7tQRgYAtxdbWSK0mbkoz6Co6G/1xgGo4lxoKFQwWcR
9aSsz5s10iY2If2oennOHRrBgQ5k+3qbXYIp1xwSI88wGDUtcjljCR4VV0Sii55J
vNzR5/YYs4ksHAD5OgoYBQ2z0kpjqZSeqgFpIu6GovNXJ6iHeGMMwkTH2NvAugCx
nWLN1hBRLymzSTP2BI3MxuHtdiWi9TUM9/mdiTA46Pi7NIpjOcN0nyMcRNUXANEj
uqpCb9Ev8pFcDdqUHfM1MYwVsbADnBfmAPqYXrGnkKWxchCCaeMuqZYQFRr9QzTP
0OK+pS9bytzw95LhFkySBG0hYy5rAdrCfY94NOdZDBn8vfj6DlzRFLWBBmhD2/sF
ReqFXF5nQVWaEXvQbeRstFombSAM3ArUr/YzdTfb2PAgcMTOk9HP38/rbV8iXe2x
+rgqMHuNS028nsO5ZqxCL2Sie1+5Ctsho/RDgoEaV6ryXkrOXIHTUIuKQjrYUItD
y8TdQX6l/yAR2PvbvBuuRw0BB6GIzHNUIvBWTGuI05Lbvxr7J9KPXzrXaiHnBw05
qang7RPKmv4BG3tb3eKFQrBO/EVkq5+w7WkVv6NwijPxv9duk10ocsqp9P/KkNUJ
ZE5XprPrvu/2yezK3gKumpYdh3YSkvBPhdT/8vhBVXgEqzBeRsXWK339OrtSNPHb
jvvXf5IZRxHWXkQ10ZoYEZlCUT1LXIuIObDGDyNkKezY3PQ1JHvlpoDyFh+PoX1u
D+Ro1W5OQUIJnmd2t6GCOD0PnwdW3dAX7VOqfYO7VbYLqAp/Pmm67BN+QWj0y8uL
yLuVuzzJf2qmsX3H1sDI1Ahnl8P7x4I/1qCe9Ur7WkKT6dBEDKaa89qsxEAnu26A
kKCdj+/laaCxlN9R9MCsZ3PJPoSjDxcx0Q2D1QI4GtGx3iWM2Ol2Dm94V8mI0FHs
RJWYc+MYg7gdzV4TT0CKliWhABQZPIfBYo/pfA+nP7rKZ4zdwlgjXW4mpNR/BHF7
BO379bQco88NkQ+NutNnUmtBJwOn9+V36hT0w9SVNlzgchd8gWcN7k9px2l0Pv7j
qV8MQvrPO7plwUXq5I92FFi70tHJVEld19Ur/tJMP8NZfwRjwQ0ox0gcKNBWcB+f
40d9EHwHlBsNf5u8+NePkSwIycZhZm6H22dc0UW/0Id/wUnRaeVuVRBFe7vaAJ4/
XLbT1tZC6uXYDjMuldAO6d/d3Nz7f+HrC3NnLj3+etzGOSk3ZvuAx+cj6K3QMSIN
UYcmWIsq+roI7GoDfJt9iypSc+mLshXGz71vs7fb+iJJdKgs0/OSIvL20gMdi3WN
P9bk0PwbB/JMD+DoMtFu4jWl8ELx8NLknkH+IdMUFAXe56Lj/VpcTNROKdeS2zBs
/bFK5a65X9d5wvUgx6jCCyB6kAQspW4xcZ49CJ/b+nnLC9MbGH++lSF+47nFpKpM
iqAFshj4NZTsRgUgted9rgBVBonXCbJ/dX2USafcY64MbprwtSp75XqT8iX/wBTD
p4U4A7rtmx+D28zcM1BvQy1rwbGHZvIdN4xyWMso3yMSiUet+FDRz1y1EBQ6zfGK
h0xQaOJZYsjd4rgD0/rjh4Hhxt+j95+KD+u6SNwpeQ9+WcPcEanDjBKYF9b/acvC
mmzmnbPh3dCs6m+2B9u46DrK1nkY2poZVidDnvoIS4LIyOc4pdR560IY4fzWSQTe
83fhqNyo7xE6oS6AeRg8BdlpM2n6ftoxwE7f0kagdnNdZiMe0+wH2V9VHK5KJThh
Ija0Hyuhv+euYrWokdNdb+q541C9R3teGwn2b0g2rky8vmfoYhEEXBHB063VAAcy
yZtercLCungH25m3nbQiwa5DaDnRQrXUU3BBA6T+T2AM7gTxXO9hmAvxjf3tHTmL
jKrXCHi+8NEJ1yUekeGwSvuUIQ15NWYS8GJkmBE4F5Q1171mp6fA9t8LjK3kaC+z
ey9BLJvKQeJWzQlJeVBD/IVTUVWGdzrj9B3GHSsxS0cx086et/wX5AQFbwQqvQ1t
eg7YepHkBWN5bgCwkexk/+4R/+fEJEClFTAuSJ9ZxYPYe4FHdQQMTcM+wD3mQWQ8
9O2uMN+ApbJfZ1eGaaykURlambr9jAeIbw9zBc3njfFcGMSnFXIZXU4iR3kxGHmO
E1vCvPveYPIQieZOcW5G7A07TByc/A9b25ZiculC6m3wY1J76bxpJO0qwCdcJeyA
aymTSgmHSXDVA1GmQcO//52nJaliv+Rgbg1Pg+2EVPIBgXEwmRssrs5PljsPyOZR
V8KwIEkRZ2OKocSwJLkZpuRNc0uG8IYlaqUywJx70OdjgBHg5iIs7oeE6NE2t7fm
giadfo8uyap5JIuXV8whMzreuQ+pV9OXae7N25lfxIhojhnOKP9Wxxp43a/x57q/
+I6JpWZaxQDr5zeHgmUcAAnBkV2Zw1Zy2yEqChahAYKPECo3b8S7V6R7gUG0sjT9
WHVYni1jX/SHnQ61NWrtmnDZmjtTG1PSDHyUhPJ9zAnmlY1OLbay2QRMJkea1X9c
AfYZ/OEESCiJ0g4Xv5cMn23+kgJwh3qrn+X6oOeBdlWvwfHygZI00Gcx2+7YWcsv
EQRdBAU+8a6FLQjPMb9pJ60VrojIKFCp0ai7UaO9T6d8/fjCSZMQx9QHWCkF0zLa
z5f+9OhRNLrarFaqUwH2qu6PokEvsbxj3pFTn2iRGnitxhn7yU8svzwk1RXOU6rM
O7P2abQ1HREKSzNHvg7NkGz+19g86AiaJdzH1we7zW2b8+ckTVxUbMK+MI1CU59H
kQRySSRxgUui1XZKCvHg6uxRTsuRvBynPuPIAgIIG65syGI3M9HWS9xUFjvdxROo
hOubBzsZgvkvtLurwXlLJrEA/L/7gCxn5qTjtB71ns/06w3VshWZ/EbxaPpgwypQ
97xhuvhUUYUORVbiYxtElD7u5kjh9NeRcpLfEWvLvIdxXlSqUJ/Wx5RXvySwdbSH
DFCP/pshI4/Mr2TELn8CM+rG7mFiDjzdIo5bppLeZWZjIkxFPIy+zKLNNwb21kyj
AZcO0nv06FMUsy9mM+UpL7pzyoODH2ux1scBopmezp6vBf9P7IZk0XhAIVrEuhsQ
gf7zP3UVvbF8Ed4yPX1nO1Y67mbdKJEHq06+o/I/Gzra80X/f3QtueG9ePeoFG7x
m1VhjBmp62JuuhTlKAA23lCLONNJQAkKoCWWunbWQlxsh6RzRTuCgxyDx+bk1KMP
Bg0keky/liBuZFGFoko1tvt7jZfOXkAPKh4Dy3kYnjGP83VnUZrwiSZPoqKK1e0K
tPN3odHywe56SArcI1K7VbmxQgkLme3oAZn7FgPUhONxPt9WVOkbWSXlC2iuf47x
kKM0OMeBH1nD0pKKrMYXXpu1MZZJ9pfmtWNVDZc4c4tfo4rj1XfZBMOEUlpQzkNj
CFoerDOt+gW+7Uho4+MW5Ver5IL8FVV+jff2NTZxwvupR/DeRI0UzcSnYbNHp1Md
fRmo+xldI8BV8AxFGoJietyZhNaQ5/4fPgzY3S2VftWi7eiaVDGIqJzVhnAiwFzv
gDXb5eZR5PSWis4c70Ryf2/Mccos8ufWF6xcsE1iYtYf+6cQW9ubyPZe7b1w/soz
7y8aEbuEo5Id+LcNwwGiSoBvfE4gG3lqOapDJbnuHVb518B522YbfdHdg3darSEU
G5MpCUenoQnD7iDrluXu5h4du0Dshn8xkiJ8SUGTrZPEHxPfE4vsiG6tX/qwK/Tb
L89iu/jZ0TxMSMqcmiV6LrpPDaKbk/W9XcXXQSFlvect83i8RJEIju48HS3PGuk+
rrV9+Uaaz5ZLL/CNWGD/onJ778PABFLkXylO3UowupPXbW6AuBV7gnu/FVaurhqN
zGjMsjusel2zqWaINtN0NyAibu8lh04w+SEzFRbQKMDcqd6T3IGIysKr8QdRWAD0
2IFsnyc6ZeItetS6JKc9K9DHfd7Udy7Mr6+ToHBg+UtzqbmrEiGJjZbBZjVt/ix5
b7d/OLSp6kItihOH9IcY8xOpowsL2YDNLjrArUdD0hX+qDJAVaC0dmsvrZsFq2yT
+ciJQJBlRicmOs2NqWwG7rtP1OuK7V/QDz7k5IRmDgRRNTB1Goy+REyaDiqpMemE
qYgGQNIPsksfzfLDXiVOF/u3zu5QJjbZm1Lw4nDgTvXZtjaxuSkqut4tlSQEFOi1
EqVimwoL7TXUwHRTYY+fqlFdlVjb+4sgNCbsk+QtvMkXmNLhW1gHvjB63+eXMiZV
gII6ZgTZCIxaLa3GW4D02IGHHlCJzI/vUDYRvXyrCgQayV8xxPXylCbeee2k6PEi
byyi4xSTczQX/MjxlzrfNL1ZAtOy6fC9UWZA8Fpe7gmogN4LVDmOPXATWc7U0+6Q
3flkYVOZQ6x62jpotHauQoFx4T/l3Fl+cgKpFgX0XY4FyniCC/YVNwNGJtWjqUvu
rClJUS3Xyl9Tkz5MJcTiMTmvZBNE3B484WQjL6HV5zUDUfI4URWXcki+6PuTmaSN
XJhdujgpOqUkluZdsGj1DVl1phLoZxc8f8gW5ODDGpKsJNuh9qu11rUg35qsskt5
iHr0cle8PKPDRfaOy32nh4JixSl8AkRIdzHaHKFbS8K9hUgQUTadrkiQNkjTbACS
sutHxJkjISUacN0qtHa52g5ohe+tjo1ZVHcQtGk9frT+UD5enTClO2p91KkJqdq/
sD6vNALRrme1vKlh2uwdFTIXrjIkHPqwEgIMIDTJ0teDQaN94RDHiak0Q8Vy7fmE
n/GmqpgzwycPGPBzZXDCulGJjZTIq0UlCpddqxrtqt2riNcpKAopU2s00g8CreAM
Pjaa5TECXM2pXPBUyQcXlfqDW+O9BElNShZUDYRSp4xf/4KACXrBO4SDDBgOKaXF
sadpL33J0L+NAWgTVMaOeIu/oX0MinH+PgxAQ0LZbrEeaofVJeqpic/hGuPGCTuW
374iwIwDIl8W1GzbQSyiMQpcdZ6+otWWVw1EBaCGdvjYiBjzTB2yOT2fxDvRvjHW
3o7mPwIjxZVs+VtUUHC1x7VmQUdZapjznxZUNQfbVkMJpH6MAGZ6ozStfh+r1vti
fBvQasMyp49yBJjHVUZnUajZ2GLtJQaUtODqgWhALaO+VyHC/EIGpzqj+SPlwQ/L
aJiqIIc8ORNiB4K7wo14MM0kmvBpRk/E+K4vtv/ZUWTDBL+3wqJLefXaktqlDgZ1
MQKttDqOTWhlF0TFhIEsBDDCcoPsC8nC+mMZtV36SXG1g5qoHcoN98vXoKgdkBGY
JC94G8ryoNIIrZamz0FkgT6muLd1Rr3ud5/oxGoBf3e5bfgB6OAKu+RvKRQSjMKk
WX7wgprsfT0xKg686E11HNHXDHcuHLwPxdKTl7ZMuWLKVpm5QLKIg+wzOcTWLx40
Y6aYVgrBqCZnij7SA76C/DDgSWu3XXw30DZKbHeJuNIf35dq+iFMIPOKqHCBpOSG
xhzNmkZHd/UOZg2+OUwAoyLNX8VeuBQ7o13TfivgBvqicQrOCXDN1awcxjUqxXk8
mhaTaGoZEMaPX7fmsUWbw20EFX6B2ovJGjCm0/70HADdFd9ISSa8pQxZSMscHnzp
eHwg6SMJbk8ig+iM6huh2JhzzrHaQeeolQWMQ1XjHf5MINjN4ze+zE5Rjt+lpECE
XJrTW8UstE5tCH9xbUGo+jGQS6cqo54S3aijzAlKxs4OvMTI3IKhKIQ8DYgJYQaC
vZ6wXa1L07ku90veAmuj5Abdn8CVbzBjrPgqYr0P7zuo4spRGxAkB6X2r252tjum
JqwpnZTnLUuMCtPL3ZQ3xKQ419/uVlaZC+zxa7kNoU77hUO3xfgaLSkH2oyHj34a
vOHtbZ5QfKgRGCBI15Jm5Mre4xfDamVjeHYJuvsgKEnBCeP1NuBYNul6fwaJo33o
y97M98WCkWiEER/elEI3kOWzXif0BbFDRwmWC4e7HbPJ0ABOYmH0vC1dVxLHnlnq
Qgln9noCeHfiZ4HAB1aty6srrU+4ln/Vu6gktYttmtfXeCUV2VUqUgQhJZY2AxCD
pT6bNkGKxI49H2QdKMihzDlKY4ZchF0+Lnuyq3bNvU7L1Ek99MS1cWUI9bOd50KD
NuHmLy0IrQAeT9DcGE4S7D3wwSbv4NTM9vuWnryuVFU0EmMsrBlUMxDKO6tPOMQp
xGjX4MXRC2W+KTYtTtbxxUuve3teP5oI0zD8hMHArLxbkK7xwcpvL1rPuhBJNsZl
6EXFhz+HZ07u2T0HuIcqeV5WjEmR0hrNodHGK9WuebXdx7JeUgx1oEre7BlMow2K
TKhUAzRFNWdseUKWHlfvgJ6MZhn7qNuGWJEijBejKPgCIYsBFKBSNr6/FDyq6Ar+
v1cOMFUxRy6g0jXVmuyQgZn8OGkgFK+0ploMo8JS6p5Ljdpj4vqCaRWGLZ7V2mb8
wBlQVVm6mz1rX5+55A0bRIXAXHzREhpA1qf6IZv5G35ZlP7zqg+qzWl2s0fS09yU
XF421Q3n+d6Xiw3NiSi9V0Etsq6LHykBtGFHxYeiBdjKJ307u/SE0imecm7rgouh
Q7v5SQfjD+Dgh7sAiBrutwhl+s/3r0eF6a2HXPtTOo1PZeVmLqDzBxBdXecqeeZu
ddT0MLo4mXb8xQPH6VDmdXMV3riCC7xXxOeFwMznS/cRVFLOQzMA5TXgqED5iD3X
SJa/qjPOnRLMZcgPSzdg8VRpZGmaqcREVyyS8bAMepAEvi9AX0ukXuH7iCsmhB8W
/wMmjRKv0VLa1hdrrr0otuSueGP+qeH3gL3u8isubrYq4ie5YTaIqPhqSK0l/hsb
7CZy9LRD4HrI99BZbrEcLm4J9B3Qg+Pue2FiCI5rQcAJ2eeoUfXya3G/XyOkeCht
vNxuv3gWw2HQJePjbvbj6Tg4JQFZqYIZ8FE7lA/lloqgJCvwa8iAbozAO+mhU7kN
KGFPPTKYN1+EY8alcC2YMwCFf5z/O4RtUHADvYmIDWAGXhWyKSnNmoPIeth9vxM9
WjT7ah0t7/xnqh1opJDslNO5TAkfo0xRXErkEym8old9TEXSSv+Ups3k7rvDwEKN
N2l8yEJ13wLpymVt++QRKb/2ZPcvas7A6C7mcBxvXja5uIESj2l+q4tq6u0iHmIA
++3Y1tVwf7nNJBlf4+HUVf62JRrbOjV5yNakRzggLAGgmHs1D3EPV9R5Na42VzIt
EVM1zeNsgX501w8sL/rebWc8KaSPAVoTBKXu7PTm1wN9ITSlKGJOR9mqT6mESY2T
/1J1NQqnvI59/+vkkr3AAuNe5ZVupuOoHE0rZaC7rB17N1gC4q8CUXZolrs9R0Ws
g67qxLxniqVV2b28aeHuvENOoWOYCqy6HTW0aVj7yiGW0pIQHiWIAXKcjK2nviK9
js4+axTw9JOtUx7rYA8ym9EDfT8f8Mm4dY4UQ5DXTh+UMZbi6B1sbVoFeLtFGMmG
p/sYp+avOBwaPHujcWxdokWBRVB8IsZLHLMGbNMcQrRkB1kJhVyAeiBUBW53rTbY
75J+CH4UxeloVbqXGfGoW8Ke3B9A0d+sXL627Bk2IBmHBCLHD8LMb8mHkSnYqCjK
yrjFKS2DK2xaO52qGO5/ayMhHQnmltDMoEuixhN+2Cpp5H6Y7ifUccZ80FgtiPq3
ou2nIYcxSUGvxOw9M/vcnVLy2d83N7T/Of6VP6W8rTsz5gy4m7BcSJTeuU0LgU/j
N2BxuLlPUAljjhfiK3Bc7hKBfWLc4BZ5KirS+hoTpVOt5NJFlAlTzOJ8OMAKL2zk
TsRN2c2hCimVAMDcSPPAp2Gi9xcOfDfbZ3ezZSX6C8kXOY74RWYe7LXRv05fqgum
blf+OWqwje5dR6FsPYMmgqcvmfoibJvZoUmjireM/Vbqfjeahe31WpttQMTszLOl
0MjN69ejZ+snOmozEIP49klz3Qpuc/TROqovyFQBKjbGbcuH+PFJela6gnhCYoPz
CRSyP15fRZFcau6aum2kJZ3TLxmbxGOCgAvHZ3HqTDtZNe+ydGbJLFWh5vJXYnJF
7JoXaaTsbg+G7yni3VtkQFfNcXN0keOCb/i34msj1Pt26+/DqnWbkKcEnr3ov75T
QsQiHIrEFN17+8P9Ude6b6UqY3mRJ17CikVPLjiAyy3mVeGlMOXohV54YbythOxG
V6dKy0VKMNiAmWRq9npTYSlhQEvEjaAsT1S1wB+q2auceuCFrdSjDRlsAx6MJE1w
4/cUd7+js1/Cy9+hf8icaw2s+XVhGaKULVQ7NEfbgqh0/jfyLOYIagSv1BpvagG7
0I4szCCnc+tfRYXU5IkPdPfR15PBFYeQMMKtglrpkFWvQWqNdAQilInZyhqf2W8P
vl2846kGSXCHeBlZPlCJ1V+JvWmc8yqib5z8/HO2xvE85+c2g3RRW0izwLw+cem+
woUiJ4H3hoEuIhzhrsslJd3l/5CWfQ8UJ/JpW6nkinVd4hgor8LWCtTKuyBrLn65
yfGodslyd/ptAPSB2PbdcOTgcGOJ+dUfiIveLjqMsnZt4352AtW2ym8M5J3BmldW
hdHzGYk29PpBXdJVdddsGMH/pyz3ZIaX+GEXqD+Q4RD7M+8a5l91PZzMKYYJ6TJr
1aBMTJ73ASBqT8d851Vixqa9Je48VgGVXaRXY88k9NHfZq00I8fVfOvzng4Pb4sB
2CGuXtsIpsRv4dme/ZdEUg+GXmLxzSyDWkWf++EgmBxwegGimBhZmw4SL6X0oE02
XoUYwgSRPblj5U0XPiy2Y5aiYl6Zuh4NLQ8HWrblA18T8w2ZUD2wfyD2rAjezyRj
/qFYw9+mkaUhGjxxUOnI0IEMo+R5xqCrBazOE2xufl0ZM3wjdlKAAGVRppoHbiNI
PUObM34S+WtUMa5/l4I8DGyv5De3vkLCteFB8NCuZi72bxJIjODq9T7lZmsaDvPU
xy9EdfAs+CaQGHNZRgw4PHz7pd9ynmfWiqBMVS5vehsesjRVisrVuWwJP+uazDBM
sarbEbQ6B/CeHNs02Gd0/IjkxUBHFEq0c/pLkQTrdpAesLe/Xl/+IvNMWbIrFnD0
RGtm23auTRRocCm9NyqIMNhPovl6FXpS445r+MdHpROoxKhowB8R177CTZZGfmYn
VFgt+Y8HDY3VZUqM3g1albxmI64aUlP0pJiuSaWl17x0CSiXhWjtFPcVLkV6+z0D
LvH+TH77ZWIrHIpB+u9umptatDexXe8QqrRBTgsniBr735bMnF9BHcQn+ihlhgsX
wE6HRZxCRULQ8SYovEwL2E54EK5q88DbH6XeiodMIAolplEKCO6VrELWJzNAMNni
h0ek+JFf0k4yjqOB1Bg4DKzwuraGk2WsFmNXLzvjD/t0eKCvhDae6ZT1sWpdqDU4
OB9C4yi8bjRWWeuBn4P6aEoQIbab7WOjetwcJBxFX8mBue9D1GJh2/9biHq9+IHD
CkwF0MFJV03BmW2DB6oECBcVh4ipqK8wsaIueJMltbojZImWuA4cELD0tPSuq7Oj
EFePXexMEJWRLVBdbj3U1FDUQJ6Md83ZuYOuMIkxxLX/+Y8I6fQsXypK6TceJJNB
O0V0p7wbRHnXCJxwQAN9iYal3hUCxBPA7xEGjMrXkzFvM36NTrl3ssWrXEGoXWzD
uLzOGEmHZBI3s8GLs4wV85AAySf2PCoLxQ2xI09t5d92IWA2TSYnSBYkPUXQw2mS
5h+XUQ9tnEUMClOOHlCOMpoqvLCQNsFE1Lleejc2ZJ+f48xwEceKl7N3vxtca54G
1BHRPqbGU+LCh83tnLUtQ+OoJXnLWFEHfPg2YYW9eR5//W6i8eRzJwJOxdW6cXe6
Y0iBkUaY3cHgQGvo0MncQDI0vfUQ30BvT87W2iX0c0NdlDjCtJaeHbwUqLcz2GzN
+WqeMch710yw5zsQfbubb22C18plLOpSsR9735yRNYz5n1IDRMqQoUup3M62lua9
fmzUlXjzZZDtFgDRMn3JMBbzryKECiSiBavGYFMIuATU6fIdEepcjgIlgbGI20Mt
g1Hlk/T0vO1fDFmZouQJoJE07CEydtm0fhpLgzYu1IIY3pqYDW8DJPY2yDqup8Kg
ddTUXStOO6cMTah1w5nCePnPmZOF1bbTVnB0PP/l1YFI538DMmoSz4SxaB5emGWu
IcZ9RoqljihBLDzIv6HSXxAuvayEGXhghdxtyGQoTYhfl3nRxXvxd/1hNEw/2JDf
jMf/bS/4Q4kK9e0WOVq4TbtHGfyirLqIYaDntWOYCwWdWZRzUJfuDpuWmttqzHAx
nxIi5+60VHnRD8CN6UlFmIC6g/MWzdWoqQj0fts2U0fnkTaUC6Y8JYK1UT1F3XVo
cKSMfl1JE4BuvEzvuhFLIukekwXRiXt7Jh7g5CZ8MQUKHJK5dPfbO0ridIll6YdH
9M64c+/Hhy109sHwEOVPdGJw2XO8XJeJUBOn2OC1xel0POQdK08a4s8IEdPz63yb
BlhYuoLW6Mfkanw1iZISRUzSsTr5Q+2Hi9pWdjgBTCm++hwcTHABd/CgBUaCDLWS
iqy+GHmmU5rUklXjmYKDLgu6hamTdzDCpzre8ctFQtQlqEhYjiqp12N968eHSXjI
L80gPxcNHMo4ZDgYW6dSPJPF1I6oKuTB0sZ82lrXy2INCoulSlgSv8lmSMJYjSaC
Vwj8kHq3dW/dRtwdeNLHLbr9ECjHRl2M2vM4sgVjFcItSYGb2CfXxUDCOc0OMwkA
SI3PGpNyNLPUTGl4SeGtJ+hYweLswSNRbDH7Yv3lqYjeebvaZLYRFYhr7OSlx1Xd
c4l4isidIYVABhq+qEuqQ7uOVtArPB7Xo//SCsY0F8Ucfg6P/Sz/8YJ9zW0rne6Z
misHdoOnZiJOfwQ9JwcWFXfaS/bYlVb6/FrMPGkrp4rbNqlbvp+S86hhxh/XruXm
HKQDgdun5QwWkYxc+j5AuFSUA+C2+d5fIxO+Sg5Y/xq2Xc+qKB6p6/0q7ofj3D8u
YbYJiXy7JKtvBAGXZJRgShsQfKwpu3qI4gOEIkMP+r63GsUCaDFc0B5sKY2al6ls
fQ+ufwI2wEM+w17aOHnjwjtxH7pY3NPnQZWeW5qRoKCwyhGGyXVhzysZRy0l42Eu
saWrKEKxrS3b/HXsLBlNzqMV2yE1uycmdmRjCFCNuX4vxf3hWs0m6W6O5/CKZZoe
YA430BfiIZj6i6QXZqp1U4VPjQMfeBaeKlcgJZfWauUe7p2agOgMNFT/I9g/GacN
l19ZRVox3Auxe+d/IuG/AR/RcAjFacbTnGyp4F6KL7d3oSYXGn+aXrnjfSyfCukv
845G7AwzFd5bDf3UEU6EDEMMOxmOKS7CwjONXHrncLpGlkgwoJeVLqW4jEijFdJB
Jg9bpJSEhd+vbvcS5AMMoyjht/cx0l4ulY8TQyW0d77bYp5ZSHsXTqxt9FSzgCql
BjofQjA/UJdcfA4if4agR1Lk++dx7Ixg/b1ML8tKJRmTjSXlxGri9EU8Ck8Wzayy
Ihf4HS2NbhJ7DgniCDLl/ZFJugejpANHqljlY0UKjWMekbLziCeUeam1kUtHLO8+
nP/3+B2e5gf2A+nNpVOVyITHLDK/mD3jX8qceNCkPJ/ChTiCD789nAPWdlUP2Bux
/jZ2rTdRaqMWPvl2sSrUYjM1T2a1rrKTH/2cQHo3V7NOGZ/YUq1XK5LjEBzjGw8Y
jhHtdiEmVhClMfwFdFcOb0WyhwBNfcIRx9Bgm1nDPl/Mcgvsu5JKeYuWPV7VP6yO
s5y/NFRcA26ALlt0gdpPFwsS9iTtqWhn4EZAaf44fKvov4dOwK7LvXh+hJt5R3w7
QXkUO+TfoN76oNXZSLUDX4bIwSzPaHXsW+RgeASLvF2bAIK87NN7FHm73pAyTtgK
WI1zziBKFMfZTQ1GydIZUUW1/RxfPhsTTCdskGozXbuKenY88lspasSEW/A1mIGM
+SAnqGPdwUfKhmPQYlYosGMJJTawodsZTFOw/k3OuNAYGz0Z31DDOM61hD7coftP
gHmD//Smp2MhlaqGVhV2xojCJWKLCxdcaVWs4MUVnNT8de0FjjjIAXtiOQW4lO2W
abKqyhUoezln4x8/vfzqLFS4R2nTmdUSwawfptteFGEMhEHegCB/WPtNxqIJaT8p
q+POei4EIkS0bOJOctAeROI6FjBaHBS9Qf+6mvkklHt0vjMqtrrDoTwy1FAkdSIp
RNzsHajexuz1swA562+/BmjJalQsZwGB2/V9oIIbVWKNoR/pT4JPyRttrRG0SVqN
xV4UOjyOSsNL32CmDVsD6KeS3RlB1dpPDTXGTjpLRBu0BCR3NZ/V4zm5l9HR1Jkb
TvbJoAtdxY06fWKY36xPA20kLSo3QhsGEHahGl/2mqCKX2o52/gl/tF3zlIXb3jq
wJqNBdG+FTvcUO00fzKeZH7y9zKVUYnM6Yr/uUJCC4JteGgMZ272bkkaqE8Z4Rya
EzeO7FzL99IJERQT0ZmVWLoBEA9ZVNHo86Dr7MlEFlwRwbIcKUEK0hb/fjbd/Ixv
G4OlOMwu5UV6gs8HoII2MvFijFp58huoUGkQPllf12x+Q4cpSzSL18EsAxt9/qnU
YMU1DVXEiEumzefbRq7HGJ6ybgIyXKD51W1+nG0uPLYzax56XR+kW7FmZEBgg+6F
4m81i8pQ9YLjBBRSd9acXhKRlPxj1Pqg12gqctSxL+NdCiaibtAoU5tAc7icmIva
vu9e80qO5/TU5Yc+JAPGnPgjaphGG68wLUJtNmKAxJt6xTV/3fgvGsytGw1AFDgr
Zx8RQ+pm9gWR6+keKRj40nSFOhnHq7q8dDnrkYGerPeiuLuf7UjUDeKVBI+9X8yv
FU8qwnfzlmEghtoXvWY+Y/umRHI3gMGHXX7oxk4B2tp4ykw8KQPzdJGZ/pzVSg3i
F6vmNCPIn/m8Tv6iL60FgBEFuiLrMNjNZ+HUOQv79ISsHuwH0scKIH5VIKI4ovWh
pFmeJh8w9bSC43WZfVaGMlubKpisCE11amfmaMqeVj6resugp6arGIdmPP6AzKFk
FNpyiaMG6wo7klbAcrKTGe3/QXshLaI/tgyQ1S4FqMCCx013wDSMWwJvrdjXsK1L
Dg2KeII5zAZPWTOsoScsHcdddCgW6FRK72PNrR3ER3FoZbI7KyhW2K20Tz9XoIIx
BfYClfG+p9XsX03SVO4Iifw/5AXxxRaaagl5R5RcSXZ2pTf92Gft+BtVrz7qRFGI
TPrE/DelTDUI0h4FdJRRHomlmCkfQcRFHX7NBf11Ufzygr4I9tQDS3UvAlDQ76Rr
c3rZ91oY2zDKgsMtbbQgPA2a0TitqNpG54NCUi3JCdnoW0rR8Jg4hCLIv4MqVFtq
IfWVT4Of76f/rKVwpZCypu0PF2ayeo2N4qMBwq2iO0ZFRfm/ez4nbmmqWEQIC/tk
fy1EJqf3ShccMp0eVRNYOZP6QHXDDWOpjYnjIOeOKLP04G8Pr6TohkZT+82ieTVJ
8+2jM5/3I1/r+qu2eb1fEjL6TH4Wpa0pIcwlZtDNcZQtLW1O0vQ/RN3coKQMXqmq
0gjy2bfMewkYFZ0TmtSAq1WgXewtQH/ALFgn1HYneOKsq/rhlHDhJO7TqE225WD6
r0JHeqEkZqSMa504kDGRAFF9o7l9bHdV/+1Qsc+RdPwxMLWL277H/E5vKfEcwgk/
YszblWW6HOkhuG5wI0llBdCdRBcnPSBLRfUxPOyswj/yFjwqF1p74g8Hmyd/280w
Q5zswsn5CxD/U+i4J+QChrs3IOq8oaYClvOAt+d8SYx2jr+4bgdvsmG84+oE14wA
pC3MWkAa0CpeBq8aZ4GupbnaGUx3+OnqRCmffx68PpfGfpur85jQWCL1LDEsRyLx
8X3AX7JR/s6SmQQ9hl+tw1CRZimPrMe7Fph1q1N+GRgJfjbrEvUJmnATtEi0sLkp
suh3uXhqh7ZfJVWG0E2vd8vD4zql3KZpUsx1lTOSQvbi6PapPYtA1rVX5cuvHVpb
nNaqfV4RS+9v0zmsY7LmEO0RCrZyDSxLGZAvyql8UOGfKS5/7U2lFqzUjOCpD8Nf
7Hhsoh0RJQhmlahAkx2f2XSFCCeX+KWgYZaQPgOekJEkFedfblHyWtlJSTnHnq+s
qpbPJxEqwOGaNo9BuU96MShpNRtQO9sjg9Bz1K5chkSbGHZOFL3iJ7XcvgzGDanP
XxWSLc3EQNnoABILY/umT0WurEWZ54J1g2DePVDZ+gYe17ccRuH2GpG5yVWA0F7b
btb5+JJmpRvOKOUYGsWAhrOhSkGdXIfgssmP06gOzK9LsfvdS6Ny1NITJwuCDv1+
MR9zEcRkHtlrZbh3C1IPtqI0d6+cUUsAm+Szafa3RoMhCdEeZZuNj9skLkCPYg8T
dIvI2A6nVgWcWow1P9JBZPVZilCSPXLw2b0e5akVHjNFQ+mlgcIJ7Be6kx7dDl1u
0yUP5d1nctmUQTcANeicOU3EHpxYf7vpGhEk+UceHYvGeG5I4wJutTJZE2C/sGUV
X+eKkTJMeuspYFPGQl+KKtOjISqdPxNzaCytd25Fb/m+9MRpYjvoSf2syaTTre7M
hu3JyDg5LK9kUres87/QpvWqtgmGTNW2ub1X7GD1AMGC6Jt5400CenlVty2w3XWY
FSryGP3ISgUQo5nOvpgBxpkSst7C1ZS2zNSkbA1SduMwrbOr3rroqcFROFiJ2HFD
vdqy1YPbkKjzVFeqhjtIlqFbPwFK8KbHWHxWIziANMMTUDBQ6vPkM4/O8uwtJtVy
Kh6i12daHgNcUc1F7KItRSazjmvzfAvzN7dKJxLc/stvJUbj/eY4IMIUpA6z2dKo
0k6sHmgRy2vNE9t3VQiJMZUSwikQKSbcH64Y7aVXxfdWqLalHeoAdmO/P1izCpZh
CKbaRaLkzstO6CQ/g2Oc9SFsTbfXH8SLUWNSMEhkx2VgUOiSqorh05fOua3ELreB
/XSsApJRtaRy/2bGnAGdXPmc03DAEQeO/SbomW/dGApLDuGmPGtB51tDDBa/6xgJ
bAlaysE6rGKFFNu7IFFfsZmdckMqFQtcJW2erUumLRJbYMcZLt0olaRNFIEWqti6
DGXIII5U4c5o1ecjJK7HcFLhZDEoP4vQBJ9ma3mbCIjgC612VQzGCNWrYCLMLl+m
TWQXBCpxity253EDuvOF3u4CmQVpyNC4U7vVrrkZtLoZatvwmWUJR/Mo5na1jxqn
swaTbUQHSEhF232cMhAURumFRhsRMF26+Fe3eUvfUcYz45/fYU0p+rnmuFPCsZlv
BkVmJEe2YI/uzDNraP7B8TzcX0tIvCZWBpfamy5bU12Q60Z00zIftfpTIcHxf4TD
ZEqT5v61sLX+6glGnsW3UJAEX4hfa8A3cGKS/6EjUcHejfrIh/FChiO9PizwVeuV
P5mnjNe5bEla0gSkkOzKABkldVnWaXOlCLQKIqxFC3IHD7D7BxX3/m3bPYGsIVi2
folNlLTJO6ZF5nGxBfnxHFUAkx3N4T/Kr4Dl0HGaDxKVpPQNijXLZ0/X5877cwNB
lPhiG/s/1IeyQT/uTxoGvmFlpyiIroB4hldSvg9it2nr5R6j3vInvDmNbF7PFMyG
WAvGMcYNjkpS0onSTLx9E8lsZdCnFPzekDKj7rd9blIHY87T/plqpKmz6sks/48g
eF0spSw2txBskdmjzWJz04pJ+yChR78UKucK36MYiVeqwUiHE7M1Hrw/oPTZOdvh
bqK5qBRln4nfxusw7XffJz7S3xt/8oe5w+QXmehRlcVx8UVCeFyjTjiejt6Thw/7
5y4yuzgwoKPStGAQpd6mrnoNGDnOj7lJPDAhGGIEYGI2596kN4lO4OUnWVwp9G9k
JyV+3ezrudbJPRpb8qUqgLsmfMm3NcS57YLss6zsm2SPJHDo1alrOUmHbSeMgyAr
2tsTOKbrDnrygI89HEq2X5ISVfZIrgxEg4Ij/QfcSfjEtfufhkiY2iuaGZ7iUpfO
a8rE8AUOuPcjVsJ5cDs68tnZCL4L2H6VC4SZ8/h+b+KuErPuBFRr9FCcRW44WLHg
Um8O+BUy+ckOsv61nDsvdJF4dmuU7XC2ltxRFZtsi5Q+xwkQ9K8Ef3GKydM8LOqN
w5thZMC5L2A43Z8t8zCPElIP4rFeAMP3j3o56R9CJhmYwR2HRCEN8PfZ6kDxrimK
Cby38CFCMchAnteemgJ1hND7HiB4CFpCUOiZ4IXCm71t4JSHhnfvLvFo2JXVaGeS
d9k63EFsyOej7CxLR+Tr+q0uzyu1xc7AywYH0CzTQ2Ip+SEUjWStxRe5ZBygpVzV
yzC7mUt6bKZKNFOqEIDuJnzpIRxUn50M2C06wUftpsTCh2PwuyD9CHBqMyuN/qb1
13vfs3GV5rd/WATKCDND2SwGdyfzEk3s/YDw1ErtJGJx8936HsidDNR0IwlX8RWZ
fxN2RKJmRySHff9ulePwSsFTtuxOs9tU3B0DD5JuTe9stw/kr7Z1D9Tmp1+wkVKt
LYlWjSz07kvsghvBrpR1uCiYUGae6N+5ZEoiqrMfOvkFI/6Ygopym2bV4eF8LHaY
W/2DTCnFzW6XS+D2qLKp9Ir86EptnlO/CV26OyqlW5adZc4F+HoT55EQt1/GBB5l
vkmt4S5ivj/FAu69zLs+25VCnS8mYu02KX+s4RnA7GCZsZqaaTyA2mauUvyJjXQC
R/5Gjy4Y8sX5QA+YcQnyfPZRPJZBSnETflz6XrozFLZKPd9PRxrvyw4hc5I2j4ce
9HCfMRrZaFWgjmkIEm/xo1RDhxQ4HdS+WaYsDWMphrsMDnfKEXgOa/akcnpZ9v9A
6zol1wA7iTsU2VdR+FfuiyuGc8FhsQjMxdN0yxIIsYHdz0+NUDdCYVPbazPxblsb
7P/6dCoAwmRtQrGDXN8ZwsRB2oilpKZhv52jCNEiAIeLhaZRnDnRc1lXCsXqB55Z
aOh/6YTW3kcTmrkKtxr4GcHkzEvBdh1GveabJ5hKPzmtuRsZmuHBxGYr9F1qJsqX
ujRv9nwXGY/Vw0I20nHDD6KP8r6zXPDsN8CDEE1+ioWOmyrggfzulBH6LtPKM++Z
iiMRPKDOwW9kNb8BLEs6yOj5oNgWSqf32FqZGMmWb1g4xl9MjneXiiZfBBoOD8ib
wVgg2gIQsEIOGRo5KvgKhuVtZ8oZDFQ6RcXQ98ZL5NCVCl2YPE36H6qjHsCW6tIJ
yzgyRJzISXeQhohRR5PACABc2yMr4CbyH9LF6i/ZjFOEZchygAdu1BgaJ7IT3ZFk
VHuiJC6OZGJnwnBZ9PvFHSYRdhcW3O2dt/g1PdCleBaVfoj/5mLTdr7ZYY3KVmyT
/HQKRd8q4th+huPFWnTSwGgd3wroR8bTtFKfq7Z2772DQHIEFnQe7Mx0BC06fiiI
Bhhq3wDO7+AJvK46yD5eCtoEcUkpP52t92Ie0D8MS9UhAg3X0ZHJru7ob+OZuh7s
v5s9Z9y66Vl/ZFN5z5exznqoM3yN0r0VlAjjX0R1FCK2DhFusF2pMcA9uPg/9Hj4
gAFkkHNm9wSMnZhdP6Qw9EcRTAVwQSn6GHUPY8orjBBwHYWjips9RFVEzbNO+vw6
YCquJRT8muZWsnu/4YGuCA75qQdnEfzgs/R8/EOaZXHOgL6QN/J5IW2gP1ABc4f7
oMY0+SL0S4GtgigOwO4TyklQr59h5PhBXCVEpWXvrn89xC1S3rx+J4LooI1VjcAX
U/H6jkPgRfdI3h71RtjX1XzDAbhwDVPnxR2wvcQUz1fdGuShq/K/mrrdgpewVbaf
jouhv9mhNVftDIoDbmcTtykQsbGsk18Q4PRgpG/ZryUZa3N/ix8YiOX7Nsn/35uw
92JU0roLzcQcOJtLUMaHNZDvC/uBthxK5yMa1cUaSsjtfCagbsPG4qnq8qiJ9Yk3
4ssHe4fy6GevVxPERL/TP/mLC9ULHc+vNQnxKKdPygPwCh+tdpmigcNmCNTCvYlf
Ocnb1lxrOnOZncAEpUxn7nTXiRrX8iAsdNHGWrgUaxlGcS/1KdNYQQLWulJrNLp9
+3a9188mnaK73LgaMqSL1HavVb+4zyxGXK+yOYc0fC9s/721pnjcmAwUoa7NDcb6
NOZZ9ju391b0/tiX5itYqRq1Mnc75Esl7NFy9V481BAxzshY7hzk51mZ2Y66P8KM
xTYgi40h/U02k+vaJFeHyZISHs9jsTRu9tHcPL6/9O4ASznyL04ADA4zADpLQDkn
6VbH3TiipCZae3Bl/3Q5BwOjvozVYEfAoNav9r1OXMaO/uYAuvfnAetg4ozXCQYm
p2vHN54qEwGkWSEknL+bnFkFEOBWzb61IM5kj2qXFYGpixPHUpqeBBc7Kc1XHr2+
XANyK9z58rr2W2WgtOZ5WijUOQKASizotkP2HGM9hukYofGARv+3wVezmUno7Gde
q6BgEOhGpSCrbpcugjdH/0h0pyMBdQpt/9pS/GsdDFJRmH6sOMmjEZ7cmF+Br0+u
9qZlR3bGPmKiH6steHGy2tj0AkcxyElLqxwuKq9eUKlhQazRaXRjAhpkkiX6JWD4
5V6KrIUobpPpejHNVRluO43KKFa0h81SD9IaLp6SL+136nLQMs5atEc6avBji+/6
liu6JWcOic48BKj3uMNz9u2pAT0Hw4rZBWviJIQ5lRKWBAGf/29PoIMaryPHZYyH
kzP7MHiWIav/3uEC99c6ByVPw2sfESK9TUW7oqi6qqnZbvzwGR6ZNdsIoUWVuymt
Az9nrXUrvti7goLNNBZGGykOc7AnJgQW/2GeZKg//A9CEecX3Mnl7pfclXkqL0lM
5FfPNmm5LSJts4XOqEWeGG9Q5jrBUmhk3tEfW0WkP2L3MTSoIjD3biivKzWo3r4D
VBgBjISzwy3FOgksKOwJwQLrIoBisuLgwuFiiNkdwSkMDNdjBJFLwi2np26bcS+p
ZT7pYJj+q+hrr7ZjxsA/jyuB0M75Paxc8ck7GkKIu0+nC/K13dWR1hzILVMq0jz7
b8iPtZxeAyW2RTp9hTezA5PqhQL+JLnUamLtMI8F+pxt/iegnsGp7dtIiHs1k+Kn
8f3R9ps+59SlvtV4uIEtJeXiHPZfQfShWf94jFXay2IqFBx1OWUHI2X40QQazPFS
K5Wfz+RC3573EhvQE6gBQhbtwKHsZlmO3UFeD+KhADqvRlZp2PtPHyxN4C/oIDDU
GO12/hbG7k0kXQ2BD30q49LhP2/Q0ZEjq62tIHso7fGmoIb4++oX3vQpyXQkmRak
D1yDldApZ20aUVCnM4LOHVXAtd1L7wunWqLFTTipHTtY7SbaIEG2YIOfYmLHmPex
AmlKGigobl0ZAeLKknPWFl/hNiGdOLZ7lG6Po5lbEGFajINwONYXBRZJYOY2BfMU
QgOo8QojDmhpROa9LtfLR13+QW/16jy6kbfhwmDQTxLmZCYu142XFTZeeADRhE5S
u8p748Wo+Pn8h5VYP6yvd9eiurhC0Sg3PzG0NDgHdEqDEQrVKN4YzECGwP04nDUe
AiAEnGQTkiqmhWVpmAqcg3XUgxLnS0Tn/TaZ8eBaEAKtSvNGkV1LsPXlNjpqk2m7
tnPAwzu7+dxifd9c6jxtlw5fX6oZD1wQm7v+wWmIzVeGOJKYrlsS6OE9298ZJFlK
dn/lKLOM7ni3PxaV7Bk+LMlwfpUh1JV6vAphd+uRag7BadDuMKqCS99K79XCEqVk
GVI+mvTRC1AEw+SjmDU0LN81kzDuptByW+hvEbkJDENJamoU3b/FFKkjUUyInfef
WH/n5BgE5l/sDSM/qmqBDtv08tbhMZ4gO2j4cgmOuxEAyzYSxNmZdCsVn3JbYJ8O
3/TjBJDoSGEpqQyAfeLQXoLSgEqJlveWZacicmPRdeuwL3HCGXGnr3LOWkLOJrww
JybE1h5fH8B1VIyXCeG84ctxNLzteniTQW+KwP4Z8dZMvsWQqL+QqI1V6mnBMkkJ
agKi5S9nnZrU6Ll06vQM6Tu5C+DnT50WVOG+8ag3UdOS/LveAuycE/3pUbzh4OC4
BFc2kT/UEyAHqH8XMY7Aij9EnwEl0uUXQ10UrTJmx9lJghyrlNeTUSbSepaeitNB
Uai7Fv4LSsdWSFSJVz/Ww0g/ZfhGvv/UagywfHHGTZBGxpJ0/bXJwCFsa4WydIDY
ombRxVDAIWpJWE59vwYtnqdvCC2gjlxIAtrqSkjUtfJAQELnor3eiTZI6uwCZVu5
6q3t9WVuwNhvSJGpcaNZh8OI3Hq34P6S4aW0dFHawjtK3yEpJi1TAx2NxeompFfz
qCqVOZUl5yojFAFMcfvffg3ujkf3gs0ErQebYxU+YGvpa8UiDMBl2l8NU+JhLL/8
GDwSbZJ2lRccZrzoy62Ah//0RJglpYHLCkrEc+El+DCnWUcu7VGh9cnwS2qKASUO
1mkaFF0o7VNxb/YlsdsktthGj+sgL2nummXt1Ehyg5Uhvozji0GV3AX6+pTy9Y4j
w/C9oD4x/rIJOsEFxzZ7NiPq3hPAiAHGTkhbqPleR7bGJd//XkQ7Gh7xwOF8TC1y
8OlaqNDWPcJkin/LnyYLj6ksYMsBicQemQsXdOb3hxgIuCSSf3506qHa2oft36Oo
DW9uNLD6BOC6K5zWnWsaKNFhJzzNzTkluVtLutlGPx0YqzRHYI3wjCPH1qaUiJp3
9KHWd8+vMrM66erAqcOL07i21BdVzWS/QP8rhLcSQlF56+gkjKAnP88IbskNSKxo
pKpCyKj8GNvVPKrJ2dJQurjKNhdhiEPaKlhtN6rbwIvu+5IOcMFILhd2KHlbk++N
IMVbTdfUsojRwrXdI0leC3UhMBacFxwv+Hh5J8p1XywK9gnmwlyjfNp4WUy2vPub
rZUdfkwfIEagwTT5Hm4dD7IWxKNgrZ6lJjyY4hDWnacwj4GvD+MMLZawy/3qYDaQ
XIAJx4hq42MqOftWkQNIF+J2aVDdaxkPZOkhP3SQMpaSDokouS1/W4gXzOUXUE8l
ZDoeInXPqTecgeh2vWUk13U0K1ZUTIYysnVtpcy0c4ZJgMQbpdgG7XtiCUpRBcTn
FY7BehvkCEPT/gX1kfLloHji5ilUlX3FjENzg8HKYPnABVYCZ8aA71VXqs/e2oK5
kDT5TeEikIzOX79f58REVwUzEmMm32bMDTXYpCtvii7JB9uQ7HoN2FOFzio77lej
//xKxSsMpe5rtrBp6gY8UayI5M57vG+qBb1z0qJbp1XO79z33153/P74PPi37TOR
+ne8IokBOe7lLgSTMqB8cb0nhhoY5leUHuasQtEwO1GbrKZyDPlPaavmWvHRu8yo
X9OhDyeTvZPZmdYBV7B7K021SxrZ96tt+FvHSaWUxQwbJls0dKMzg4wPCJibNGrA
hjYc/4XqIkJPZu03wvwl1BtPqW4fAZmuVTN150UIaP7GA5tTAoo/WutH+nmst2kC
rzB25lT5tdBIcR7eWTdJSA8xr2Lu//hYhLugJ4LL8JuDgkRFaOjbYMKP96Btfl6M
F3oNdq7TArEskzxCeDUNlCo+5j7XWKt/1AmpooCV2zX/TvIAfqCDD349paecE+jy
N2GZk/W/7AzXpG6txC7CcKGbu+kf/K7e4fLdm28BRxGqNo6cMVWo+mzSBDMpqKpy
u0InnKAFeX2qlr92WP9DTXJB/X7jtc+GCTKtVglnX99VtVswgO772MKw8VGsMJhJ
keXxzmVINS8rphJbPpFK3h482AjMu1N8yZwjFztpclHSKkHwnrn1QjCV23zFN7xE
ZAkeGiZ25mNXySpJbAox8bV3EIKehSAXYuyUMQFL+WXXufC1yciLbEYxq1SKwhog
+y+sfCUjXJy+ukBsb0te8Z5G/J4ooOSbtZIIg40p6rxBVZqVYh1MXQtPR0hbODVT
miqKGQ8uTuVJcrYXNY6qVvzu/oASqELq3ZSeiTSJj0vFT35tp4h41W7vIh13PnRA
S+lhs6cwJkteq7quyF9VIv7XxKHWs8ZWpPeNdyEJA9Ce5OF60mOrc+6MECVQrStr
8kqXosNgiWf89UOQHBBUTWGFKzIF7sKsxm6ZmeijhuTZW9kU3h+D56Apj11kFFj+
nmonwezpozb13834r6ufZa3J3hpt2jCz7dLA4Oza+TfuPF4ouAscd5ID3l8OrC5p
fv5gf7Lyygx8ZVyeBJJZGluICCXhutt5Q+RED3WK+5DQWWNuPtXnXPjHd4DwzZ5P
XP+/r7fh1j2jWK1hpQxmEmNKMkSohF4dFi82pjjS3yeYcqnXpohIJrICH6lxfasG
65nJ0PtNGR4OkSA72iEz94fxXa7lxnCBu5AhvSfgKRUYvl+aTGGGKM8SAuOkmulU
WOZqrWGdCN6cP5e005fzoRnLMPtAl4q5G5y09CR5V+h+D//YN5/Xm7HqXlUQKc5g
vAWoK/U+Gtl+3h8sokdTjH+NhDsccDOEPPnzeaMNKL2LR7cMxl1mCOxz0Y4lkxPq
zeTWorFOUafnB5U6DdYBVuJN3wK2L3APG2hIb82UP8zmE/FPcLauX8hStLLUHSxZ
QhZx4I/2fkYW15R/G22XTDSWqyYobar4qpj95+MNdgxpINxmtsYuLhCvy6DIjjOo
WvSaXbju+ipH50OQpsw7JmVtOK28/5BtpAoEFLR9lmCDRgOmbuJ5ETcOkb5SBK8L
Ub/8WLK5348YZznXdTpo3hyB+u+lBWSE58Ujuk/OpEldg1M8VFmksJYU16xdbFjr
DqlNROhr1OYFfq0z+Xt9z3X47hj8GsB60+1LuusOeLpBL20lMGzHqIzckSyXgXJr
T7YePjeZD/0RSDU8Ov9gZiW8b7Zv7UNlscMEZPaTbjmpl4OIRzanQsQq8ohCeJ+/
JC8lWBJQfaNVhyL3ULB99BZJAY/+Zhh9Hz2TsOFw/bdJYDQBhzXv54lZbONQ6ODJ
SOvXVy3jAuVcIfsdwFYlRVy+apHSLUEHopP5JJw5zGHaaccMtezQl3xgIPpHHoZh
CRVr64w1skOfjPHTIloE1LZBqtj0OE7QZs03gDwKRDzcveHiGLgTwy2/Vz5TXzp8
7jNmajGA3sydNd9U3qOCeu8UZGVdN2BHRokALo1hv5L7egtoAZFkzR38xF4gSweh
czaj7tmYVyyxOBWjZVfv+VlZ0rEc3JVrGa1xODNzZyHEX7JARkvF+PuTepS+xy3N
/PmgSO862snuikuP2iX/OBocIkhuoCBbSytzu1KpVf65aJ1CweNYqzhzUleQAM59
6u7rjn/5MKhyNz1ULeTY9iFQh5sHcWq1uQoeN8SIUZqbHophzKMGx0kiwXiZEL/n
Bvihbg95Ut00aDlabYzL8VoueL/s0ok5JIwXngPNZNAlbuggbW53TOUvIT+2wGZK
dV2UU6usR+AbI5ezi7snp2quLl4iYa/Wr9lgTOftejhMHEjqY9VrnedaC4EIEJnj
Y+uucjkel4TGq4P9/fHJe8ANR42Y3vzUvgsOfUjwguzJCcmWYp+Xkckx/9V+8aVm
3T+O1XIzwxDJrhMU2itMYkcga5CVAN8e2sdVeSPATdtTuIvnBz91yI2E59tw4b9C
ohLV6KumaKFUG8rnOg3q0dP3Xohj+FOVmEV04YjH/bqDW6MmWeJml+NIa796uA+7
xswOKC/VizusmcWv3Og4sx4uTcfzTRDhHbjvCAeBF+jZ7IeecHXsTxleiU5wG+/D
YcJXfqZd8sQN2zat6UiwEV1dzI5D6oLkkSv5Lu/KRBWVIa63tZ6wjiBFAe33BEqP
y1df3nbAY3f8vEUzk+s48knyJKD774dJVdITfDC5pm6Yem266hao7vL02pic2DU+
YDOcie+mXpTQBc2gx4boT/IlSdG6TrV0v1n1dwl+4BOHQLqMQTMc2pGx42U6wbsW
NO6djtBEvGQ68bI5EmW/vHNBVAR4utysZmg8An4VRjFiA0qdB91umOvq6SpDfkkJ
57LJw/WTygo8HIHlIuYJp6jNyjTqlPCjQgsaLr2s/+dM/4YUQYJXSf6O1Y2mkBXN
5ieD/9rKm8F3vwxgxePX9vAOzOMRx/jXAuA5HIJjOZ2HKmr8Kp7L69yytTYps2Wl
vIZ1KImex1OixVr7Ni6Fgal3vj8RI6RXmYDaohqjdp4EDpDcxK8m47LgikHArTwZ
wDezQULHH5j5yz0ppm/lkldU0aQWir3RcG6NR7RWfgeLNm53FenQGankk+VuG9WA
YM1utuH0PM6KOqX3p4tdOYpuLcRBtKvm6KhWADf/SJ0Q4MHwqCzntQrEKY5Zmfq+
IgBkT4/MOC7Y3q0Dt42+SD3KWRkYjAK7mqEGVJQQewJjx6dvilUO0aU5vXdk3xIs
LRjsHWbX62lRUGZUk/WldNKUBKTisuoBN2qeL8zuXZr5haItmiYWWguC0IacKizM
xrZIBsEPJKpQT6VMLfm6uElbzoyPNKlT1SNeAyhv+GywcUuxRTJxOQBmzC2anmsu
7HoCtAeRlfcoovej3SbS6n9nblkH3eRG9RZhxzMY57TEa+9k0TjomMDV1F9U7o31
ReWAKHvr9ABLtcyevRD84ZghwLirgmqD2OkxTGJ6j7NG9vFoZkHUVylOdRgJQJZU
RN2fHIq/nLFtuYyy1iZITl81kmDlCj1Jzra6KxtaN3STSCVLw/5Ur9T1hFt/VXP2
FuTAvNujpK0HuuxMqqr2QeJ09D0f5JS7eQp/yq8Fgwgrf06PrWrJMT4wVexWJYsK
ugeQWEPVqv66sChIBjX7DgGqhHgBAmRINo8e1Lwct8QRMfi0XIwtYRKxx9ivC8ga
quw+YgEIRyk2VJ7A8aoO5klqtXyaUECQuCfMysifr+MOytST3QYLDgh6RW0PiYGj
fu27DpdxubHdyNMQQaczDApt626CiHPKGLtFOO3Sh215leDN7hHQbjyUyLoTuoub
RYaDON3l9pJNjP9zLneqT2kHM0oBliZ6/95wak5rS7KnF+YEyql7GrD+SnFo9Xex
HHBC0aXENEaHd+5jvdbS+rsPm1d7pwUtFma6qC8XqGHHFQa3mCBKKpdc+hlXL0iV
Ob8LazocC+zEY3nG7X3K5nZRX/twOfSTLkE0wbAhgfoEoBJAZT2KvDIukEjVJUEM
Ijn9/qPP/5sXggHJJ9jAx5/YjB5F8tDqv3RC5hkOLN5O8oGfnCfQurHJ22CmqyGm
8Hef4xdKq1jBAr1tmOUfL5KFjFUimy+WCp+Hn71c9YBNZ/HP4i59ICW/zZvVWyDg
zF2lfr1PbuBvmvhTS0Vvyuf6xTUGs3leVFJKF82VvFw5oyhuueV+FGumLX40/z8K
lvZtl8xGwPTNw5c8p2udyPi5IX4q2lLv2Nnfy1In0VN1UwN9O6U/ApC6EaqlHc6+
6OTstpbcVzmpl2+4yaPHb7hnYMd8lFi0ZsFn8boFa3kGcGMS4u6SGD0iepP95yVM
25AUoaF1+A+bDixn7t2hJ7j7MMhlhFfJyJOvdmsmRI5riuRgYBEFV8Wstufl+ISa
2JUwguP3RIqHe9uSx/DATFfOmpjipjzFP2Y9CbEry8xwCi06n8tbPVPYaXCTtEmB
MkC0hOC80RpeaSA76CGVq7ooVTSDtmaElP9AIU5ZXNPtqQOZbLfvdA74RjQA6k/F
idCiRIx8sZrhO8mWGW7IzuS2XeGYTNO7jrCsJz6MMqZXIgmKjDRvuAWRm1U0CNjG
hY2S8/oBesnoIvwJdcXZKUz9GPjcURo3d1SrTgHhSFVgLIcpZiL7lZsYuNHzOitZ
nzTrGDNVOY646oZK2wHz3iOlgxkL1jSzly4kg1SkDt4dm7q1SVgz/LMtmjQhtq7n
h7lZy8CZPr1Ud9YmHpjNIg/02Nbdb4cfRHCxW5dpnx938bmP2bSL5DX6MwHlnmpd
1nupK6YXnj1+9zPWSKya+yEWriJl/2DmiTpWHwgfGUfYss3E0k9Ehfoy+utCY+sF
z5kol4OzqFvd+oVV5+Vvl121NhfzFKFzc3xSz67RaOpH1UN2eruSnVvJDYer6G65
/3LrPPGCwhoGpCAZud6tUxijMbU7KeKT6PmXL/zrme7YzBSOo+2BHR1d/t6rEBmz
xPe25itDUq4tPD8dcJKjGcnFyecmuAUBZo8f8uxXo0qiGxU6uiHGUhiYAwkucOvG
d74X1nJaobt7xQdgWv5RvKYzZ+kVHytNXnI/iZRqWNPOwMpFMdRq7SKhpEan56gv
2cmKBvFCoezPrXFjEIySZqScgczY6NLPC3LyImtW9qzmM1jwps7oqzFg9Sc5XGuT
KGaAGHEVoT47oScDRvCH1L4Fd40iTBqhsv1/xOlPOMh2uXMuLUADDQQFK8G9n71q
3wp4jd4qZbO9KctJjhgNsa9Ohs8TGEgyKYoAh+JWienyyieRvs5MbuOs+yEQw9nk
LRC8ZoD2f+OEox3JC4520UD9j8Hc/2b9GWyfRrKGvrC9CbIEEpXrUxcm+L4Oq47C
LUFpm/w56iOKrXCQKaohY2lcEFKqT30cENis40V4rSg7um09ClyctQ15K58N8dmt
JiQu36h1M2W1Dfb4nAjSl9WVs8VJwSl5WN2j26FvTHIXjkP5hP9/r2hJI2XQwTQp
vgvytwWv4mE5VNMvjVdxG4rS/4tgw3KAEx65GBPYelX+HBDxuLOnqwPsuwn0tcEz
RxlUukTEySWKrsv0cLhsUov802/CRmdUho7tNE64STqkiirh1z+jA/rBCbLwOS5T
CAFoo/yS3oJ0a01eMOqOP9CJGRxElSvy1Ul9wXzG8yu7p2svgpixB/B+l0YrVdfF
sH3VipUaxC/tuKkVNwO2UaHvciFjT0l2ePYI41CD/k9FYhUYMiJ3k1RSR2OaXgoO
9JrB9gTJnwvpPL7Jw2CNQk+nXFfsvfAWlw31cZRpgZD+c8ceXZAIy+3BVgOzmJMX
hPVGC+rnKzzKsMs9ng3azol50lOfuGfpDrDzX5POT5jDQPwrYiDH4p8fp/rAuqi+
J3iFjK8SxLwnK7QaIfXnCS8u+0CIyoeKbWB/cFqT2N8/eQqfdclU7+/T3tsRiniu
rD6rMXGE4zYWWYDm/miiryg6l6mc/gYmjo21yP2Yaz8+JpyN9XbBnS02GzWcmEJ0
P6iw7FzrEY8f/1ye0nvqA23ihtiwHa/jrY6kCddvmawD60dC4wUTzUd3iQvmbDcD
MnfrKNQtaWwXb4XQQmquP+ha1TAAex0H2+ghPdPUHmcoAeB5aFrhDjx3JZxiE3R5
/Ex5wI8JcdF+KrMdowQTZJ29pjSCLQPSCv1iEhr1nyIfqiuZzG1RTSgmdy15jR6Z
X4cqVLCkfGETTwsJL+eAgSdarluo0YsaZdWH7gOCsWLKqzH4VoN9IWg0rQ4ZVxoT
GJJk2ZHYPtSF670Dbc+eDlmrQqa6iAjkEb2uyZ3oLzG7POdMyWgUrnQxAVe10QqG
affrxPokD5DkWYUpcDvpNHtbzedMXHB9EZkQ1hWuBYXvFWGUlV0hh7Bphno3BDcK
Tw9q6kJe7rwJvHQdImKBflA06+Fk9246N2L09HONicYLIWG2ASt/ON7xYxlRYke6
Mgse1D4q6TX8OKhUEAlvfNbf8a7ceAlYemKTUHVMO6JDk2ynT5MpZbfH71VOHlwh
Lzgvg0IoBLq+NFOEYFTPaRKjCozsgl2cv5D/YUpimxdlTpc3OJEFKPIBclKtO/Vy
RTcrPUYv1lt1vqSgufqRBAJu5U7ztfU1OrZZFVpBiYfRnSBnJ6c1K5SPu0vBAj7U
/KQo3l7H0ElRxLaYa8LkvJoyhBaAW7FuHZW7fKsPcMaI5BY4YvEMP1DTLBgQ3P+B
PE67YlXMxsfGFNzsNsowZQHtsJTC1el37N1lrZ15qkUZEpU7znhW750FrZA2O/aa
ClTXmP8rTuvQ+6ZJtf/G8xwwsk8ah8kxtkfDI0rkQ9SZNImyko569Tcr33pzJvYF
Umm+1idd1fsXJIbj2U5H9JIlmE23sJjRUeywLiKCruylPslYciuji8aex84MWn/D
ay8+E7xoP8nMoL6HKOIj0WY6u7FSQmvFtPgGE8GshGbBGxaLFUoYs3sjkAtz0hYR
6is73Ty7aZfYBjKe9bwuBPOnUZRrQ8ywivKCP1Z17D6CzDqAGi267Yda77aoQD7y
umt6kO6LtpdVnWU/hL1Q0CZkNsH0c0c5t7NTFAUwSaMMrqxx/CY9wiOVty1sOKBk
KP7Rc2zXzKIrxDmhRkrNOGHssngAdfdVfGxDl8Bw8pxOHItvrZr6v3kd017DfQgo
B29ZAhw2hKoF5HuJyyZ/ftyWWxUgZkzLuva2wB8GiXuUotBpjuIibCU8q49RDjoa
gDNI87KsyFyaQz3nhm1oUEc8A4Wm5VQk4j4gkoYGWcn7bkso5TyVEyPR/bB0uoz1
KXqqEfubV+TSFNLZqAd5YrTVsy/bUHVuFQEqEaKCWsBWCTg5gFKM2IK1pvlYzNgz
dejvKkyoW2KHr40h9jAMPYzccE6HzuLmPJMNGzmK9KM3hU0+QOIxUH+qn3wCCO8u
rJTqLAw4ODNU4ZE0L2gJ14Cam2I6Fk6A5HGW0fBmp4gLIr0paQ82hIuMb8jcj75n
VRYZ0BKec9uBbD/yAa6RVh50idiRelB/Oiq1YEzUb5IsK3m/5Fse4UJkkIPPPQgs
y/ey4ZFB3gSUh+rBKFzFjNSp3vieLQMhxbBDgYVKHfRGex7llZzt8g7l3fAnbcDs
EzFqhX0NivDv4guzS0p6SCnDfP1J/3k0Iz6eSnZHUgIJV5e1aJh5TeG3duLcsZJ9
YRvI316qUtT6IlGFLAva/oOPUvZPKNXSqqnnGh36FTPOYJ+DZ/WLMjh+k4FkNv4d
k9VBBYFfXHALOUw+lmRvyGRWp1BkRGT04kwsThdbUvd8qUWGyO0qP8LkKg70K7e9
u/fFQigHFwQPygQr4BqCpYAtdMw3D5CCa5pdeLmrgKxUZ3DTMdM1R5dZN8V8GPE5
cTFTYtfuDXFjzUAmVRJycqPYWk3rPaE1oSUJbN8bNWCmD31cY9MkDO3Kqc+ku0lR
0rGzdKHPhv639Dji5ai0/HoOmIgGtssmqWl71eCtrzstQLgakj7U/zVrKRRs/hvq
0gkrhoRKGNGDtVlf6bGU/DIb7bqJSD8ttjT3ci3tN4Vxqt6r7Mg5tv5/IJIWpIYc
LDgXZi12W9byR2eqVyP9wk5LkuddUSsLXo4/zOUyb5LDqnlQl5y9DR0/4FfYmQi5
cajYmY2Hs35c5Jn76Ie9GnKQhtYq4GS/mKxNN+gWvufY2TcZ4ct6DyR+evaNnAQP
MVumv3RuITWHlleTeFAukomhED24U03Ehy9cUwBdJ3+u2ivyMBUWjt1za40OalBq
PexwumCUU/Q60dP25vdBuXmAcUHEJKe5Y0hdxg/d2zrA5Bv+6ec1wQDyFWV3q8y8
5iEBxx6e/rB+uIpheG2WL79g8Meal1xyLQtfQoLz9YlfWK9yL+Rr6vcsdcuuviG1
yyOlNadXRR4WKWr6CkVVJu2RMAM/OpiIVvhH14fCeqA2JmX4ASsYuFQZHjYV6xCq
MdWvhgjIdePGNO200vSppmhcfhkobc0MP19u5ssSvoWz+T0iI9/Iy01Y69npcEn7
cLoURvHEXn4mEyF7mSKJdI2ddyaNxvzkH+iRmpxd8J1BkGmWtKLi2OdeXcUW5R2k
4Oz/0GswK/hbnjQESs4U+by6GpZ/ER36EXym6aJwgJfivUbqud2Uu/DVgDgY9tBb
UvzfO+Y/GGP1q/CXTeyj7SgHMF8XUkJR3n7O1z2eNmjVvzGJVpiD0sbWoHQbLsma
hFaCsLpnbjEvVmRd1o1zMvIUBYBzACdC+Mqg+C6H46odp1wPPRKCmP7dpNoZ0Ygu
YBaBkxnFCgslJjP/lOQANKmKns2Hb/+VMaKt6JF26OtZEBd/pxkydfCp3A7fDlIS
c6Wz1BUk0gti0f3YxbVrKWuh39+K6hPn45DeH7+Y7L2StoJt9Lj176CRK1N7/sDa
FRW/NPOPtEh0QQF+Ff+xHXLvfpypgyv8IluYlfkMp0hh+trdG3g6fcJVwX0O+q62
T/XZ6Iau8I+kiuyq+jhN0uQp8zgZHBFchMKZxSY99pDQB3KizDF5x50W2MTSX+5w
QMSBluHG9ZRGLkiQ2suJpCUkYkxrwljh5zc8iVaKenxMKzrRY7IJ9v+V5hjIEGkY
Oahgh9rJEtrOYa0dmVtfWAjNsPlVvUBbOemqXeWUqm8mu+UN4MBLdtKAV/y6QcOB
U33EhjfuyU7VN0ASsyAkzG9DG9tZDKzpR85YTheSd7szVpUEP8zouGOJNpalmRVr
Fvf0xXzsO25NAyf3TUvbfU8664esqtBPy3DDr8fmDAV9cGMJ5ArMeSE67ZwC+mQb
qwHsRpVQh22/z2mioLMpKYVAks3Bcu+/UJ7xMJ4WJ/hC1pm3tNxmj8g0eATt/G+I
Kg/BBddfAY6ysoq57sMqo9rR2lJtfyk0On6/ECV+Z5j5C1PkGG+BYrZxCNWBCUTz
QADcoN/ncO3oj2l8XRfjHvrzKZ7UmgePd0ta4zjpaEPuJVPXnmRg/YKQO3nB9Tnl
h8ysanAPH+k9qc2sGzhkbJuw+2BwKepYBKR7VmDHhpbuYUwo0efKcRjFjO86IJKY
Uy2es/LMI+k5DFJrd+lT1b5kgwUH+gIGCjcYHovbFlCxGRBBvaStSZsDA9k+hUdp
fJkcyCI5Mt46GhVvI/yaI4Spoun3aCENm0zSXt1QtfofY//2lL4Xz+Zgw/HOqhnH
WmLkDgYMYg1+cpOd8tN2KNvT8f3NKKjN/oBVsc7QBIap0JG2c/vVn/wGOaJFAgc9
xVZhtTHfGcYwGjtL7h4MIOGG2TZ68xTE9wSVZsS2UG1Hgd6nly9R1PuUO/DkW8z7
asnegq9qGhwcCbzZPnXTXSMG6ryoWgpQOvKtOJtycRbjB0MGStAknyYFK/FAlu9y
BoXIPcB93dAusNpxkcGkbHEBf/fc5RSkb1E9lBhh4VR5j3pU351ixIwaa3BzXLQs
BNscRnnBRKssb4kXzelEtbk7xHN1jHUP/hFfjdJ6S3tVJ0D9iWSAEDWlSWkBzylb
eb3H+Ralc32lgm7BrQuxNFygb3wnhNsQr/4lA/PYGNqPHkOCGFGvEOFuAlI2qS8B
ZzFqdYaoKyb7s8Oeic+Map0PIvp1ExJxJtJyhCGs0dXBW7KzRsAEl+s4C5+cikpO
9eSHTLZkHdLQlj9FWlX5rAKxMq9DCPhshm6mQMzoZidn+OVa9qiZDIU8+FgKF9dW
ebu0HFJ9vLeNOKMI6WaRh9OhralvLKMfduL1j7oJbIQM3VAzWcBZvCyXuqOL/pW2
vZ9aosYl0mOVWlodY5e79qnJJD06jAtKmz+/j5N8TANRG/I5V+DIv/yJEzTAUP24
mFzx/FrSSGhB9czRQEVo3ctHtmBdaz1O3/38OybGLAG9p2cU0ZxPP53Ywbu3mG7D
h+9DrzrYuNHVkFBGdKqQUygch4L8l1pAHNxUgQzs7SIEpkCeQTNRQFiVVGtPJs0c
hU/SRokcR2tY+SxfBsSvemt8oh8WpHz+icPRApXkAtpo93UK1iUl6ITFBwgQmAHY
rdYa99IfjAQlOZ4xlMVBrWKyKbcM40nKnT9UbJ3Bjxw+PqxnLrsHqlNI4dVLreSZ
6ZX6TQdmRA34enSw9cqjYCgeTBr+VUR2BT2Bbj1spnTceFKNT7Zw8A1FGyA5W8pj
/U+L3UGWhqMa2n295CzW+sWodRgVL1DMOXhHQrvLHkt30GTqrPi70DKARhoX5p36
tDi96anGBcx5lSP4vfhlzna0EqG9kxpKvNIsQF/joZhYiw4ESnZfVQHVbNZSX+XZ
9Clcd7QXViMvbGIy73t62ZxeJsgVeFdtlybIbGHrPJ3yW5+/rPQjeTiBysOtNrwY
sOshbPrn7Q7+3lXF3F25ivyiK9dtbDmfuH+DMZonFtbyYOcUe5pbSoG2mlUJsm7g
pQeUMXtr8cdWZkWfwSl4NhIea28m5+1Oj7D4pBU2PTit6D17IYzrmX67r9kFZB+n
I6NF3sf7wqqsbzZfQuM/P+0RdETkXp1R1aKvZWSXTR2yR4HjiGfAIP05AzThrXQF
u+7gx0o0SSs9j7pb376Kew46f6/fyZtD9ugXVLeQYQCMsVZCfWPwmto9LoyMYxkX
VQ1BSJ4ZlxsLnyk7aAKVuwUOB/5rqO0vBJDDGTFuIeYAAgTZil6Wzt3AnZrbFbv+
4M03HFTHgM8vPhfOvimOc49xTkFn0wF65vI6fqfo85NtOSyHlKcSe4uiBObxVnXS
xjwJ54qFCnCIasmSI+zg+4LzzZDiYHyxSyU4N9WGDa/yMVL3u76i4nDRgZZNExxf
dBff8+K/2wOb/E1gu92M4m+7z3ybTDLPGlvLsmCcrysVPabwbNmJb0pPz7iJfPmM
PCzq92FRBfRq/6RlFSF1XoF2ZTAmOC+nTBFiJFBlYnhq8bRBLfUG7hUiUBEfnBjy
agwowBhCqAC7XY2riaNOrOU20klb9oBpy/f35AKP06eIFi6t3ZxdSmWEmGvQ7xs0
E1ZAbtypD6MK7Ih64Hjf3sy+mF1YE3bqUXu7rODNxLrMQnehOkvxjiIrvpaA03lm
MKAAktWY4jUE5QEBi4BwEfm09X3DKyvB033hzPmuGd+HXz5V0ilWnFAzrp9V6NSR
vMRwHcAh9trLwcVgdeu49r9KUXw0S1qiBKbu3umgbF3TNnlHumLoOPsqXVW4nTNP
TuoRqx3eBDcKerr4D9RYS2nYR7TTyosz7hMGNWLB0iPUkG7238iT6KKG1LhWHp/R
R6ABm8+Bvi0xAdXTCfRSK3UiptAClO9f8haSDZ5elhnnIz99Yd2ZjhAIPOHmNPvC
r7zzhta0hrEg2V/TTb76nyG2cgbIpQCwWOfpwPcv04CFR20dQwvUSUIvFgOPeyee
KgwBeIwCMdpnexBURrtrdC1kjYOqBj/JfSOREJrgRnYo8tsOQItXCmArboI38o45
LlaGdP7ZbMpndkSLz5JsnkxhMDqpGwwzE90dDTdclO8dLvUaUE82Xgtd4/KoMzVT
uTcaWsRsNcmrxht/53roBA0yVnRWJsn9MBE0+GODnXRnaXFPQw6Mv33qJAaIVibe
ooQ8Iw0YIFAfb6Y3TaZX+fzZAvTLpJBjgIlWWE8uW7JFy7mTDYTBN4stGAIPs/da
hO6scE102VgjdwYAHXnwNC0AAnK4ohyVb7S9EldxtrD4xCamW6vVk6ZIO0VdfYH4
TIXDbOIAIonQnKycV83UW9A1jdBST6emZGITsKOfktsua/MHCz2z8DOqPO7XGWAI
bLnWvJZc103aCNDMJr/MehuqGmlYbTvKlK7+qBo2FD+Rlaqhycr5oQDribzbr2zk
djsTfZSiIfCRdtZmuGpkismKmriSpN9Wk6Vxg1OOw7L/j3O+TsVSLUGaR4nAQJOP
jB6+zeAJALs4hEcoLwVhhmYrstLvruVt2AArgVD5wM8nGivm1MjM+bqo2/4TABrH
GF3dJ3NqWMJof71dU+XfIcxzrQwR+r5JYLD4k3yFLvUJOOHGE3jqOF4LdcjxGHCb
iaZKX/HxcBi+00BNqZhrTBZcKKIEY/a3Ovwcxbi2uLVhoV3w/Vuc0jGj8pIYHjw9
owKZaIELG5rN6jeHp10+vJHU1vdVIq2mw0OcHRIKW9ieCJBXxXK0aAuWYCx68Uoe
fqJTVFrqLcanWtTQfdY9zRCunQnLp8cDPbPCFIvV9c4Uzbh0h6rja63DtzT+T3o1
u1Si/WynjmCErectMJoPyGtQoCOnq/JzNVI7kVBqllF43MsibJ/wlFaTW5DEDPU+
ft5BrjoBvwTzkclxR3CbnLSHlGrg8ZgUefADQNOY8HhDv8xc4GVPdNrLkd5UimQc
trn91F8mHJ7wSnaMnzpHbFAsjww6Ro9MYkhon+kpezw2pHIS6K3Y4vlQlpxu/N82
yPLjfL4ZuXr132vdVbtisvcpALm1pNBuOZ9zq/nbWkX8JXCy5H5JfKLhq00b0KNp
kfyDShawEE3dL3wmSCpw2JzLhFyYKsd4VAgupA83aTRC/w4oN4JV+xjAA316TWj0
xTtEuf0SyqH9LBDZcS0iAugwU9tvHilc7s1hp11NS+0biQcQTxgDSPmIxFDPjEjt
N+UKUMzCEsSoslP2I0HWcwRlE+HjBQoE8cRP45z47RKQcRDCvE907iis/pw8d4Jh
q5C4T3EEZ8yUWYyYtx+EkNS0VdWHhOagrIm0Gc0y8MDFtH3WN1BWNQZhAfJQyd1G
B88pwAkHK+Mny8t3pwq4gYDxseP+Zwrl90ali+TKYLLD80LeB0rLhJW+brAsAHPA
486dE/MYlzJ5x6EmHAe8eaxCILrAuqtCgmIJm2CqOrKo3HOZNrikjmlZfDsS61kq
WpbYrcCsqqBpBW0vK7Q4xIoeEvlc+IxcVi5iM4HsxHN84mXDIDD3kNiShMOkmeHF
VS0llIwE8U6dEeiqBRn4E1lo6X7kqui8/ztW6EE9P1lDTG/iRNL0zyIcHs3qJuIE
aMavB16ZZm2xwmpE+/yoQbKz2J+KXj72XfTf5YhX05KburoNzI5GvHxnXsbnmskb
N2EVn+XuFDvX9yUA3Khunt1GgsQNdn5mcjkWctlvLqXnsqI5CAno7e0zbxnPY3PR
lfQb2clGw8vphochYIh7j+4p+h0fyrfo7gxZTF353zQ/jX0z0zWb5Aj+75wg+kwS
BF9d4RG3fsJ/T3hqiwlOpoWyfl675ZKlrLqWLTVieTlJWDIXU5QIamrgKjiFwElk
nzC00s//Lri5Vx/gt67X9U2Ft9QVPqd1KZEgCcVZtKzcbCMpYng9zN38KrOt3m59
zS0wjF7n7ZjUb3X/94+Ng43BPkxoREq1tIKoWE+f3/Ug7wdryDhWsRWnNZdIT2pd
CWwt7hQFcyzr0xMixWLlQf46FhLaSdHOLLTjF4gOTzDEB5aJ0AccP/F4BSaTXX0N
5eqqaTYTiBHh1VkOA1AZibaUkp+1ondPnSeFFQA2p32eKyUVthPun7zWMa7k2Bjw
+ubPK8DZHs4B37dE22DG2TCrGyqcZu6qrzYi7XE+BOecxWeauAJCHSJ6KQAc9x5S
uvg9+q/gCrxtMaVIA79bBDAqH/awz1IfoybBxGLe0Sjeo/cBmmiR43CbKAjX7VF3
Lj3S857BXDs+yTssHcg7Z+2uQ5ReTzSOy7h6BiqwUo4I/HJkuOpy/fyKJBNW12ZW
wWcTaWqJONFJdRykpfHQW+VHt3kwVfoizYDdnFYm0JTYAeJ2JM9SLbY4u2ujftnS
TDsk7dGt+Y8vBfabth8Xb1wO525h+FCbzYuL6NO5qXT1B71SjiwnajgZxioZRo80
tOVJTwZl+W8nqyn4nmD6MNqopZjvlrWR4GfBnL4F1LD3cu3KACaM6Ivdl3hER9H8
41yx9qDqLadA4l5lfiBwNSVAXG6bxaRUsCMBfE8S51sA5shqFMY65cKWCk1sNq/j
Gl8u8WMt656Ax9EEVXEPqudV8YRI2NBDOkXv6sZ3kd4QQLwhmHfnmfMXEXRu1+af
kYjU71XXalJBbvunN/01GF2ph8vWKleUWpgEnZKajBaxV5SwkdSSWtCR3wC1+5OJ
PeLYr54ex3V8gXI/DuPwYQIzScdk/uMS4Yl/Ml4edR946eIpnWwjCo7olbqBpnBN
8xXewy1F0ROeP/v1Cdxcg1UEW75JuJbejy631pD24sHUBeta937/xo4efybYoxK6
LB/PHWzSZOky1+LTWO0kqhZA+rhPw9/Gkzev5Gv/4DJiVPxjBKPEPkiPcT/nonai
7n4LNgB/aq/wZco87edDJKDb0QbuXy0ibeXQqLyTyv52QtJyZK0IOTL4SLNzN0Nm
mFvH4o3SjP/xHB2Ez8lEktiYqohN7vbNvkOil/iqHeKzlCC/KK1/yj9CBPLpyO2P
H6ueHJPWN1pkTiWcKCj7oYxrHKU2Hsq55gq7389IYC0jDuZ/w/vEK4vWFz16aXRF
Eh43v9Mi1zOrjCW2dgrzUVMhwrjMEm0BFJu5/AlM8gPpGb1Mt0BS90FT3o/LJ3Mu
RhqU6tGKqXTwwqtWY5naiierrBwG20JxNVrpeg+ImAyh7nVmunFX8omLs8W7iTiy
e5JQ2HJSRTHKUw9wHiVYO0uUDBKcwpTUjuTnOIeT1uTX/uXqydXuyoG2sDYedmSG
J8JbdOcUIvNStgijHgppvar5q1mHaaYAKwrnHPiWdQl1OiWVaYCAnxjCHAovAaNS
BOH61iybUc6Ug7rnvrEVOXEz2CuDq19befH8xr8q8P+eAWNlsKanK+goQ9oGMZ6G
DdxaqSonLfZOUWDAOQBA+mEa37aE4gAGNoTJPl1w0iue1uG9kxsRV/i0mlH4S6n1
bneWwP4Y88p6zs4UOKc1V29y0xNTuGQPc4HI1EHNWeM++HCH7ehwDkj7wTE8iuIL
TS/cl0pmzrF4W+KhyifdkM8gcS/H9JJL0Yo1/wH4ejnaM3LVVS1wrtBf5hueLz21
ODVE4xO9ERpH/hCvt4+jtDFf2YzyNVSXLmKcwOr2Pad/h9roZXqfL2Wq1kTzu6M6
Awv211RzJCPN6ocsR+tJfR4OaaeOJIFD4VtvIKZVSR0uYxcGT1asQtaZ7caewU7y
BC6odrAbIoCZeeIH3xvswu1/nzOMV7vCDB2ES5HZFaEQ+V1kqIs3Tk9Yh2pEcE5z
9uVytvY727Gnp4JKWPLH4vHF3g7UKv0lLi1NumB0w7rrsJxzWBhty9cwdLClTRNS
RNeaDJQOkxcurah0+rfomcLtzd7S6LCGy6ElTDU+Te2Bcu35hm+wD1oX4rZiEniO
5nX0DqHxtYEGLqWFzGEmpBimno/wKExs4zCArdIjw0MfB8cE3JQdk0kL8X8F6+8a
auudCHCBDo+Z1KeSI/vfoGl0YODIA3p8SlmMwjX8q5rNMKTqp1vSb4bjw6nfIONP
6/lPTDSpxn9nDTfhiOjzS2rWGqeFCVMruHSHSg7vrgqpYowhDFCfjbzbSRzcX6iv
GUCof0WdWgkLe3T/f9nCusphr3vDs6WPRrwqpmLCWWN1QulvP2S3Df0uuPBG0sC/
vyLp3Izv3PViXWwXpTdgPyinyBuw/9dYq2lASA3LVIre7rixJHfh4f8yNkuGBaEv
Ok+dWhkD6FCMIbSZJuW81ciMv/zGXzNcpL9n/dD0q8vUxWEvP+WKCjY7Rr0gawUR
vxaSZM7ar/5WKQFNfcQc2W+sDwAwMrBH0zpy9SZ1xGygiTZDwySPM5iz9+tOIP/x
coy7dziP9PY86IFR79Zna61L6Xpa/kEiPJ5Uf60R+9IrvV7yUA4I/v5O3gbD7YGI
EHpG4+wJ8UeJKIAfvFXxy/wDL32eFg+1Enq6V/HcE4IVFFmPxo0W9YjuYztz+gRt
NjhVhmllTeQZYOhie+nk7mvUfWzmfBPLf/dd4AUH9DQMbaUIw7JCcTnDwjH21S7l
laiIY6uKujx9huBRZxcno6oXbGp0+44S+5ISj+YGSZC7G8WI3c+QVvxoVr2tLxfD
iKS36xvP2hD4CrW9FQNJM8mQH1Ebt+Gg5Yr27AlDhqUg7LW+b6Wya+6jihjKt7bq
baM4GjFTlaNordyzAZkS0HuDfjfSqniv7y2DJ4A6RBIS+Ro3lsRc//bh5bj5mZ/t
0DNpBFXVkcHYMGoG03W66uh1ir929EEO0NIlbJRPoSrFAjR4HXmK1ybpn7mY2IhR
5GmV95sorDM8j+Tnglka6cwoGbc720SCrNOeKXrVscMC5ky2T8oGI8lYRlc0wOch
pxnWroXd4Itl2svphcNdpWgfS3ti5g1KQO3wnJBLK+5DU7d9P57F7vU9wMYamBRv
KNwysI8FMDPbfj4iMc3Z4pr1r6e+BIQbN7dmduDpYVjv/VzJ+1swJ9fP/0ZTehTJ
dLqnpeTkK9jaUoVpvt6o+QKFqA+z1PDK0AWBEkkAg3WaG3SyEyvmC12R8JsIQmI5
yVy7DzmPJXsgTALyUHNgR5QBmUwF1UTRoCN2RYaFLfLydlnUxq5oOhEiy1mM1Nym
fgrWMZiCJqQoQtb+xj+M5osq9CHm5ZSrCmIGgaygiXaUMGgiU+DDTq/gt/c+nhI8
ZXLjKD/MY7qpWQQiq5UwOvFBArZE/FspwrZ6IXVsHVHLBMf1mm0L0JIAuB6GWKZm
ERZWRZiqJtH2YbAnwTFToY/qKfdBTsw0rk/6L94xMlI9swIEaAX30m0GZ+RPxTWa
14KjHMnAqDBGFwyc5SzJULs8FHkHDGgu5Lho2QvxmsK/Y8YeEhvauL37ygTkp7Gn
RtMjwWFTHRq/4hwlLKgJyTXRTZvUr7JnG6IaQpEnLe3m8Lc0Zeihz9RmT6L/u2++
/anRQL5PZWJ9J7e/MUfct69i+NZo8is1y+QHtYD/pa/eWLhj2CXNtRzpAvoAxqFk
1RaQqwMePIxALFDOgRVwWtsakdTDZdHquKex1/xE/a0FrPZXa1GMbk4rOGlvT87C
zrw+JtDbqGiF1PoYa/YAk5mIBMgnIwhf8NvpJW0DssibUDGo7XHF90GY9BWRf/jf
2wbk1RKHkRA9ae992Qk8WYE8I93XOfl0RA5367XH+m/Gut8HDSs+Z7oCtIBt2ozB
5voYJXG0rO46TchXdo3vwRc32ukHxMp6gvHSrYhQmZSI2HlEcczNulLM6M5rsIhp
Aj6hrwiACQjY/OaLXvEktgYoZWcr7YPwzX7y5X+73iZj3aRrAfhSYkpLkQhYFjCT
wn6Wd3fwLBLNiYp1jxBxFXZPXsX0oWRlYuFTcbRK/jlH5H6ZpsOaIBnI7VkM//+j
bLkQdp4T6GpOOiADzapCS3Wht6rEDsTm/GlkpnJC7izuVPQDOt/x3ljdUJDEbuD4
r/uZyJYPPIPkyA27bycd0pRBRy2I/NhsFPxgi1KTIUcPavH8PpUMY6Gx/GG+JlnB
5NpootoA/bfS5jUkbx7Uu1qqwGr+aXBculsIa6doWYE2uM4R05wLJeXCwudPF4/b
QoK0AUXBrgHtYHThibo/MERDEmHsUZg02O9IT8aJ1IR4TN2qQTvM5RGZh+jwhLl7
utvvSWjfHIPJuftKDfybDY11oZuTdVer39lyWRDGLD6t26sbM3srtOKY27sZEkYB
7d1gVQGypfmg5MyutTRTPAogx/l5AJ+1LSv8oKZfVQoe+cVXg9ZT3ZVCuzCVr3HJ
nQMqC3QnCxzM8bDvwZr/WQK1w1fwWKdaVrjAN860xA31q4su7Xcx7PblRsJFwxIs
+Pf66W+vlkugf+vb3aF6Wcu2bbPKjbhJJP7F0piPQVDB0G9QlSgVVjr+ArGuybnE
ikf03nVP10aQBJ1sxDtCAANCtKniXNJSpXTtYI3OfQl15rsQIvMpy+mTbUmpni9Z
UKP5LwYcvA9ZZ3JIiRf8chNlv2sGyxqYWkknxuql30E0vZ1dhyvsGQQ25e2TpYFy
y8PxVc+tPAzcN5Ip2xEsjZV6p3sFrUV8S6RMg8aanQLu4FNr33mHOTR9IdfN7hom
BSY2kZrIQ10mW/zfJP0Ar7BjpkdLFhoEAT5QzeOiG9Ye2hCH2HvJQQA8mjZGb5EC
En0Vic1T5jLTCTvPkxIm6/f9Cohnioec4/FPC8yE0IkqRluy1PX4zfv3v9w2pO9c
03bmrdp3IrzWYxwovnT77Xns5MRce5cHSJv5HIkGyqaAAzUnHAhlH4ilCUDPl0cx
kDvQlXrixg7W6nUUklGf6sEEhexFXC9Wqb3ArJK92b5Nx0sU3/BdyKQ+GXoRVon9
K0m/yZ0GY5pBmgHWYf3GHJuEae8+cqfIKg8EJIPe+eS8JIaxCeizza2GI4Z261ol
tw6RdUgsVlSn8pzr84kQUHm8aHGwXQNTDDBxAIj/1Rd8AOil72gyaufI9ozI8dsI
cQiV833o/ldC/dvrlGSEPdODO5W6RSOZtSjbQZ30pyR93wMPGK4QxlhopWc9VKhi
Jon0a8jlr9tFVB0m1PrC7pPKr1JBVcEkvJR89gXKdTgEiPH/t1eAsTbeckeuXQ0e
BvdkM8x86mpvR/atbr+rMV1uggWPEy/caughO/s0NQpvl0Yr5YEZdhxE/rq1/12C
ztd/iSiCDbWbK0vUCKpWjxnobNFcINzzpMTo4AJomSb33d1y/4tvXUKN284J+k12
/c8xU40pmcacj3nxgeuA7zplU1mM6NIuVugWrCOrLkLVMzhvVsY7MXFxBeM3VIEI
s1geHSKOQBDYpeqU/JKpwp/HEbJ2/NZVKMXkFKuUnIfT15hubeVWslCnYcaJhDqq
4AgIkgSoLfWDVzQYsaAbqmgkFSkuwULdbY0j2Cwj1dKXrkuwPnFvFkji6pVVcsP5
yHVwHUl4K2VfcmjcLjgFRm1uBoLp9EjLdMQB4VmwAnmUn+jmo3pYs8PSmw/rJjAE
GNmbWnzD8k3Gbz46RRMxzh3fMR8InE9SeCDx8XR0mhEEy2MH3lK0/mgCVmO7PFFd
qvEbNkWYcQ66HtU2oeUuF1d+st86WyTJfm9kHDS8fs3xprSXYH6sOEErhC5eWh/E
d+B1EYmMiVrefsNb4QRLE5AsloHIj09k8HJzkNGO46FEU9ThjcIiyzxtJbIMvUAZ
gx0PECqlrbYDvF4PVP5WJNGPgKTJRJGBgvnv/6ZhmeRqtWmvHVdVP4bWg8R9RMhT
m1n2kcgZZ7K2e7Yz5s1laQJH0oWUENBjR93ipKEXu3D1uUCeI8jdcVaY9aDJHe9p
oS9BUjlddS12jNd4Vd5+YzZy5rbG2kSG1Bt7d/hvCoOB4ZB+v+n1rqbfSaNKbm9J
FL5Rl5oO3nAb8zWP66bhuSTdX78Bm12wfzRLp3nhONpfEZaFG4wP4QFDjcXlU3sB
EDpckoxYLwFSLn5WvSSX/nG6jTJxgpA9yB2oPjCCICkmfYmUU4f2hVH/PJINub5F
61B3fgSh1ZEekLb04skGDa8V9/hqqAF0+cJUMyl0rN4FTC3u/CfqCKHpZn1wiRkl
1RphgVWNfNczPXJk52S3OZvG2o+1Ud+KjV3a0FIJQ8p2JNNs96QLU5doYD7F1yvd
uryi1l8lz0UF3FWwbZA+826dyiXWSX61M54f4adRC7uJmLF4Lq4aSC3KdI04PZBc
h93t3K1SQrPnS3aLVJ8HxiE6Xk4N7B0hc/AFvnHF21lRqlM2oYnRlFC0EchW50LC
ao57xH6zbIuEwIM4eSd/ziiMpjSUzZnzCeuSrALBMaKG7rbjIEfF8fNOEAX2+UBo
oCgoVPkax3kFutfMdnaL9504SX5ADu6BNSKccidIPAP+86yMd5060yryp0QMugLK
B6nlcvAU4E8zZxA32paEBB0xprxJuqgtTbG1kbyZfWjsA8S+l0cjnd+jqT02bRsp
pio2hplTtzCiSECkPYXF2n4oc5ktteZBnkJl5JWwTvXfNH20Sbubp3jqU4wm3G6o
BzPsdpPHERYp4X+7HWox/C/UlNmjF9xWmxKC+o5KnfCBsum0Bk5dqPfp5JPrUb5k
63QVHzeOWafTYCHouT1U0o5ttVTKcZ45oT2MLGyVKjCdmUvmh0bTD2xeaIpVKIhl
7JWyJg7TnBMpFk+WXqIx2EjM2/kdkskTvEfcS2us4PkSTyvz/a3QjriYGSe9vJjr
vhEojMCfmC7dMdyO8ueWkmU1yV5NUmIjuVWBPAcYL6RLbVGQPTiunqnwdijE/uZU
V2NDiKOTZ8W37okdy7yKsyGvzU6ZyuPxp07Mr5BCjmctbyo3PnxMzOtCEOBxK9jJ
ryXrg1PY+HZzEylhqvfuxvdU2wa0BM/XmcgkRyWG5kk7eBqUhtyzM5NbxOLFDLEx
b2pvuAo9pInlB2ChSqM3DqbDItZFTbZSDzZol3CYY8YglXngtpF9ZKMth3FAr+qP
xlyoeWHhk9Y+hb6NEwNIFUGKac/U+B28b+b2/tKFZrtykPShcB5uXFDHfSMgVY+8
dJPcxkpMLgXDmGwQpVOQgPwG41wqMttwgs3yeSuio1jaQjYKNW0L0GQetwPzmYBQ
ZnUfersx3W0OASyfGA8zBUYDFc8SnIJiiU5bj5YS90ct8bwcWPaC3mYdW5WCYOoP
u84SsHPTjXdIe1aYm/HjQNsbv1j2qvcZ3mr1lUIVjJ0IvrH2NqBAhkt5Nej9M1xZ
QLDestPTPArWJ3iWMsEz57CiM/QCa+nh1QhmKNXkVryfBTLSXd3GZOQKUacgG0wo
vL9V9Iu0w/IEyvLLbABzJt68H+W8ofD/MgJNHlpAciFL67l0+/J41tZZJaf+EPJQ
8vivHgGFPqcVxfCp4loRKquJgg9dPatRZdMXUXrrhuckF7if0L6gcoqxbg1y5Shu
T5V3hu104KbdihlVfo+uozAFpOkHqA0XVRfhk8kFn9p7lF++OwtUVkSXcTHL/1ea
W3GW28VPTBFJLJOD6dzkKAvQeeDTAoT+A4S+2QbVoF8ZJsEiVD502bGksPBuB4fh
t/wkn0plj9DiUMnNX65cWtO32RGuBquTJTZ71XljdZj8ubY43lsqATKx7my6mIQI
0Nnidwmj6h2yDjCSlubLCqHELrihesbBStjWQgggF419J4F5US9yEytPVNJdz45K
EuNm9eX+9zRY3pgSbctc/ClGS53YbThyX6ftvErAYHvjxROSqX51wzpGTq81rkeC
ZzZi2HOqIxvkoOtrM34WDw4SHmlE3j2K23hWjUhF+eSLqbmP56Gp+XVznNWeSM25
4RDVJu+dtsgj6yFXg3GFDGcfw0glN910whzsF70kmvzlfFgAPjTqu4t6nN5Mmj/Q
3DapQzS4DSAhhh7JwMmk7xIKHa9gD/H7Odelp3A/J586Zijg6wMqCseKW4BPiuoy
vq3jMaD7dOqed2RTfwfhmRT6t0jeXXo4+aBRefk36mNS2x5o4l9twATcVmeTGRp7
5RzwW7VRdlcEv3g94K9iDwSekiFi4DiOUyA6zxPBU36hnXSg6+/w6U81icYKwY2N
3LIRbxpBregZ7pVVilhI2gdjrpH+0zZvoa23yKP8nCuBVkkhLDyLegSotyDaE8xw
ZTNR8iY2P3HC0PZtU0bvLpUatbpj6nY6YX0N1Wv6Fhy7w5yTfDcmF1NnKKdD+RLT
lSUHMRetc3ZdntL6b6iiwql4UymFr+FtUc37uEq5J0rK8N3szKPsbgwAUDGv8VDD
glUrugJfKxnK8lOktXgcHqGs8P+ldk4hW2/6YLd1lJ/y1KNQdaUL3rowrb9Xd56R
xJ8IHmQjfyRsgDoQhkVz1aUwd/ZT0jL3Vp/8Q+VqKVdohhZ5G8zYwSkoyQaxKzbt
Y7f5GWkKwF1CXzOy6j/92OlWNViAwfvFSMVhd31S/qjdnPJfiMsjI3+mFaJnwwH3
wWPRfhNMdhiiUkFMFbTMB56Y/agZVmmd0C26SCW40SA2dMhx96WYWSfKCo5dgL2M
0s7xbA8WO99BAjB3QHiMDHxcwPTthZEPTMDu2ECYOBlRnlkFKpIOXVoI7dNeyIhW
iHHjXBZ+Z/qfn2TMBcel7Tr2XouRsiHp1/LaPARUiGcMCGu0WSxxf8ZgNaysGBdn
ttRWfbU1CUuTcZvpoIpmVJjcSOil629jJuPPnlkzpbDOW1ebaWDd6vo+40nWiRyM
4w6SAKVNC7JVmfNuRwzItVglDfcggk9G66kVNGz7LiqfnEnZfPGGzTR2Ma4mye7s
bV9vlSCY5Uv8fSVIdAWZWRu0cIIavukDcKmlt6WGJL9aGtTAdZY9WNL+OcTn8s0S
apflvRXcOiwf149Rk1TjbnompH5XlDkusKk3WibHgFbpPq3BVjW9wqoLvJGmRKr0
5cpcyUMAvfyHtLSvqm2K2L3Op/GXfp129nKTs3feDLPgyT5CbKZDEbsvokkskv0E
dRfjTtIk8gO545dH8zHgxpheganeFNj/ypwAFQZQC9tebLJUP1dWCJIK3BCMcUVY
qdDZ3Uo0P4RkfvMm1HPpC8QernQGrRwX/UXBO8Yye/Xc/0G+3pexWHTYjvmVmR/C
mM5vKrORVg9oU098z0GT3qNE9B/lHoX1rpcQOUONSS7CG1Qd8GCoYWyaCIs5Fpqe
aanzG8RN5O5W/As8V7NzHx6xhmsMjjPfVolr+5s6FygsRkughHWo3/xPiZURYSik
7hDXVU2o4vAu7bGitw08OoEl+eVeEypyb7LWxsQf8r+zMregMfND/ZbTfNFNFdaF
REsdgoiBeM/hzmDl9j2N4Bd5PZFdpqncUabt67JlQM2YGiJmwm+/ENF77JNTKdZF
sqbTjHlUixb/0AaP0czRRkt+/WZGITIgNpvzfZwhAmz5uxd0O/EM5keffZVk8rIK
giXWM1fyPRBEoDPbIqq1wrOb6G244CuRuucALiDQ5Og0wYYVfn4RKF74jwdBOzM7
G7x9XWRSdxgisOZPDAyXQg4PASu9axG2Z95wHEL+whSyRmXPRx/7nbgYwydJYb9t
K1xm0rxRHmE9M1l0rpy+dxYgQy5VX9wSngZ+6HfelLe1Ta6iMbJed6efJ42hYHG9
RPTHwGv/NYO3clkiLVu0p2QdcYPdgzvmFKCdGInCdb4hasUawNEsUhELqWnTu0oU
TH6Gh5regx4EvggyvlyWErfzK56LhOKnrMpTGD3dzq5gR0K9WNZLoXYHu/aow+mD
sa+5BTqcNrHI87wePBupgnK5MGDsXTj1sVOJiXPeoNGAzbMGQQsaCBUbJvY+sK5d
cBkKegb8FhBwXyPEy6iep/jUAO3XAZdp3PPj1PhaLBVYSp3sG1HcFj8/ZJ2+32BH
pkUzhKuQonLOz5A7HM4afJdxRCA5dDsWdr2AlEt9htarBJ6kvcrJ/cy3Tn2tHBkg
aY7cdKcVOE2VjYMMinqHs+0BJON97erjhvpS3wG2+wNAPzH6TmGE1roJClkhQJ7i
zFQZBb6mQ/+BpR3nebxgt9LV+u02VghuBf3Gk275+wzQ/BSKopXNhPYwN2rwZKxi
w+3f9A3+UMP42kO2492u5R2uefsEOl1np22xIzaAauaos1n8GZ5r8k9Oom3pXuV9
0k5BfCMroQhPclPoAqkh/gCV/k9wU0CIgiiv1GoY1FiG5IwXo7Rn4ufSnJIK7Iq3
mDI1oal7WMos0iFzO5IC6pzT0fjec62QPGixlSKF1hCGX/Sv8A37CKGoGTjwXZ+9
/yCo+xbZA8FPE6jSyZp8K+4C31lvJlne+n2ctdahcx3J3PcHjLYGbT0R5gSAQaUs
Yvji6PfFdg2NTvcZa9AsucsLOiKgeK0EVKqkelRgYc3YAmosU5hVCjSGgCK9zkFp
UcCGv0eEilMTjOMoPFP3JBUUhVyIWi9tYf/U5RfA4htN8Mi9DAhiF2Tx2D8dXPlZ
CHB6a5150zfK/vZPCPDss/45iYXw6/4DRPheZ2yLRiPdet1poyfrnQ70dhamea8j
N4tGI114yM/bvdgxxb2gcZkkJPzZEFbQXzhkLJvc2dZnSxseovdi8yADM4vr3/nJ
YmdOFjPK0kf5ibsc3AwQq6iDLPiu4RmZ7V46oI2jhE4+7eShbF7OMRoElcPa99MP
u5C6kgOXRxidLJhZ9ctF9RHlN2+nUUnAfLviou5OvD85F940YBuVne7GZv+68iFe
uvRB7o5kkaRxEL3Df7mFizKolQ048S63rYjh72piPef66uicXVo+sLIQtIAceQti
uPMlXkPxNcuf4uSbRvaR2acR8YzimhDLSyIRzT56MWxVhkC9E4yEiaRseqQuzbD/
78/NHUdi0rPO9x6SXj5FfTG52qbtrqI8sXzzE6SyI6/HgqUJEDxyfZqUsnUpo4nc
KOdzuUVdhsxK4RLgqFEW5tfgks15gvzKLnHS9+zQihanJ3e0d6cW8D6L2aFIsUxi
pbeG65VcFmKnf/0xD2/glSuaDOqJNaGjhaWgN9rADbiwYheGENMlSi7WhnAH1B1V
kkiOU+0S7haLJoqpNDuBUlpzL/WFVjJ+sxatUeJdog312UVA96topebY3aF6NBl0
WybLhNoG7Yza/bCdSzk/rLyfVQ346fq/dlLfnuw+kt/GAvvreCTUqGZmUTCoC4Xf
q/nMZM80VaaupOSNp6dB9b6KHpLOZjUtXEx3eSF9vHizEg81vjVOLVsh20YVzlyK
Y7W/Xwed7Ge35rN9NW5OxeS/UWgzvKb7Uu7qUs9JqT8PagJlPiQY08pJOrk4xaD4
nU/zZc5ZZ2w/d/Jp3HDlTW7XMe8Hv+FVU2xoy6+KNEE1DJFmTpkxNmDaZGq6Rej7
yN4MTTV/3StH98Ha2IeGywCWCadL8kpqPGUNzW0g8/8Mca70IlxGC7Oz9p5i33X5
yXSvuy64E7tbktjCQhfKOH3jUoVvnNxHWlJqjrqoeg16XHAmrtRXqe6JeKf1u64h
MQlJW3ypoKLRR5wPTzIDWjbPvGIL1pe/m20ppeAzxDE7nnwS3BtoW4KbMM7ifX5y
+wxBgN9RmGKFKy1NgmHHhS8sJZTEhT8mXNAdHaXKiUVRdqjayjoZn02bh/K7g4zl
hwYHt5DF2wGKVrajBLumin2IrBneusNfYgPEuUKv4SvNxGdEWJ208vNufSJRpyEF
4/ugqN9W/nzOtVIwhKKvLvORZ0+FOY2ksHUlnQWuwKLQ4rymLEFjZ4SsTLm/ltNh
h8Pqafgc8t8ViGN/gyOvgfPQNkZ4JdZAUweoAvS84XJIioycsMC4JgvupYH23749
zW48Lg7/bMnJncoT+8hs4PyreFyr1c3zKzBPzKFP0x2v70DluK3Sf9wgpm9R3/wn
6sK7JTjrGj+7lGKe3IP4L/4ZeIJIeKNfeVkNS8rWvyv69cDb3KRMeWEREdpZKQsM
5vLtcN3F81dOxjBYon2PNxy9Vsc/ST7UZFRUmYaJLYnT2XvZ0rUU/V/XSf24isOW
PS+mk2MEhKO62jJ/eT8FnsnI5K3OO3hrVocaYlsamwdk1F3fMBWRCZ7gkwhtfew0
lz+e00TtZXit4NuTrurQZPEdPbbnp/dTuH/lrJgpZgZQ6+Ytg+PJyEh8hm/rWpQA
7WuDT4nGKPuEX9vtGOe2dfjkkD6k7u9Y86ACPEJ+W30TMh+LVA4Vp8RJ9mwVwZIb
LBk6m6bymXdxrvg0jZYrIiHSEhCP669qF1DgoeCCIj85DaUCQgr4qaRUIGZUefVu
BzP4WNQLP6umT1YzaQjub+VDcGfTE1nAoNY9rJauukxjH2256f88A6U42XMqDM1Y
ev+gp4bkmFNyuAa1Lh9+4Xa5wZ2owEimqKn17lctDhwpsOXAOPGpNAgyoRaZrmJc
DcX5Qi6CnK/b9NEA3V6BEYCUU4a1XcTaS7610MO/nHBRiCT4rI+szPdh/3kqMqet
QqzsUsuqNcis+v1RtE/bIeG5krHaAcMA+jaNL1q74o+shbS8gQPYjXR8TWgBE3Wd
pzym0EryKjwpRj+Qt1RQtxq+PHJP4Wy/rPsJKigDcZYcKvHQ14qb+MhQYnRPKMzr
J6XI2wQuB63JjBRwGiXCwI51sz8YNUPNxlWsmyakyhYGMUwcVAUkusG/MNkXRQZ1
wPTuHtB44jJ4fRucJ3r/awpfVRRPn7GQYN0x+KlLnUcjEU23+pdJ8NFDU4qCDOdl
HqoR/0rtGpbGVPVVN+7qbDdax85DvsNObdON6db3DXXwPRXaE5BytmxFNjnbCvio
wWPfhD0hv8nMhPg+TZ89qMLhHaALXSO4mSkyz5oB5ecP7uVKrk4nY08DhUpGi/kx
oxMSiL5vMrefklAkR43oae4UxaY1NCJRd3zUOpCwPFM+w5p125s4qPBcUKa8ROMc
fdv7sDm0fbiMgqUYL7KcLEaANEdbGb+no17GaVa41S6ZUhLYpXX1p8eUGCopGRk8
LY5sTyRYnKlnCTnFanD303nU3hhRNA16E5KEdhK8hqB1O71sOYeuj+aUjN3dZpOm
TjdhQ5i8rNX+5JOkqnPWaAMqb/knp/dXZrpZZUXFvpRDHa8Mgmg3J9ezQsJcFNDt
uxyqNnGQ328Vau2LQxNPOycDoPFWZ+ebNgHXj6c1zZSbsmlxT/m4vNL4AvHDT5cV
5e5HcLNd3XzFeH/EWFEHMEq59F5T2s7rNNJHkX9q62Tpb1UH7pUGjQMvkMNAue1Q
m/2Tak7MH+q1c1QpqO6AhV8TmLdRHyVKaknPbsnDOdx+JsnebEJGBv2gEEyas3rU
3RPc8+GVgqjeONt3AxYrwSjF6chJMGYqLYCKTKHw2AXCOI+Z3ZxmH9R5lnft06Py
WZWEJTN6mFcMOS4+cTVIIxgS9mfrZqFLnhcbAehvfKfgOgqr6LDNpQQxmFVSMWM1
GYsIm90rDQm8Mt+SpW2M8djjNQkLJ38nyA6PDxEvwHxywfYA1Iula0/dV4XFEla/
D+rJOuL0lwFAt9pIBcjou9mYxdBwXfDE09Xh0fJmP8nT+VaOdtm5wf5p6u/d6YV1
h22L16/jMV/N0QzBK406AM6R7KermEPeecyHGObPsSF4zp+8NeFx2sbPNcoX26AK
q9aLoncRZ1zvPv35so9YoyIksjazKn99qEYopKQ48Ej+4s4yNFdROlsqC4IVAhrN
Q3rwBGv3SFLbPry9FICBufYdIIXGOfr0XEMVfCefrwh1phcIl6bsLavlwRLfUlKi
pGwtYjArPNTnKFuUGS98P+sAw43rU8QGLKs3oELfZknkY3FHxTuEQ+3Q9qfnoN2v
mAPPoDbMdv5SDscGc3sKYA5bEgng4LtI2PENdqoen4ljY9T45EiY4RJuqjGJo1D0
M/JYzgc0oPbeTtJrWATai7Ztmis4t77zSPmoYC722vNEBWDgoYp8fkN2IuepcLuG
R0r+fO1LWRf2ghW9NSQHLMnMniApJMiCvjIjxy6HrsFXspV4yOGzB5UoIip5wkaN
L3CRGEwTeLODtKtccdoF7ZwMGBJ/5GoE/XswiZMXBIchE2JOq198ffYKeYW8vV7n
fFs3WgDADhW+shZQljIu3tE/nI7U+7mrf1PNH/MlIdU1c+in5ib7N8tb35HRuG7t
H6wrxoXEZKTNAwbTPi0+sFLsY8MGMe/jHALKrLLIh1uLF7c7l6jQSrQSGwSOiedg
9q13zCGTda5RGtCM/OBQ2JVPxwPRTtb5L5JC+KHPq3s77Nt249C6+Q9Lw6sig/o5
uvP8esgKA9nyrsA9WNmqfibB5xvPH9cIv2b0VYdKjo8fTESpM+6dK0SpwXkPDd/T
N2gqn5LGrXGZRYb7n7FlgYS6Bw++miB11Jy1m7Lt24UwjzgQYlwTJLkzIr3q/zHO
3m5ig6scQbD/cNI/4k58maaXECSBtwPnCRV5Qaap2ggedXhLpQIYQ1bl1/yA3q2R
dEtdJMw1bFhEgVQSJUBspdGuW64JxCMDoOhEYeIQr3adSVtqKloox8w7nqCrqawv
N2JEBBvEd6/SmYMoOj6u3OE6XJUMZKOF1KOV/jQT6OGgm+7dgP7/RdpwTAyzbBbv
mjIXu1//66pjWAcz/8A8VHVfn83IE3v97RxEfZ8HBmucHl4qkHIaADR+W7XC3e6g
DQ522Pz63aD0CDD6LkhMOQTqMjGeZSKukph5gTCN9RfKCIZuQTbLOEZ8QXMorKA5
2UflzB6gtjL893CtKD35zjJThspI5pO98WbRprBUzFP0bL/16zQW7wIRdTSi8jZF
ED8CzWjrVYNo6lOFsY8IRLcUdInF1QtilLpnDCdEU1Lw90bHVEKjsDuKHkCTuLFx
XMO6sI52CKF08tJfmV9XyfwC9jrMj1CS9zr2tjRp+tM0AcejeyuX1KyFemZqAdMX
Ig6NVSA5GW8RV473wJa3XSHdT9bfzgZM89kx/7Zm9H0Ke5T5McPrtqFSVvfIadhN
F7dgU92PlfL0cBbBF9F9viSiMDUuMzxANtCFwVgyMpGid3K6uJJ3cPZMo8q3Av1s
G3uBedUySbaAH0vs5xptazJlCEPb7mKrhuS7xNfBCE7KbNsZR7eeL5VJalwmskWy
b0KP/rDE1FGC3eAmDjh+xh4ulhkQb9fBnbl8UUIe/3bZRbymK/r2DfY1xpxIP1JU
4vtxlLO7HgoXQ7OF+TXntWC6vTUf0+Ev2r+l6KI+NYNqdlw/25Px3QxMbz6SIZi6
oVDHIeivzM9G1uOu9FcEAxk/8a0Sf8AFXmcva3TUysU6HW6SVsWvPFzLqvca4lp3
usoBl1MMaA8T5nbBeGCBURJLUBxMpZknF3EhiCn9FzpJhNqiwVfsL4vfIIB8KBRc
V52bvdjrePF4CGd0Yzq6aa+XLXqbWpcmy6I5Ra+GSkhvREjH+po+Yd+1SX8dkfSC
KX8eI7Fk+YioloL+2rje9rbFogNHCO25m3kSHdsrhycTJZkVN1ZCKTae7plQ1Txh
iSW5NdMOYVju+B3XxJJr38WRNDxDT8xDoLSSzI6p1SPHvZ6H117+wHxPykUHFuJ8
s1XXIkPK7VvZYu25udJkIwbKJsupMttqK+D4fv3O2ML0NMR4RG9a2527Ivj+m36j
TB8mtyxt92v2fUgzL1n40VMfD14zReJQNOFfs85aH1RkwR84v5LMAuaLPeA9XeiQ
yWENUKJYENUBWq+khL0q5BQoyyw4A3LA/DSRCfCp7UF1a7kh4wwGasDkMovEQDDY
4KCtyrUC/EzbSq0A2x70mSxPrDKH7sfc9XfNYca5p9LOygtmBCd4b2TveoFvLlfs
Xll5UjjUJ+RGMPFud3CX1sOf0zD7xwB0XFVY00YNMPk6VVJ/QkJ2sXP9KYZqy1Fs
Fkv1zoEAizGbSk6dRlddfJvrYxzdgq/Yvhb94uaLt6pFAD3TgnKuoKKhwlXmrlxH
FTXrNRwdFs1y4wSkS5BYHu/Css6tzxrHNNXZACQEXSfgJkN1v81yCwvUlsDJ4/Hr
6MgrBhRC0/fd+OWlSBOcnWubNRPell2yKBfBSVAWUEVqW8Ktgo6bKn4xoaDIpJb3
7fwoX4HQ+K/JsAlqKicegvjrmZfzIUiBsgWye7P4SBv4jh4Sh42x8EuRVIoy3Zm1
kdp/afnHjvzOfEEqC6YMNGmOlh9iflqmjOcGRpd6ZKDmSpil0IUYamjvAWMmvKgf
V5K3Jq0aLXhAY9HcF/RQcBTedX4QrEa4iItl9VFRFmSUojkok3AnTq8N5AEndqUV
WYQISdOJIyo+9awx9cFNBktcgOA7uPNatj9vJJs5JItgL//9Rjf3wv1+nJZ2RYWN
5VqEwNSK8Ed1ZmQp6chtONQ5uqXMryIxu0nqhgS5snM6beqkzkqtWWi667kbo0VK
sCQRXPPeSJI0F8MY6B0dJCxLBjLsVu4rlGodCjvnlezBA5b2k5cH+bfaqFBlMwlR
GGUJ8XYs77+bZP6ifhVy/Cr0gKn6fTnOPrnlY7rbmUTvSDqg6tvLmPOLn9f2NtPW
Je5fcBqqLwPQOO/cXdOqLDecCOvIrPK0xArikEoefuNRCeSY+LBJtuWbqc5+Ph5t
Wju1OQAxdMplGruhwqOdnx9ByaNzEvialIK/kBw+eE4bNy+hCJEyR1sb3zGzFGC7
BEY7f8dHU/bO+J/UONgBsBZRdl5CtsWeQae/U5okB4CtfrWlqXQBXFGSi5nqgAxk
Tsp99gS0tYLYOpo7xHBmaomkeOXpY13PU96cS5v9RmcgI3mMQzw1Virr+RbsM3Vv
Px6y1MG/HB6VoQodaJksGi37LbYiWVAXO5Qy5zSduWVDLqIEGIlQYsIbrnmQI3LW
XMuNNoIiK0Y//zPKRBMvAVNxQCTpa5r+2qdyo415OskQQmbK3N5ZVuTuc5IbJM9s
GT3oFYAH8PAlZKVBuxSsKmF/H3oT/lkRmF+WGKOyuf7BHN+2wix/T2sUcKDBy55J
G7UXuEKgCp5FT2G5i1WAVmPXlgx3X03RpNYgIGw6S1vRdQuTgwi0+5QMHoNgW0u6
/ECyVWTq6tS7Tw0iVLPpajjhXqUgHwqatNAwS3bgjOUM6kjowCuLKUXMmTULRD4F
4MhKzJ7KGWVorh7ukxBzthuzW/m2UkGk515DIUxsuwi1U7r5NbM2kub9qXswgsnP
UXi/+G5iOP0WizNIBDsRAgvY0FpyajQ7YlgHJxg7bojos6X0zWetBOlJGl1SLCPz
5U07xQ/pW+GD9LesUsVljf5Nxyjuopiifn/Aj4wl5vcrI6qp1x+qm+N0tWGzys1M
5LqiZPbTCAQGz9K4xvOs6VRWKanNswbmZCOqO87GJtTWAl6oFHLpFyZdrXG6E3nT
9UcpNBjxfQPQcZWVHvLTjSVtnf5ZWS9JyeEkqFaoywtb+DkanCxpQXCEYrsaN7KI
wG9Wl8wd/mbG8R7SQWxUm7WijBU82lz15VlEBT656z2dmUE+y48P9mqUcuLCyYMC
NJWFbdomp9ZMvOJFOQu2lDtQnqkfec5Sd5V24ToeSa32McgEak7t1BJYrXZRfH3+
g0xVlBNDFyYiuLIibGttbhPH2YGHad7aS7fAeWxA1ypblKSPU7zyQRw7dl2tud3d
gV9c6UnfOoO4d10ptJmqoroPBzUVQ9aUUJdCDHD8UdX+6RArqDl0RKYzs4q9W8za
Sbby3Bd8Ag6Gr/tGuPGVpzv2WyXVmeDRLv7FNy+KS//vT36yIaSFr0G2chnRjHzR
3cxPPjxUQzvTdPXyniahDegSpaRLEgkbU2gYonbuHlhBonI+CBh0b8TZWi9aRY18
FI3t0deNzK8ney7Ly7LEb3ooFGVXqj2s/h3wOH5CNGNQAiJqEdpEuBN5SmGpK9ef
RpxAVW2Ka7ploPeuUEALG84ry3DmnOktcY4IJh+1THNw3Na7FnLAGVErXt7ilD3v
zFMCm5CnJDEd9DIW+jU/J0wYkC6rYi/9vqkKY+3slp1KsZYX3SFj+n2rPkFqN9PQ
dh9ou5GxbgO6yTcpgIN5r/byn3dvz+eB6pI3ynDqf+mR7mA5oJtNR6gAf5hIoKeL
oisNn5bMWCHksHLBoGbnSHLXL56f8k0syAlGe6brs7p0wjDQLeLjeAJldeYQ5kmw
PCzqrglOcim5IQnSM9m4Qm+BgA9kQMlI1JK3NqveMp/x7MYV7nUrIcM2bwm/M+qO
CG1gBWqD1NkuTgICiJRLc2zhe+3/8/mYCMvj/iXclRNWMVsxtKH2uUk7ofVpcBew
74NXXfnDtiVInGnsVAtteCtOTGFycilpBLCkzyrSO6m25WnUU2WDX72fvRM+nTm6
8NbYS7rImA2vjAR3DUixJzlxZhiZ7+YjUrN55XntA33FPJq8/4kO3LWkU3VlB8VQ
/hvN5JR6+YJjaNQTpRcuI0L47o6L+NTqy3D+em9aZzVfsb4zC3o/6Wp5sOdF/5sk
BsBhXxsO1tkXYTQnpSKy2TezurjqNjNWzNnKcuYRnUlZiyHEa14/rKDirSATD3xK
mAx4E5aBqtOI7u0ljVlYlfSuP0E1ZYTpquDEWocbLTsvnLcn5alAZ9uFrzwe2lS3
8qXH1jld7u5F+qRNcQ8XLBdUx+FdrGu5mNJHeIKWfnlHrLthBRZDfAMfKwtdxDjr
P8tbnl6k/DE/9KjzvkNgLp5VCBTRitTp2vboAi+lAYbfEqtMhI98kydjtueRgJ5R
BCer+1rfvxd7B5LQZywVjZbJY0L435tvGS2qm0Y7RI44AwuAq6/pCHXJRmgA3ot3
r7u5e3egf8AKAxRb5Uu4z41CYdIgHrbZOsZ6WhzRdsNiD+3m00vwABGjVMgwX7rG
1ayG1tmDah7L5JSERL5KTWtf2l+VySuJX6qcFssacJQV+zaK5Bafs6tLaiO5Y9sQ
rPnlB0VuEhnBQbEF1DpIgLvJz2Yot2z9yKCygrImOAzFD20nITXU403lCzosDFy1
/oKzxkE2Yr3uVmpxr8P2djdjM2VOHOwsO/1zmZ0gCs7wZXHA6BCFrJX/eixN4vjs
WinuXZbbbTFmS04yni9pmgzAlHLMbfqR0CXS89VRytwRFnV32PokGRCkUCky0YNu
LzyKrmdPHCS+DcJgOr3beAeEpjhi0cqpeSOUza95AAC2Pbm2+GErHpmiZSz46ysx
ok0eUCxpCerwuRRzjUBQQ7OrPoyM7cAEHXbp14ST9SUHHnL9ak8VkFKCyhGzyM4K
E1Zdqq7cQps/yXHeMqeaC82czD9+j7QUgzc/n4pJ2ImGHYNdweVZ47UZN2B+F0qM
ZtM3/p8UCfgrA3KER7WutGyB33RfQ+bEzwcYeoDfIoREN1NUlK/S6jeNzZfRDQv2
s82yu4HxEXiUmBZkev8KqxMibDR2PoocNMnwS9NtF+Y70m7fxsgFw0NYIz6Ipc0U
6CoC4CK8dSg8SKm8KMjTV/av/e5LhxHg4aq8A7XiCg917wZ0CGnpUIgHMcHcMuPW
IPegs5bD5q9+GsmrfUY3+M5PYShDKTt5BBSI2CXisOWd3YVKHyzMToCERU9hIeSA
L6dKoxg5wmk4VhWh3IFUkNFrXP2vjXd1uju6REgUiis0N7tIIFuuSUMHJNikEqMQ
J5I1WoFjSz3B2a4CXuBVPLlD1j24j/SmOPocRouxm0uLJQieoNkBIG/AjJuQclLC
y/dK36e+znT4prJVl5RlfJsahgJn9BqMUXtnSLIdaAwNDlS3nStTyjROjV3M3D2N
ffmn6Yj/bJI1FlMl7s1DOtKD2VanB4tLU4sRnEF70f+AOgyYOncKh/SXsKHr8N5Y
SYPBG+wG+T31slLnAJnLR3Hklru0tA0qxmgjH9YH5o9m0PsUsAC7qABcD/29TfG3
VkwoyvyNx/d/p0VHJ/t5Xpb0I4cAM6NQ5LASLpzgOZhFD4fQ8ravnl1qw3uXlzZH
/t8OG8JVJOTdWCP+F4V3e0n4QhcoaUZEMBUyjGXF6dgDIYl69GsI/5O38F0fLM3A
oiH/miA/PlpFFP9gm4Xivc5LQOQH6JZTH9LLEr7sQfQcdUrxBNbCvlmNfkx+KZ4Z
M4eolZICdYYfIDaJqRHUKMxJSFLTsX4+tN6lxRcUlHuSCRhzlV5EuRTA/b4fyrqR
iWq0TOYL/ZPHuztrNGT4h03LZzGlkykqQt6+SEvFqjD7Db9ZGUWjsYAGgKfFeCz7
8xbccL2BaY8f9WzQ4/+xBjxWujKcFNdtzJqXduxQl3bFAg1ILRQKPcc8Pnl4kfGe
B/1jydxx173SwYTaqjL0AbogPU73DkNr32aCNytHJtwE05yr9+heRTd/rppSnS2K
AqLCCl7aNY5xhGnkc1VD5m/JbGjhNAvQIlhV2PegmUBtNuR4w4jN64QXzh5x+4zj
gOpu+dn7B1RB/5PGroM5+0kqzwVjAnJ4aGW5X/6xT115J0/KefNaya2/jnB1TF+H
uX/JVCjet0m8y/uxzspzdO4vW2uqQq2Tat1gQQc3PHU+Kt7rE3pc28ZATxBxrt+G
ciB0n86FL85umi88Shsv1Lrgc05NpDM3L7GQSWvx1+o/T/IY+s5EPqSUFs4DcjzG
yOIW8goUBqf7jcQftir7nk3OQ+QKHciXFaH+fQRitUW2v7BfR7i9znMTkwStXNYY
4Tlaqp6sH5yKGodidxvG3ptPEH3RZWP6K4dckkB2p1sX5L/LAZWuKe5NNMTAag91
7ldCQ5Rf2SMZfUOOb43v9KOuGJedUsU/6ezx15jY/vEi30vxp7m9yDsq+pOCwX0e
24NJzXfj7safgkJrEQ967lRRbjX3IY7E0b6/r48HT++UHVWkWoHm2q56OtQ8dmp7
yIWB3c5jwPLDySFtR4HY4WB3rpxwPFj7HKQgPOxdJcYT/gJ0nBE4LpQuyC58/hZR
ZGHpMxfhZW8GqenA1O9LOmWGLqAP06uHguCQGuZGWIxKgmPXK3tXteupBLbtSVVr
2A1X8PGc8Jd+a0gfxAYlE1ZhHeS5cNe1D9+GGvHEUYdV31tftRSRTjiNEnLuVrjN
mC2XT6oZ0Xl0iqf36FM7w8zzXbh+T7ePwwrq5Mg7C+T6nYwq5UFI7f9Zrxw70gjb
BI7Ghr06n+JWIUOysARC6LvPhaSJPdrLkMBZVKanBAyWLgHHg2+WG/ruPhD+SgLj
IqoGvfXuRGfcBo9Lly97JxwKflPLpwpMTN8DX3KPpMNbv8JQ0Kxn8sn1xUlQmdBz
oFkfKwK6yywi8U1i1GvPzJnVzS/7Ry8BAbJbXXbUKUzVv0RxrJnJh16JoCZuSxJX
CDii1T5voBKa0X+UPb0J8/XvwHCoCBtyyLaBTy+NarQzU1reRDxv/4aK3CSViCh3
Y+ev39RwXa69LmG05Qys55nVboqScq1lh22bSNvwgCUnTSQyl+dIEVb/fZjcnyMx
yTSnXKme8OWvJplaaw+CEAcgInao9ufq0K3yvOvTrSr27QubjDc6fAamEMJaQkik
TG90hjcwrV4s4CsKdRlJX88C1GW7rjYPYZ4Mn5d+DUb527YOuhmuuMn4vwEgFP4H
fa0nJqR3pLEguydJC/JBVL3tnYrGInUiisSBuHtJHvH3ZhxwDKn71uygZTW/OzO7
muC+CTJjAl5JFfOFAK25A7UnYGIio4W63ZAv173CBr01G5xLMj6Mmb+7D+dcq9zV
TPRN4iNNY575q9lVxBSXMBpO7ecE4k297Ui0my+CZtAw3ck787G+nA2dlK5T4rG3
0ndG1PMXlCrSozFwz90sKFt396Gb8dT2zKub6Bc5uRMjUYh05oyH6mH3ZBYOEPr8
cgyXtUSnEB//c5NretrExFX4iUl6LX2ZURqaVxUVOw/rDCf16H4kizdDGAeK5nfP
3dur+eQalNpNlujNNxS8797HchYv5VbwoJ9Jhh6Y/0ElKr19xH7l5mAm/vDFWS1P
/3GauzmiF8ydmHUGkZ31VW5ZjUQ4o/J9/6X3uVjgFiag9zA6kf4uVkciiNX0fuUw
AzGCNuXkQ1qNHVkQdL3siFvsq/b7on/vbU+Fb8wTqBJgulTyle3nzxm91V3PBV1W
ESr7FmczBqn/EVdASfBEZNFnTtvRJBFULnfyvlxE5NOrVDxVb0Tea9dCme/cfE88
znmEGV/NDZUuXycDx3FO8t90Z2VntIZy0TSeEg5/lRqC/HVHiTeyqWWRLbh3oCft
KRpyh5TqB6bVFF6tHld8DAyvi08FVv6VH//gZt9ig4y5p0u6UO5gH4BxPW8goiI7
rn7aidipTLRsA8mNvyR+UULYd2jnWIfEn1ZGMvPjBAbLwwVvXEtFMR22KOb1KBbC
aKp2LoUqTr7rU1I0+VWCq6lCenDIzzyIKFUDCWDYzEWO+z17kdOiPh/+Q66xaSxA
jXGf2C93RukR/2tgL7WjAedmd6GGIwGodLYapVP0ocyJXVRGg4f6ub/CURCtBcHH
YH4QQJuiKFnROeLYEfDnQVV5cvKAzm0Vf/JZAMLadcUbACmUrTtgJElwdIqZjwKc
1pzyt7cnnj/L1U+JGBSqLhYZy4xe0AUxZ1nifM2OgDhCsCMM0+KPlUef9dHGE2jO
sWeJ+zTpbjjADwgCBmHqBLGsTw7PxqoNeSOpGW7EDtfkpKOoWMX+AgOZfKuQVyE+
SIl9tl+P3YNHTj+I1GcBu4RBJUrfhon3wmiM0rBV/Iw+E2WK6RaCgQMdpe9ajzHn
dgU6yQ+8sErhq87t0zVJ5HQQA/O4Lu1OzNgveIiUlquSEmVKjBlDw+3cbLc38FUb
GhulO6dEtVnf1jQYUs9VOROoFBnK83LOmbWmN2pEaVwax7VLTUMWpIhorsXfzpBe
dC4XzecAMTISuDhuzv4FPTAyKrVNkW6AK35P6y/PRacCxl/nNMPRp+krXRZvVRsf
G8Q6vcOxfg0FlSq/FU26rAnpt+E+QyyqJAaqAagTUljnbAEGZsNCbWpKG/FmuXuf
8Y+42XQt7MSXo/o2KCOd+19teu2fVHFlHLScmXKBhkwkDR6o8/hOt4rWXOZqcTYs
kFsWfYDWhLp5J4QrGpn72JhpFQXaUvzfejD12zD/cETls/WQ7v/Q2sgdbQ+EVUBT
/XeksniE7wQWAF5YQOYBmdFibhp1DeZ/uC2BUzIo3kA0Tj/0XlA/sgkDmZjLWYQ5
Dm/Icom8rB88KHru2jnmI8SjsO8GzXuo0zwNGSrNloJBwsR+KXunBXuSTgWW9sWS
MNrP4bDKN0p9QKTOgg+AdtLgQ1InO5iEn3ijgq0HRvGRZB1TMPonCKXLizEg/YuB
z1rO6JQ0TQoGFLk4+rYgshsDpML8br4IcEBAybyLvwtL5DC8fdjLrLbWlycYQqwG
zlsSiDZVjSSXzvvbt//lKQf1E6JKpjVHidWtqUCZDWMswatQzDU+YIw7mCcS9n67
Iydy9Upwt5s5894hr4cBQ2tpXf+hRizIRDdVE4B8/IZw+yUSUeq4z3ADPGvdr8wZ
CinPknjwK52tz40OVhKvFpXowghzqUxU9YgnjzNorE9ypnvgquYHmWkRKRol5FBF
E/MgF6F70zVRQWvkuaouzF5RcYoLEnc2buAYE48Uqdv6h/hlr3pJ4TU1eaxZIA7m
rk1ykb8uGyQcdVHfGWGPJXY73PBpsYjZAVkGVj2SRqsSsNvC8Ua5zMpwll8yfQpZ
5fzlNx5n9ArYmYggkyloO6hRaK6PSrd+ZDfI3oZI8ktcSdXbbwMP0OKTZQSE4tP4
1Qym28pTqwFxlmpbK8efk7JLKY/M0ghOIqmt8nCJnif3bqToFqEY7Z7P5nRMI0DP
dkLinFgmdxIQ6384JsZDJUT0yULeNegp7696oihl0itB88hUPOycFfHjS9KjME/H
KDdvLdWheRf5Y0i2T/wC3JFzOmVOhlduLBTfabvS7YSg9SLmd3XpbzZOKQyTd/29
diIl8PoVPOa4AOhTJdqXmsIKEYU1qtCkYVNBN+JjutesoCC4ftPOzIMLwHwGaXXO
o3IIQjjxHKknit6qc7YG39NVvvYUhzeKzVe1A9Q7zzqzsgLF2Ne5h1exS91bAZSe
HAM5t3PnXOCqbr+LfNVPkL2ooPiE0gfHdUPYrRfMjoGGqW/MzexlRn71bMatQJv7
NUa2d5O5DJQzOSEgoLXMpdVqM029SyZJQpsLwpRsOY3EL9uOxgOBQ+pNx3/zkimS
2Ioaym9lEdu1vX917ijb/KqVQFrH56KQ+Xc4UoXsp21UEPABqEHOLK7qhursR7cy
v77ZfCZUFGoIOrLa1AzxsQiHOU23bEr2NU4yoocoIZ/co9ZLVR7W08XRyGY0Nlxx
yx/wU62zEQ+BqGF9RRGvMnSZwmPzok11ut0MwEXvFAegpW3v2kqakW9ynQemGBaH
Wm6PPLNmhVXG2bJ4rK6Mj8+IbBBbI/F2YuujKera/Piy5BxH1z8K2mT7szic0oRm
zJCUfpYanMj4ZnGQYoDe08Ui0WfTrkYdMI16VmNLAvA9sNgnFk5j0WED3SgS30j4
rEaW23O9h7zIiBZ3rgIXd4m6TrExH0KLUQ+Tzr4aOJ6hcL1wiHkW0x79v8HERGGB
KR4+gOKw5mtS9d+gHBMrxOkOJG8XVedUdFW98b/qQyjLLlVVcCG2EK6f4DNzWC90
7CQanLo0r81Qt45BC11XO0+lMSlUaOyGgGu8DhDzSuZqDxq0yWGwuq8kSLwH59Bf
XXJKOK4MEa2bDKjx1oc5jF982jFxzwKpkaJqKaY+pGELju+sAS0cHk/EOc4CrOBd
GoTJum/j7d6zTrBzD3+6UcmvnyZixcIzZNbtPIJ2ojUyckkg5WPBuh3NzoX2fjbX
asvl42nid7sxeqI/AhCihBlaLwvev14H+aIsw7wX2+c3+G8gvzmNPiyVYwlaxONV
WSubfE2sTPMrBc2bnQTv3CVshLH00lur6ljOpvZ5tqYlwltsfGl8QQkMsPTxz2lp
ZXgd5xbccCkOm8VERRycLg7yGmfhYBFOqNkDJyRKyfO3fF+6ghbQFzRCRwXwmMDG
V7Pqhcn6XwtIzgfq2ZgI3M00lS1rUekIwtg75sWB5X3p9cboyMPCMpDrDJpr361k
y1MvUM9feDCKMeNZYwJ0Rw6HcX8+rJANS6ONzENHW75kA7ivlA0JtTNPQOB9hTQR
I5sPvfb1B73QIX6AXALt9+2o7N3IhpnnxhPBznhnjymZskm6RMdZFyJKCXa+euN/
m3U4uTQM8C5acZFKKz4q9wB585INbL8O/hVPnPkSZj+bxm8lIRkNcXBn8GA2AVn1
35SJ3forgKZX2DbA5yi6BMePRtsrrXGg0Xv0GdLibuJXsZ2KWKNaEyf9UCduHTc8
zDt5t74qChy+6A+mP6suNAptpzNAvW8fL0RioNxmC57Is8An5E1y1JjnNYWZmBTp
SfHLcmV2oZa/+pSyPDrXk6JVYqBRF9gbBuo16bWT89GyZ+Nzd+9VIIQW39Jg+rVq
oMJtoqAOyMrmzr0RamQaNnqyZRDbTUkO+8A5rcWCXFVv/oTJn78vBnb3zpcb5+1s
8sDjrfTrJKKkuBHlTlPO3zqLvFryNQ+8CcQFudZne973jdR1BSwhDkU+RpzYwFo5
vfAVe5+44lAHYv94S0xBjKruXqw6G4v9slIdmCWNcq7WSD1UWlnJ4HIP6hv54+8C
3oOTmz+VoKUxhfaHKTOlE2pERQdobBQb7z2nMDqo59Id2UEsROcv45Fj7bRXlvGZ
0xmg+7M6htHfVEEMTrnRJnRMfjd6k6eL3LLI5yIc9/mcmwGn0TBrnAvrivOIbZwq
FknHiOT/ws/HKKnRH1dhqHRwVmbIKE7YthxDnUjCIosGZMicE8iqQ+V5ueEyL2p7
dhdMtD396eFkXmm/U9QP/5asBtfjYrqb97QJ+5LSSJuttL24shjSPJ/hTmHjCxXF
/cfyOdnQ+VQEKpKSYguSULRgtHuFMNsbbS9EhIGzm+8dWxodJ4Y0ycSEwFZhWjYf
YojC5mHTM6L6eLr2Sp7gTBTfeEL9xUzLl/VR2HQ+4mcjBWejJYeNiyOFOE1v3LHa
DmfUDqKy612qigQNLJkO6qSygu03MyFm1F3+SVnGAocWNhMsOHRh4E2qB57QjNq3
eyMJcw4pyhnsBQVH+l7ipKsMOBBTmO5O+A34Equty+3PnVNGzFZvPQKzMYolr8wQ
dXrOfAym7yC+DxcKqIDLmXC++3ttyNHzsbdLoQn6Jjfl0uvdU0jZ8gsOunoEAVoX
UxY2eL0mKIZQiM4eU/ySLYu9GJz2Y3Jvf6Iq7uX39Dl4xoIhu/BSw3iip3mcwe0w
9wP5ycGVjMAN4i63VGDNdQEgIoexXLWQ2Wh2f2GNPpaquFlIlIzZGmpJSnjao1yJ
/uqhfRdXH86Ut5IZGTE8WLnSQjDhEPax0QQgR7mc+b77Uohd3Do86KrKQyaBfnk7
EH/mdtTot5MBQfnqlDRzE3FaOnfnGV0n1l4Ta560/DftvFfW0b6AKW+VnzDRyfPy
d1ayWOo1QbTyepoEQ0kcYbOgHqB/GAyEyAgXGIDO/gu9CNR4Y77gvnFikna7E7Id
knHCEXnyxCV/h+VQUWfl+vXUhSWoPOqZYjLlsnGfrgHD5TYYFom/PGpGatI8BX2J
OX3FVCcRHwoE7HKQ02i802MqGaN921A9XNWa+PqKIyu/pW5Hybml8wCTC7VAkrph
eIQ2lMVEtSRAaCMtAwx9g+Gx1obSblkHd3wliq7tCiFwxjMun4RtNOJyXWCIhUit
KoXqM+EUIrWFGferExTOT2t+0iyAR73JkiEZ+oyLHum22giL5dyO231XhdbzRcpS
z2FMNRMp104S98fYgQ32HaAFrti9NDoHNHIsXOsvaiKYOe6OAl/Q+lFeq2Tji32s
PVQ6O/WMl3cgwLpuDEIvqRpMzqB7eO4o5KPeTC5Co6i1981eGquH2Yubf3sk4dzm
CdUcodV4eFJFV8aLcHuhkPcEGENDtMfwT5Z47SgF2uHu2NGVyvPaKs+j0GbzhGY6
7qNQz7mxVlNa6ILXsqkP3wxxfjscfbRUskhVanTXTy68XzrvAj7h0fD56K2D1JmI
CV+U5xLq0Tbdk8acplhGqwCtYAdW1ULNJ2Ky3G7ucsTNsQZvqMMWsgmuNSRwHnRJ
McWp/6i+Tr3lvGvUo5fVqM8De2I49r8nkZ8Do0vKe2FvODMKDpHjaEArPgjbOw9s
qiAByi2rAcGYZyHQgWXexH/7+TAt/4+RyXPR7+Q44yliNbl8X0s+UyhRlv+9hYyX
TKCaQDu2pIL4vNgMSu1Nkp5LnXiWPm+Pn9yPD9d7/9cj7VWb9cthiL/raGTUeoxq
kh8AKtmU+9Knzn5SNiInyeckoizEs57lDmHlK4vLsNOhDMvPdRmSq/MELZXWHZBo
7b/OnBKVJT7Gh06mzpHrhaZKnyBPmXII2vD1e5aGA8JGsTTImGkSRzhnziDpUnMW
nFOsE90Q7Y9+xVOjm31UB+vQ8OlXTq7D1WYGYxh4UQ4W8zr0QEI7iJAP6OdBt3ER
vNeZJQOFHI9yIGxCWeqEno7P1mYERoCt9p0qJofI3YypAqg1FQFFI5OCKuOqLTE1
Qdk69+1ZQKv0DrW3TuX4moyOCLeqUnOoe0s3AL1CbIYFKAq7VxOU9buqSH/U5LUS
yG/Js2fjejUu0GOvKOeGcpiX8Hm/0E/95VH+sGszHy7cWO72RU6n21PUtZyd1dUV
EW1vvDkvTfudBMNjT/4FBmaPOZ6eUFgffxklX98E4kRgG+Bkn2tmG5Ogojzeq+Fp
SlT5rAHcN3FXIKoTRNuuHksw6CPqFmLas4MnenmPn9erovDAl27yS0LKRMLYyQ+X
IOZGR/x/lL3GsXV2Y4kcTsFaQaP41FiphQO81qaYuAC5f/wYzGd5WnDfyk8JzoOJ
OyW42TOU1b2nAECq9xuLu3hIGgBg0ImWG4dNWZFBjtlLDsvvAfiWGO2lejoBE5Ws
ai5LGowcbqS0tsolIdJ0KqLZ23/kM6C5RTLDoEMSUsZYmfQr7uceHgheVcUSKXhl
oyJ1ImvLArkcYxrRwkvpV1gHOlUJ2IuiwkttfHyw+HkhirYT0u46ks8AKNptOMDx
AvBlBF3sLR1OJFYDnUFoolwn7nb4D4UNAHk645B7D1z9AlM+APDVINY3xiMmV6As
+DtHuD7dZ6uwZKhTDFR6vXPfZMN2QwVrUQj2lcfN9AGBQlKfnRwq8adRVdZ6m51i
tGpW1Ftyq745TvJ6FaUo60SKHlBwW3sj7aF4QZfC6c94nX92DGGP51js2CbHZ2ID
Q80ZahcRr1lKysjLyx8e6mR+oBcRxNEIy80b8zchs7m57SA0U+NgVOn06AOzz2gW
oXFCg/U1CDMO2Kb1ar5kVnQ/bNOWSF6hV7nJkdgC8x27mcjoal9KFkvLbAz+8K6S
mRB/MZRKHJ9msOJG5MZJKBBFcEKWEQ9/Yk6S6MWQPfGuFNR+862O+0p5tjvVepCX
lx3qJ+WZ9kPLfxozYyNA07RGvg2GR6XW+IJd/6h7z1ip5sVsUJj79MXX8NKlzsSD
XayM7+7KIxRB9xl+SYIqH1BfXjfdTZGS416KNLeDeDYLY5jP92+29H6ib2aRxkot
cP1JKBLEXc0aggz7KDcsnCuWArY5CvjsL4u7ExpCzxTrCkVr0IjpSUyL10/GNPkw
SPY57dq5yZzHo8WlQ2OeSbXtmheFRnk4gEeStokM8mtprSuyZwKve7bhcb91D4kD
S7NRqErsElr2yNwlr5/mQEhgpLeaEavCg34M4d//lbQsEIAYsdRfJ4PyR5+eMu8p
9nYd9/rcwywp2TlRTENOo/LwptMxaemsSpdfz/KsRxeFFW0R1WBPcWcKIoh1mQXq
JBrtxlnqli4HFsHWP+iPE71oJG/vGTW8gPIyZ5szMGyFgQiyL4y+XoXoNb7c3CwU
TM97Q4DGJNaeaRKOlgNcOiX28SvMGhF6NVX2f3gxYwxogFw4j8frHcN1i884txYP
hw9ATdqtBpnUkushbMvij4HFxrHXEw7NOCiYllhiMfQWVLgJ1LYUeJS7l9UkJrHx
GZ/NYhGWG3aCRkI4dlnpmq/knlACLPdpSsrC6MpvKQ+31jo8mkDwRkDPjEPerE6j
CcYsnXVKtCYNnSu82mHRAZQXPDjJCVvz3M0r7zfRtkcHEXyr8v0MW2G9KlUs2gbD
y0pl+8DASKbCJL0LMWAdxBRs9WPpLLk9l19y4Lcpr79ZqMQWwoyZaigRXcKiN4CY
aqRnr808BiLMUXXh3h7xZihX5tYFZo4msaPnf1JyGxBmw6Ol02CrN+/RnIp1fIrA
bll+lnmM8mlZnHLyTX8asfqfHUV2VsX9yi7HAfB6549D1HH9lPOqg2UTHQcLXm/z
LuxxstQ/8DihtGuDtdTMbd7ItuF3xNCM5oaNjQ/Ait3BTKtNnS1dgMkMiyEgxGlF
auZzk7k94+bx0h8vN6ThscXxgQfwzEN4H8KKWZY+MIIJS9xcMxswGLRHwPOahqpb
zeDxC8Q8ka+pe3jpGEA1DGic7xDkJ5JOMND7csEl6u2UwAnkTTkCVypA6fcwOy2b
IdslanBLQIIz6/CJUSAq9rIOo/cS9fxVDKzmYlfuEhB8LGZ51UO1Nmfd57Va2TJO
LAWINBOqGJrNak6f8y5Elrhu3RreDuouaOycYUxpylQ78Gyl/FHyfw7GRVsaguDo
EztzCW1Wjf9dsyfFuk+TwgyIX16Bf3KYMv6NtjqEQDCE1oWCBgUcPmyhx8+8G2hK
9LvYDSILaSbqqAPQvNZsr5C4CMAAw+zNjEQvUxWaugO9og5ed3i7THca4xX+A6Y8
Pi5RBx4HjZT/F3yiTmsIWYdG5HVQ58eoV+f+vqoQUtDxnIibEvQx5jDRITuGV96s
EkhtOfmSE7L2DpaNrJkIg/WdZ00uyCjfntBIzOv/TjYlAtdMYs9lviPQ4kSfHHrS
UIVE2uaUrnW1I1txAJlOGpbFkzfzWmEFZuAq9P3s7XkB0W4OmQKF5PrU4+yxJKAv
DExG7dbwJZ4T/rLBbLFxe2cp7GSGft4FECtShzZGnhxb/PpsVu3EQFTfEMo+bvXG
vFktpLt541/BSFVAg4/e0UNfYQ9KVhEa+N/PgnWst/FzON5VdM3c4mPcq4hNQGrm
UnWluOgpQ9p3Gl9wzyjBSwFg9UDQDkC0Zv6yaEM8LpicvS82y+UqmWQIy7PdobDd
ddyhJvqZUHyqXw1p2gAqzxrpyoo0W114NV6rIbY5RlxGezPitFRHKlev86k8hk8S
q9HZ9kQCpxaOlQIQAzw9ZqomhyU42fzHCZFYt04coiIIj8rWxeRUUrfxiqjG/V53
OlW9IHSI8FvZxKLZEcldQF+mV1przL+0CWLhcNtw1N90ZjfrAKAoj6E2pDAf5nS6
wEkz0VwoJq9+plYIhYbhTQwHjMnSPcDOmgf5B19PhLI9JVvneokOJTw4NEgSqVav
N24LdtXd97je2WKFq7JU+ByL+a9Lqfyy5gybqznMKTT9KbNctkVJTvyqVBJRxTol
U+jSD4+OWqIdWyqO7YikHMF/3b02StxxWNe+8ENB2CdR8xdtwZGrDpsTMWZWB4KJ
Ycs4VU1xTn7agomafdZPQv2r7qIumlySlWAjTZVZEgkx2vB6PFilObiGytaEAVZK
wj8ElMILtcZXxSAl7+Vkl46KOxV87FTIMnMIr5+4vi2QJn1irLKSvWt4wA+hXmcQ
cDP8PRydmLRNuscwjGt9QCNRCyGEYC0ASq0toEuK5vjqIdoyhT50+tpENv7M2EjM
aP4mwxZaP+3fUcIHXCgtsK6vEXOjmSMhvPdQ1Hl7/S8lBrFVoampmp5iDnTruEup
CZ34FWJTCZBan+9mH0+wv5wdWw17E1LjQD2y6FR8vvClesf2UdMYioEPnwfvQU5H
XRbW2EYV0te5J3CSi2A9TcpW2XzULcHOqDgb8Yyk+K7sZ8topd5RyF0ii0d0AK1F
I3BUWQoEqCMXiOIYp8Thhhm54XR37mVZvTb5ELkhElyoPyHDWF/ROfgLFZDSxRJh
NdM734cirW4DXSX/+UGGvd0fb2pZi4fIXhCHdAuZRPNSRxaPQfdJMs4G8/3Wrk5N
aHWWloG46kJW9k0IQjgMvdVvWISK+w6+QxfJE82zRIC/G/H5z17u9kAkcg1Jqq8d
Tyfri4qC2Fns2fEHOhrJNqrMMhzQTX1aWH3zS9qEP924sl3gCNHCahh7RMKS6NTS
+VZI0Doc2OZqhj7/+72hPHW+63K33BwsAAWjB/qhN2/ydSJJ9R3mUqb044ujUYdB
zyFM3BFXRfWEihUy7uuGK+NocoRpO1tv5upMoLwk5EphplhN1BLtJKRi7yjwddMG
rfP3AdneqwhF+RFrswb93vxUZYunztDkYmXanxTHC3W8qpbp/veYG7hAe974POhB
oO8A5D/P73B6iGRsQE2VkD3XmX574Vd2czrtxP2+1PQE1xiVWQyd3alB7GEypjrK
vu/ilCsC/xGPDeH3fiYbWG3I8bnViQAgzhZjP28P8kGSoxMd4hiseUptfeDCmhEd
Iu5/qn8IkpRr2rWsbFJCAb6ozdOL4gchcYUHiZQNBVL1LcnThMEkaDP9RF0LWOlR
0b2hfr0B7ewUTC7ZswPVXnIB+Oqud0mfkCzWjzTaXAfKJxuABrjJncentUZ3hjoD
buAJuoMVip2MiM98RQD814OvWNcJCNoyhEXdu6K4yPbN9py4YSZ1HW042DCLo926
7kNpA4kJy4pKxkjWcfpkCPNJ4faqu6xLRXLxXZnajHwa5W75b0fMHnUP3s3sQ/M3
5R6qOqQ3pr79Q09sD5QwiCHB6Bijj65EyFrxdjeexFZP8CPvseD/Yh8m/OjGE/LA
Sn54UUgdDwjcXaT1hgTy2eVumDmHMfAD1BTz3rf4XNPpsBu8R6T29/joY5HsOTkr
l+aAIykH7ULKYSPTOYGnfS6ITkB/NjECnNx4WpODsqOmyd0BiFvecyjc129H6GXS
OVs4WEKFbKMyVc0md6fUtiHgKv7dbk10BzW2SzsTuJ6kP1IFMhkA1+U4f2+SdkCS
YlN5kKJOBc8kcnJy2rplrU1JgYuQ/fd2Bb8LZbaeZ3GcZo/Sggb2q0WH/3a+EKGD
vbkokMt3texLetWeXeGRiVn0j+rHxeiADmOw4Pch2iRf7L2/Xu8ODNjfKXddCgrV
pAOaSAM3/KAyvYhgRgtPg0n9zDs16bdYjVRbUKhOEBt5+Nyn3znrgSi/MtuYPPMV
RDNQ7AlFxY4KvHsaZgQ8+nhBtPIwGNK+ppU/ApP+M9qLrmNfQK8JVaz4FQFY8uJe
dLJJbFmdme+G12rGdjAmqEPB9IqS6ozMXnAtobx5hfyxyeozgSv5wVgmlsosa6fz
qRuTInGYSfYShnG7WaX9SzalNCLYIM7R6iQiuu8Jk2+QBD+8f3Ew35Kg/M/9keDD
9SB2gxtR6X5zEmupIviAI6m2crqMiMMvoBoBaI4r2A63ozxDUueDRJk7Dv2dkD/r
/1TNwbg6/YEpVQWROTn6bWwqAhwjHO4Qyovxetok5k2Vn866QqDccB6WrJL7uono
XR9enHEBZRRljR5wW0nZ5l9RyHOEK/n3R3GzaWOJMaAtWBJWguEYCpDTX7+vzni1
NAOGaM2uM38rVk6PaXc4S8NN/rkZQOGTe6pZAfoOKdQQMPYCqfRXDEzymPKZiPYQ
w3KsGzlvehKAfr5GvfosCaB8TaTNNdwfdkd/9TwPOSv4YgvPg7TLZRn8kUTXB9pr
y5ZDePC28fOk/PZ0n4IUVh7j1DyDmfQPEy/0RFHSwZNlmmIoosueE+i40CcNTCC/
te4CflTRspnB1BELYNLsONOUZ0CULDVNPoW0upSiCsXEyLB6J5sjJRrsyKC5Ljs5
UlkgiFVCS9iXwSlJSO/4uQ5lqEYQTzvE81MEGRD8PlkxyjkwsdR6IGJiuj2QqVTn
mPuR+G9XS60I8u/rN101/DWKKU6C0TCNfIjQObdbQTv61zlooGtEsG6cF0SvlUyT
F8Aa7eRmzoMW6N9aOUKkAoj6vd1+QR3u1YAq17Bgf/1VPkd1gJ1QADY2+Y6RqMUs
y74P7UXUftCmH7ZqdkKfeSlj3CLm3j/6Ri/mWAqafowclZikrTG2XxTOAXuiS9P2
SHfpA7J99t7pEcSxda3BJPIw4SZyMENluKw9wj56WR6XsLuf7tf+O9nFbYkvxcQk
VKbuivmeuDYUQP2ZN9E/DAcYiT8hB7sIdw2o4mEGN4+72pw9VvXQCHnQe9G4atoT
9UkQDnK+2Zrf+1fqYu5zgRD2nr2b4Zt5n0ktmk//tE1ATTUsgI2QP7qIZfrj0JTd
c6lkXqOkyc4IfZpOQLZSuH+Ykah6hU6AMNQlD6/R8pu6H480+B1r99DRiXqaUcoA
KRF+4Ze+WB1f+IOhC7B48/I2y1MG0JmQ/3uPNf0iwM1KEzZHMm/0pKshG6Ht9a6B
SK2ziEfBxjwDHHT+f5KL0PZs3HX6Ovlay8H94qVPOR4fFv/5W/+7nI7OjgBToFoJ
YdvEi1GuzUmBjfkapuCMxfqLh8z8AEG5k0j5HQeNKRrWWcLtX2hOuWbTGQLDSqx8
PDTRTLTj3HFlSTSL41qdu+HURGsPE/bZeyTmCJd2hXUUThx3vWkVwR07oVoMEXDH
tgddYE9r6yP5IklYuqRJV0Otvg+UQsMFGYtHdCUkPH7F3f2vhA28TjQoIiqCXxgc
d8fLmTxvZuOV8fOWKVK9b2TREkIZq4I69vm+rWFTe06wNoLum2/FV/FKkB384krQ
uTcb7kHUjUYVy0BRN0u6fcq2BKnGdf2tUGnGnyiSiTddNWCu0Ha0begzolMxGeiG
EUUPsB5004Y+uNz0h/j9Xeb8+sC4z40pJub5/Ca/VIly7EUFRzsT5iIBempoayaT
o6+pH6aihFzDk3kQL4VfAACrcKdmQIMC31+znVToFatNHTvVZUjqRaCj8xc/TnqI
1365/NrnSaC0bQ4kqWSmA1t1Tj1Em3sMEbeimEgD0sNIUTpesLSPnAdAz+EIDFUA
1H/VDZwSA/upjq885gLLcjSae47+5RikXczfNFfDtC0mWGKGO/rM0emgcxwCSfKp
We6B5PezGHKtHxb50zpKeYfAI8+pwEWRDGlRQ32gxm97oNi+B95gWtPHJJL/L0Yz
lEPsAdpRvKE6fYgRlGxLz703SH87tEb3PC9CT7w9Xo5sxhrPNNoKjyO98IodkyZL
ZQigKVMjyaFHNUml2dBM+YMwSz7KRtcsK7mM6hUP3B9v1p/DRY3Hgvl1eMK6iexe
gQdrm+ToVgX9H6KNEq8LXoSf3ePYI8Nc4UEWiLdDnXThOsuzfxsAhVZYnGEwAN+s
7AU09UVOno9+mW5MlGSt29jV9Sm6J/MnTUwNd/AyppkZbaVet4iiOSAUnnYsCJ+d
d1Go92Mt0tYmIqeIeqs1gvmzzqL+g97AlkoXcYdEfmx8thQ9yslQCxnChg5nMg88
wyQj/QtgkfJJUVo1NFGSccmWUIVD9mljnFAyVzn3rlH5cUuCqWMdmdHeh2Y4lUm+
OmDbHqq0hZDXfhpmsjVuhqIKq5qjcMjdb7Bpdym9d68ab78J+9n36V8b9FmyfoGc
Itx7y9H4fXBDNcXzA/VHHm0y3SwGQg/2gqiXGCFeITnroqGQHkpckdt33kX8IVI9
V04fkHVMKAkR5QE/MT+iAOiTHncGwLfIgQwD+PqTJ6KW0aUqvkgyHbJnW8KyHEzV
MxglziwZdtXBbU5OiRoxlHl/ZL/XLLK71Mb7Mq+N8xToxz1nojR+FpysQjBDKwpG
jxGpTc4JLtOMbNOP224DzUmR3vJY50ihdu1KMuGkKJl1GIQlZOjzzSdSxTCnGuy3
SsX8bgwWt+FdbI4iKbJT3cOPzvEC957odceGfz7Y05PHQfFqv0lY45K0eJj9hGcl
7lG/yqP5NZ0gK6PCNXEhqfCVEfqJ5vT6sc5jgWc0IQDGCwZ36evCGlQ8dkfhvwOH
wEX6Ik/RjD8PNJku6eKeRHSn7zrL+BKg/ZUm/Xpimha/hpxt8Ij6tcZu8Si89VH1
z0yoncQgbo1SYf7zxx+WvYZC8a2jx83Mm7oCW2a2vkoziNsKqR5YRxfoT7h2Vc68
wCWvd8CD1k0vW+PATPUK7lOGVLntbzMxgyHSKM21WhGXsdpS9h2j8aUoTSBJ9FLn
X+XgKuzl+qW3kN/7t9TISXMuZ8rZ7WNoCuEq3OZR2PR1rWJeJxQNK+9ShVwluATK
I32iz/kdOfWgywlLNedIq3zluZ//Kob203APGccv7A07rEO+dwPTeFfVUpvVj3Sy
4sU6HkEDtPajjC+3M78rnRavpnFFTJgOcJOfOqefYqgpqX3QOCJ8ZLSb40Hs4/FE
UXV7QJS0TjnKjpZ8ixoAS6Z8y24zFfsRUwOBXJ7zSw2VG0d/vvT+WqRyOJPRRudA
+QA+2vjRjWOSDFos7fgxB4VxsVPRbixkLGIT8xlI5orRjjUfoHwUGmC/nwM4SYlI
K620cvchaCFqWouTEijv+lYr1JemKdEriOCRB44NbGInm7CGRlzdhy5pI1am7MWE
GoRIfx+AT5bA3k+6dcLrB/kQoBtegXdc2X6Qr7xIeXc1y2P+xv3k4/UM+wDFsSXs
NEDBCmN6NlUSkWh6YpNLyV5D0w6NMfM0xv0TMs8alc9mpXseqQq8J51LY2bjHsIl
YOkOHvUxQG8oanim2IlGddlHReMXR76ZWVNn291xmqwjL5EymIcoNtHIiZDY1jyT
AsTuvxbT8/hLIKOBzDpoiE1BqojBgGK1GNMEJoZJj2IOUOVj+BX0u++JpAMG/H8e
qSu1cKKWtE54mIzl+RFALlZ52Ma+urTvzQYjyQOUFywg5Q1sqU/ML1baLjrWOAiJ
hIDdPWuvtveVFLhU/0gpDsjq+NzdkyZnIZFzv6/ZNK/Oa6K93hzlGMQWqg0GDUlI
7pzNI1IWvHlF6gtVSBUtVjIOzd/kvl0CPHHydvx5fyTAoP7gT9Cw2GHyiFbdX3rR
3qjhGg1UpnzCIwdLhAF6HeCTIlU9Si+uBTYibjiBKWmC3Vt7ar3NNdMGOjDVPVWu
LAYBp5V4/huCom1eznfLqjZq0XDt1v37VPZZU7gTUBBmYfabHl9NjRWMxFPztH31
LrLzYDrJSH0BksWl7FF6kq3IEYiytrPucQnTSAnW660wOeSLwTiFlxzBifDhx3iy
/QF2v+oegLSgj5trG5znAMdsgEats+2CsZy5oFZBjwEbf0y+wWrXTFAlfaomtlV4
5eEYxeQ5tfggzEYaKasHTZXYnyKAEfxayH03Bqa9HZOUogPQbe/XsZ6dAClzW/HN
JP7bvsFXyz0rXWj80MKIIMpj3qGMZUsvnWgQyy20Zkd3Hy4Zen0wT9LlVXi+c6Pd
1JQM3C/r8veW4WrJTH0D/2P9EKK4u8FsFVOGNtiKsP6e4kPtO7i9tdPdO9CJtwfO
oBQmQqNvHbF34p7ZGaxUjglogi4iGpyGv91DDhip7o1y2FVr17iUSPGfarz4FiIH
dWL4rGGY1iTRYQrBXrRbSD2bjGizHJzOxlXFCGiw9fyM4mQOM7WLX2llXbV3uACg
335UXBWgBP74lrOmEtgOvl+Ve46AbyCOCQyvhMDKHL4oPhiFentQuY1vyYVgAn4Z
2hJBLh3ZSW2Dfanr99W3yRFlAW5m99EOkvZ3RWZgMwuAVFfidPihummjoM9dqEue
llH9U3lvTJL2XCfsqbm/wONROvUNJIPeJh3J0oEotV/9ASvtDs16e0c1LLlzsYpS
rx3ZjBq/aG2SO6EgzJo2jcWqgXtjRjCl1z/BaMvJVVsiv31MvswDEJKIwpVryW56
FmtuKJn1P/K87Fzie3Lu4IXvjLO5byzH++tgrxlOFgy9BBMZm3lviJc5rapjgicG
mKLNJUo9gxcW8ixKQ88n5nKoSgrNaO4rynexc+tXL8wYfP7PocFn8LK9/M29Ud+m
H22RYLGVWt3qOGLyfoQF+xYwuU8Rwq6rWWlXMgUsi804Qs+UPuIYgcxpRhBfC2w7
naHaAazn1EjVCWG2L0i4+rFS2L6FXpKY01YAnlzvIsJCBgGp7RD12GqRHcuiJany
7KEzV3ew9FAkSs+0xemZ68h6M1ufCD3inwzPS8BIiKJncHP7+jgnRaSoJyB0WiAj
JGKXWkyL3Q9j0ow1Fa5vYc1njiXtJocWKPMeDHUj0BRKAltAZQEhtuImAfSM5pB8
2075tMKHZV3xlDzIl96qIlVcvKvolbq6zhTABbz+6Hy/wqaFgrr7bp+8BTyqjjhU
7iYBL74pMU5KCg4NgVLEMUBaIzwKaezrtRormeshRDwXB1x0z+ktC3huitlkOBZK
qYV3VtQw+ymWdFlODTmfklIzMHpmVE34oatq14ggTHJzFGSAJ///V5FwpMKr2spP
aRsK5ovZqcwBJNa7eO8AAzADLnMZqwLNnJmJiUBZN9RdWIvzxXOMw+4BN+dfpSJc
LGMsRv0W01spVfD5LthgpXYV0CnH/Lmq7e/fW8Gs2+4YPIuFiV9bZcnidGLkrA6Z
UdoNRwR60Yi4xpx9MfSC1ZetV032lj9V6FnDvQi/lMA4kOWLqv4YEUIEkgEoCozp
AJNAxfr/sI8pquxF0CjNcHT4BTk4nuJKpnCsCT8m+uFOt57rEAOJZzWLQxo/vESj
vMpTXt8QHN0lRBlvllUhL3n7DRsbYerrj4hVe1c21/SKWDQmL3fGebWH4WAGFEHP
vSgHQcQCBzGYXZkSpkja9hIXs+SCeGwl9BoI/kK4BPev6R6IWrF6HCnYLyl8wkhJ
ED1p2NVm6a4MPn4rtvsd08/lGnNgaIztdOR4jCTeF/g/w4BVWU5L7+nr9AT9jGsH
w1hyXXSv7Y/5VehWKe4OCckkZmaDh7x0FC+/oIahIiZCx45Svdx5OQmecvU0tUUV
P5IZhobIS9B5I1eirMUgHisfqtVL2eJeDgnvevmkHtgv0DL7ura3thk0+wSpt6pk
2KK1eooCLWo2r7GZeC6jmQZRVF8huzbU+BcxRqXr63GvOLosgwgc5k8//lhlkLFE
NorfZf5D2LKCoMADLQI75OENW5fTRwYNCahBRDNzGiGR9vyKXOK4TfWdLIW1EKAp
cWcq/EsbB4fax/sTQOjiHmU//++XYx7Rljgz3NhkO+ozvxmXLCdOVvDF9NKCwssJ
FTbgeUZnPCIuwriNqc2fV0M7W4uUxNeIqPreP1vzf8w7nMFuo/5bwgMt8E4cJiH9
KXkM9J8NvHh1jas0igBSPLKrwMYVzn0xR3oTLHDgON858hUYdtynmlU2+U3e9+FX
PjeVbL45WJpzVIE2ljf7jGiDHzucol3StcgnJba9CQPdz6AOVXBRCn+YBvwMN+yk
zLfTE8u4/DCZVaREc2sJd8OgUbBoe3dWYlaJ/+/z4hoWiF0b2t4neykfRQOGv3Pr
y5d2NwFyAvc13L3lg2ZHu9PpzCmvnlWDpS5r6sSc70xfySzpIwxNlpYCoA4lNZYv
UvRKS/gst3wDT7T1eUT59CkI38At9rbVqnfSL8ieLKDuUi9VW5QdDqyb+JVwe7eI
mbYDTLr92Kd551B+lWTelutbAXke5HH8X7ArV2dpc0eBcD7c65sKa31y+f6BlE1F
1fFSc8XjHmWQ58++OrgU4fvHkq3dhmno7F+Lht84W3kpwLGyCzJE7pCmX93wURfR
GtD5bDEcKEntr2V6e9GSw+9nAawIh5Ne52/XOAhztNkXMfDGm1YipgxOFaKSpVtT
PqAbypvD9cAtbS5z0DPE/ylILBNwxhNHe+kgwkOVV5bvGhQ1H6BGFj7lbhoTUFBx
mP/CwtO5DkrM5xBM7Ug3gimT/tNGNQda8awbrK/DuNpw6NMHKdjiPTRPkf/9wGZt
DS7x8ctNrIeSZMUU/+uy5FqzNheFTaMc5Ek+9U+OXtIUHdWtQVKsvXxk/3EciBCB
uEHNN2q1Jxhy5upgLnrwnPjhdXXbRt0zl1DizyFXQqyoCEQkhUaazcDaTVcJGhQw
qUEppRm66uj8xfM9cwDNBxsbANSxfXhJ4dzMv35a8WIs9weUoKjiKWJlCZE2fUZU
i4ssTnisEbYD7+g3Z2krlUn0A/8KGYcZko/hdQptxBRZTXHCcIijtJXDLvpCLiAd
l8lu/Xq36p8VE2JeHrQ/bEaMML8qDdIbq41CcBpj5uV/b9M/pX608RXjfg3tge1h
r05TQrWkuUrECTTVij4iLCDApZNIjk8QplzpS8ettmi7Kklf7MAerH3eVokGrpDy
4HSfLWCO+ibmtWEXWYchZilGXxf9dtTRurXGvu9kK5z/HePBo2XMcvcwh246OnbH
QxyVuoCtWN4eZ3VvCyXbnY/wkdKHHn45iityL+rjkiDt/nP3Oj7polVVgnTxr9fq
blkRa2FpgvTW8s1T0uWUQm3Ws/ynkjVtInpASTBSbMIio8MqIr/OzUvgtmn6QV41
U3zMwyKNLucPHmkx49TCGLp4N2lMnsHlrgRWyVLf1qLIeAPVQJVxc3+2Koq+ojsE
/f4ZODW+NDxuiiCZ2YFmP9kIcpZLqoo8jsb1V/O7FqeifN+lv9zYnvHEED/rxlBa
/LfuXEE2//BJ1KXk8PJOtNzzr3Q7aXdc9gSson6Yv6In5l12NrnhhQChc3dd+Ldr
VvFGB9fd4QnVi7vyBOKiSZaY5MU3jqeu724e4HXcUE30YlpjQ/PJbx0TpkSrYkkc
7a5zRIn6wdKH3IFIcifXG3IiP0J72pTSMd/FXUp6sz4v3Y1wDErMbMcbCEGwqCsh
AZRJBMmTb4OMK7JqAPZZUlSjTveVPMYpsXWmj+KA9cPaH5RaoOi7XDJSBtxeKF2p
lTmjm9vyXSWtQdylEks5jFd9Nj9toQJAOfeXxvvvQQ/4tEQZBBYrLwS3vBEQYnWc
bDYsByOfoeZHsE27hcZp0pMgvlg+69i6J8K6f1Q5h5xsVfrpECs+GLRrpYm323n2
xTzbzi/yYIKvqjZiG4E0bzaq/CgbhUmOu2fDtGG1nVVFmB3bnLBRZdCPFgstEJzt
JYvlL62YIbd27HH9IBr15lRDqh/ZoCTTjtyTps7QUeLwboZF7Yqkh/sbU+ify0+M
IUSDwScWXAmAYQStxFIydsamK2vuVWuk033gMb652W4HC4zbCz4oqm3QXBHDB/hj
0pef3Oc8OG7XPk6DgpTbyv7SKuf/UA2wjjqveshnexFqT4aCZrNxRTVKZ5bc9QlT
Qq8rlF6ND4E1r67NvgzrmGbeK1n6STcEZexiUE43c4Qx5Iy3L+ywIDGVuQCjm26+
EFdI8WhNoumpJQvuxC5TEl73B+AqbgPIngaU6JWjNQ16ef2YQMLMaSdTtbhAbFUT
GH5jnDbSwL+CKLGgM8J/ZZhPzuVdXHIy7eklvUSJflIFvLcbxuIJuZmPtAuC7x1E
blangDwGB4uYl/7BNeJQkPxTCRxwZ7KX/4Bne9V0/3zZZ/CFTfx8uvJiqehU2Nd8
vFYo+W2/D97CZvQVRP2ccIcWPk6tjkEerjzykG3c3ylvsE8SG+kXDtpyWr0Jyh9E
jvtLXmzTb9LCOgAn4G4cNpQZ4wrbp6RKzxyawGVeRquGqc8Ei99cdBb4DewDZukw
/tWgbYPLFJEwkzw/CZyr5BN+B8uCZJB51P8/94PyWY1pzas1XWRwiE0qvCkcxGKS
QwdRwykzfYRknclCGzKvOLKx5TsBfCWwfwAIbJ3aQJ0BjHrhLf9TIZogB7GsEsBX
eGS04Cqt50Z2n9Y0U4VtPR+xUI//jviR+UjsRbGBB4SKrzLinkuMbrIPAsdcjQrl
JA4NupTlWXf3Je6NoFhbocWJCJ+oxmVU9NCVm7dlhaRcgmNelZETV4U4U57UHD1g
a0+174ao43XFDjysIHw27xmSLgaBVZl7UwYQJAa43Habj1/feO9YA2ZskhFvqPhO
ImgOaqdoEofwuIxpYMB+c/jmkY1r4EoMEndk/E5T7hw077Wh7jqPOa3I3sb6FiDc
GYnX5y7TGAe9vNUsfPOYQpF2bMZz7bAAcoLDvrR4AesT9jv9hb93vOcIVwuZbo53
8VKaoyxvHD2Zlp0fLXOu2ccPeLQ8P4TA8yL+FBFK3OVn/JH4Aqi7bEnfvy2CSizK
hKeV64NGc4pWY7e53moftE/3pjof93/czQpX/7CDXgsTwH9Ox8FGqLOhAF8Ki7nM
WRxRR3lEhYwnLHxf4Kmn5ZpyWLcRdX0yPi29caVOb6G8te/pFK8BxQ5q16tGO2z4
5QTCY1pcHd3126TfefoO9qcv1/wOqczYnQ30HGUI93PwzDZv+zbItFmRFFE1TK9X
PMcV2jZFZoOO9+7ooG4TDO6nR/RZY/Bg5bmXwMoW2JmyqkaH5l1We9aeE6Bvl1hy
bDp0YrxS6tPAr+hkLFSkjCDNIv/FrlzPFHZXkt+7yTSNV5WRzNMtWmZhcDf/gR4W
U+av9wLvPn9OjWWBXUxgNbk336/wkrNqNuxv2PYZPoZEEjHhF2HHJeHgCM9J6/mg
Yy3qqnpWNmkj1sX3veM2PsO7+FLYrQJGanOaVExBo55wkAemLY0ykMIbokLsrqji
aP7mHWV4dYTSTFyg4UARg1flcxa+zw535Rq9oP+IZFAmLjv0Wuu23pbXaYXz6L9G
scEq6qRpPrJ/PAwZL+Tro/miRf/RmimTg3n12uPRSrBWRsfBxbGiPzfZwhLhXzIT
KtH/88GHR5GuV9pF8SItAIsi2/sadtN3/nBm0BD/dNoANOdIZcBjXGfTMimggJ6x
kVYT7+umb2HgA3mg5z2Djv7df96He5UTEpSuUozhJv0D18sxPmADA+lBqdzWM14h
lEIYfUyWuTlJuMBqxiAXQmHarrGe07ibzju0ReFroJLrIhc6csBFpaJS4whVKrU+
v0eLJKG8yf7CLFEywi6WkTrPkubdBzyEnk/a9rbYROsE3oE1fhaAyVB0jiLnPGzY
9KrnXxszaUNuyT5OmB7/7T5llxEwU++oh7P3M8xEMEGYYzZjzSrfaOPKjB3rqUiT
bNIIsr7gDgB9mNW1WmMvmzIsabKtFiJRi5vp+r+FIZY+S7NijQp+TBhcrBxAVAZR
aaOQJKhR7YOeWfhbHFNy5swVAzTULsOrL3sHEXkYqn3+GADxrGRUuwW3SmBIHeHd
cqs5HUgGyipP873+nyv3oi+PM/3ZkH32LEbsPeyyB4ljfc7+nHtXVsBfbKp+ZISz
7yDdCYJQZDPAFBF7fWwSjQzOWwUCwDiTy7aCJI3z0jJpN4pZbCnYF+7t5hIzFXne
kzi34ZTxYKwg61a0Z9haYZqYhg5qDYbhPriWhZURXlcdxRNAuqZcHjz3ofcRP3nX
le9LIQf/zJSLleOcd2KYH7qQDOgItKaYFHJc7o9OmgRojzyXPvE2GKa9/HOswG2U
aMQa0ryE5JS1aHpjMyuRav3kdc7ctNRT7NzqoUISg/1BCxUNCrkrXhZMkRMELtQJ
2bgwa+ucA382GgPEAKiuRibN6fsK5i1VOa9ltq1N9tNM5qC4bGQp+eObs+G6snCZ
VX3sxMAn1Ppck8KbqstFlZ7IeBkR58r5qYy6Tbhma8M+3dCjyEzm5YHYZ7TumGqH
MvW+1iuSnWUnfUjnnG7krKlayDjORdN2mZm8PFwuB0u4gU8zsqLo3db+CWcGz22k
1lfPCNneu2jqaWQu+ImutAjKl6aRQD3VYp2VbN929xvfSTNsni/xU+8EfAANKJCT
gWIo2ic51q52vLKPA7ERWPkaFdxOTQ4tKqKk8M9c6y8aZqFuxT/YeUERWAj0tgef
FpRlyVjR2GNUKjyt7dFXzy0s6qbLgMOZ0NKpo2nem8IJy+hn2TMsz2BC2Tczhj3V
MlpWQjKe7j8UGzRFJn2OGoQ6Yxw+rruIE2PysXSQHXK5ZQ332F2bzdBcRz++8XP/
rehvf3JdFQsAf+aL/N2WN4vchDgfEqobGkMnHCV31ebjFid2trRRzF9lo4aW9Deg
vtqVDSmMm3MA/rX/RMc2b/eNWYle6lwA1Q5SXQDNGuuhhOv3XvAfcIgTB/+4rhcg
oUmzN26SHLNddkZnC9oZlzUAEJJJbjKAfzz+/zoHu3TE9vZ2mFxN2c0scpifSZpr
kK/xU69U4bMur5PNfuJDMZ74ATPscF5t4EkEghlnJ477Qps3zj8+qJX0YR9w5Z1u
Ct2quaN6rfdlNLr5eLk1NXL2TgemeEcQpqIYXdnNUJ1NxksTi2S2hiUgHCW/vo48
HbssOiIp5cM3xrvYnTlVCfBTcdhrxfgE0bHgBdLy81lLIP/vfBbTUi5R6KC4F9G0
YeGYzG1LlaZWS6G+02KNguaZZMFBGA43CWcqEYQrbPaW60weDyzZMz2UZ/1+hF93
q+zi7+X/31XeB6UtYmJA/jYfla2cD05z39X6TtVX/wSt+0UqYRoONm+a2eOjBtCu
s/rMUbZ/lcofJ/ifKjgm4e8uGojRJwqn/c0BvTPIUJE1NdqWUyL6/nFsltfQNdLk
nzi4a5z9Ve4u2Kr28d4M/c3XmYoc6llsSTneuuqcPJw2seEif/j85xOB37HOEhZf
HlCorLre4vasPVw85/XLqm5Me2+ouF9SvqsEUgvqr6p5I9clDjY9sGNyCSw3Kw3X
exzPWdl3Zr3UsBraN1sgHEEQFZyDc/3Ens1s8EgFrxvp+kjGK8pEVi3bqkcrt+9c
33zU9gfay42m1I5S3rrm/vjjthXp+cSKqdxava6UTyPYLofLLjWmMjuTgFZcp+Kw
gRv9U296oYqRZCpiZD+XCa5QXzGOrn0WdMaFanbKyB96msU0TApEan1TQOsGTp3s
q5vG6HgvS2cIiBIphQqkSvuhyYWqwgf3fCp2upHWLXOOGe8jvmyP7LQh0FJVC3I8
ebjayRgF/Bs3Gt9V48fgyRyE6KW+peGnkTpKnPxnDsuDrvDF96vIX4eh2l8BpYN2
1z1yX+6oWotVDO4mYJ2NlNiS1dE5J++nXY/2tHVnYRjNFCS54ixlzyoibKUuHPZc
lr9zvugb4xu9pR6ICufOTQ9/irxHoxFI5exzc1kcj6PezvYfWVlklAZ/C/aPrnfW
VN7RsSQHwPdGOdWfi7vOudq6AaaDc8sYknXS7w3BAJysLU3lYF/i2yZ70DCVI3aB
1S/DLiJ9Raa58lP9CqPszv+VMrrwuGzvhctlpSaij5gNuGz5giukVWdB42Xeg9Zs
XEIBX8mU0271L4vkNIHc9cz2O6PBX6okLLN1I1l7UwQsjbXhpHXZOhuXomDi76Df
hCwwMucDJXyKCqHbnRofE2ZuSNDsbIg1lcesa77AIReDu1usbnyyKgmnXtL+092p
8M5P52FzBz0Pa4L38WSkELLvxOZn6TB3oBAly2fsAeyRah72IUjSPOjKM0lB6Xgi
MCtMhhgNJLs5q9J5AKjMp+wa5dO1XyhMApafSL46zoMO/2L2NtmMT2nv+NmFOfSZ
WpwESkDDFZEPItw+1GDCY2w7jP+BHPQQApEt0omgFS6pP4OQAAMx15ZA9D/IFj+d
uL0sfMHatlHqT7nbJhG2itkRJa5W2dOn3om6c11gtNxJMJpBVidxa84IFENxEcFu
NnHlE8U0yVvGNLEkHXEjKSC66hW2C0X0tB/twuDjuubVDJJTd9T8/I70xIccE86A
fzycRBjnHd0ELcbK1i86wwXdv/WKzinrW+AESFyaLq9i6ZITawWVflNWqoiMzczq
sq9/CIsWwci/lFDomvL9Q4HwMH8osz2f8dSBSK1Rlin+E5lDo5tlTl/YQsa8S6FZ
HinZMu2WxqZe1zvLGhxzHwasIi5kW+inyPNozIHUAMmYBAjFhV0UfILlDgx1Osgp
BYI+2K97UXKIQKeFzoDsXrjG3TNxfSHz5iD2507B7Y3mypo8u0NjCsb2MWwJikh7
JK5tI8piFzOMYrmjxJp7jsXEoZLfWS/GOXmKiEQugXYwaGqv182PHxkFsTcW3oJS
aOJFVFiE3Ai4KBq7H4mDP/RcHb90vz5o6Tcw8w+RpXsmjnc6EKIFkify7rpuzFIL
UTYAOtFfy7nJEvZa4qcB8zIsVvRuQs3UaXjKEn5bs9ydgj5mUsuFHYIFL9AsR8Eq
dX8rXiO7RcGAfcEzG8GprmG+sZKw4xM8oXn/riT8pxLGcPbjWYY/U7OPAEwszZ5i
3zZ6L41bpM6v43nX6pPj0FunY2E4icHzzDOVEhh+CYRjr0BUwYLNeT5MDIFunWVg
nSsq/KBelo3ZjTj6HA7Fyr4unHcVhwU+UrX/W/UQ1XGDLcpbTgcavgHWvhbLmbfC
InwbDsE053WdBITcjh3jSt73RjvjRmztESQ+26FQBStHo0Dv0IZAj5QFs/4viGS2
pyMXYHvd8R6cq7Vk7lLtc0q91nczHkugOaD1DslngvCNi8nXRpPyuj8H9M8DE5OJ
m6fK5tHW0FJwiYIJKZ1ZgUAVWKMz0ZrpRMWDu21HTdRQDufkG55B3SYBj2fyYmxV
DgN4eEQ+rmQEuNsW/Q2LbMGY3QpQOTI3nbtoFFSvcLYWsIWJ6MbkvqNyU2dgRV5K
8rpgt92JKLchGCzCtxCv/6+RZ/13nDLtm4H71RieiNDlBh+ZxbbfG1qY/otTINq5
s24FKZodWpk1GKx1BUAvOl615Od7c28pij7m8sm5LlyE2V38xvgpjodmc3qL2Z+A
Rpgz9qjHKA7Qt1FlZDOLSJ9hFMgrGWq8gmIYLBwUCsnH3Mw7mXVmoga3u9Bx/6HB
EZov/wLK/ZzL2dP6+j8ylVU6ouGliFXMGDOm0kfzV39pzqqAguAZ21BZRDoYrn/0
V6lq6U+21YyjowhLwzsMmpEiW6tUPq1G0/nOpz/9K2zCSFtaVJvIhQNECUrlROl5
S82dS/0t7uQaZygYdMtaZrBQwiFobzTiyg1jxTwjhugBupHvNFrlgkeQhso27ioi
+DzmQz+cLNy2pWq6LMtWkNRaM8xFWPBNVd1LFyWlIQ1rWPqj0l+AtdFMwlQs51zC
tojLFRi2qatT9tb2NhDufrRV/e+Kj9i/cy347qkpTHReon1Am9vz4fExtP+zrC6v
JLjeyi9XZOu1gFkZLevvtSX/zpxlFNeXLQaKD38JCvSL+MRPQwdc4gm4m58W9GEr
0hew8ZVKgSol7qHfpFSXhHn5taXt/b1O6/+hReAPlVCcaeCxQkt4xWBtZpz79sjm
7RhHYupw8H4/A2F7Eh/+Uoh4EZmQ3/CwZkxvFVgihyPSQyEZqbXFE5PAoRKgwf+C
mmxIbvuS/zWPv+Un3FPkrdhl2c+Ty9+JnnStMQ4Cj1n4m2gD78DI3l1DQ2kP2yYY
cZ3UMKb8dQsy1AcyyC+UW5oBgc9hZeF4pO6rWZyNljChmlZiGKGpbLXa9EAO4sfa
O52/6wFbXPizWRZN1rX54zgWF6Dzmatyxh2R7pqIu47H/Qsnhar0TuGfsf1S20Zf
9Y6Y/8d5Eoo3fS/uiwv6hcC0DSt0shpliItyLxxHfTjm01sV7rBCtXKzACaguz2J
5n5IsxwEh4CYiGgXcRoU9BJyZbsmlc+TfRctMaVfC0PHevVIHWWXjVZ02FgFxmcz
AXKjmgw8o/0zWYoQU0XGpld90gZfm8le9v5R4QS42EvEwulJxLkAx5AjzliEdJeD
H4apKHauDWZHAsQcRC4/uU28eNAMVwqvLbBVONk0wzmG2y/qx1cbbtFaGXMBVC2b
KAJpknIcX5dWrfUp0ix08DQO/PjZI5olCKZjRLsZPcsZOXxQrIS04h2Aeip/cG3f
KMIbtIcWdmXR4d166NQPldikR0rgm1KVNGLJ7wXQneluRkPttO7+AiuRvDwOQfWZ
q05Ckzcwz7G1VJUbp6wZy/2HjJY8/Sy/14ALKevhCQgVo0so9ccmaSJX/MvMQoBu
Ld06azxlc+6b77IhDUgweicAvn5LfY2u+6EoG9v4cfWpZbfGzAJMSTDJGyemi2Am
mV6Efqx819fiKFR9l0EOoLtYxU27ceRYr607T9W/Ya9GSaYm7eyDKalOzRvVTKFI
oNKo+dYEJfySN3pMzOpvsv2oYMnwGU6DQmBBfYy4dfTe5P7cTxUljGUzCp6+Q0Gi
kDOxCqJ3SsLWq5hLTyYHKI3cn3RNV9lCybvM7TGRnaORr0UAgc/50xNDcFE93jHC
WKoZspddTfLPmlK/AMMzjz3laDNF5fULFjMzy4xpr1VZ1p4SxjrwsCmOxGlmNiRt
hMWJNXGWDyPfZt+t57GN5HK+pcWdXmKaJxrq4r33sbxJGVJjVP2kkvgsKHE/8Crv
RwHOisilFDzeZntZW92iXE+4VXhPfLvIe5ZSDLqbuDp8L4xakdjpKST3MWC354pw
dSip+6xSMyiiYwTKCBSFuPdmnwG1+iW7G7sCPUmkjhsVpq6ZfRf1zbJ78CNJ6/TI
RM89OX2U/sfKw+LORc4C6QWxNM9TJNCb55jH/zYEngFoalaG4HA0zymrOhKjsaT6
J12ZClunREtshrpkBQBmOI41QVpJc3ONMXJkdKvoSIY3j5C6vV2KdBPjQMkiE5Pk
CILL6x9msCr089sMEUzt8Lr4vlJVg/LjhTsN9KKuULd3FJ1r1UdfJxV3paprYxip
YwhWj43akUSnDavu1vrhM284cY6vAshaxHQkRS8zIJpGStYVET94zt0iMm4c2LI/
KRL1QGCwrQkf5ukBWm8mfKDfhCt1Pg4+RNgsFq86DZ2TPsCqxmj50peJvpP5ZDD5
Vgu7t1XPY1yCD/uIyd8HYN5I3A1I/V+6H1/TLEIURxcOHMcOcmOvi0XUnl7/PvOy
3kNS3F5hZ3AwxVzOAmfLKjHCDqgDFrlcdXgJB6UCEcrOC3H881PQbT1qIJmkrUoG
taOoastaRx6dYqLXi3bjWR1AspbFAa4KDKLIXAd3ffv6jnM99KW8ORi1OLfO+c0Q
5IAgyy5nDeaQNwkzPhMCNaT352uFdX5mHxfX2yfp6GFgtc+oNgdW0QXgQ1AeTFhk
fQ20XaQdOLLS4dLnBWb0ZUocoY8Fqxm/3HNUbZdzWkzd4KCCvXW+wQGynNFduPUS
NlW0obTSHN0aaYLuUtl3W90fR28oMCQOkRYbJjpKwqlPh9hzU9VY4CrjlkdBsSj0
bKf+Rdeh/IOuhLdkChz74U+hC+qdTXUPxLpDGn+reafiWnWLUpRDAHNgVIPk/kd0
s7s91y2leYCPQgYfQzWp/ZbZZMQG+xSRrDpmXpsa+wcaoOW/aYmXaXMcyRZaPh8z
UdMH85dIl72fXLZS0Baj3jIjXav4XDo+mn4FWdUZXKppJvluXkcqoyT9Q3AH2Vpa
Z1cYiS4v32Xl+CBY6m0E3K3BZznvnJnSOKu6d3+a1m4uAWlzRtjnjZPdf6xHoYL0
dfy1Bdhc+2CAxTWqTgtzN8uWgyekIuaS2KtgCP/okdrJF2D+LK1nUd9tLMbLoPWR
nDugQ36t7z0Gfmyt3G1DuqmAkN+Ru2Wiv1Q/P6Pgoms4wTtfcrdCL70JN3WjFq4o
nwThpWTmhaUTvbIP/aE+sieo5idDlHOdvt8ocFrKpxsviUtMoiT6cukpGgU6THMZ
cxvXbqsQ642Wf4vnIFav5ZanlswhndhuOCGBopMx216rKN1X+OhhFHPH7dR/lzt1
Ml0+ju2fu6ufSZih6kuVAG4XL7lbhNT50fC/X/LEVrYravsMp/pDJL+R9WghBl69
X/fLIUa0tG/ahLBk40BWCLIaQ4TPwtwrDle7p5Hmv8rPgJG0fze2tgKOZAWKaLtZ
cz3G4wEhiL1c4nwfm76I3UyggEe7EkUXF1qdqTugObw10xKdBSBhCHQ4jdnT0yGs
Gntbx4BHtahfnmq7zqF1dbo6VHnchJUdsqzQ+CXk54kqKGkEy1mYT7obSti0KRii
RYgU6910+sO2llVV89hesRgIDL84FfBBh/4oqzxfnLN9Wni9ufmMqU+MxowrZexz
17NttADWyZirn9eHRjDGwDPfEvec6f/ZPW5puBmBp2niObM1EKU+ykWKTfM/rmIT
yeDz0Jl5PdLyi+163uiq3KBTcUDu9Qj+ooq1sq6lxJyVIm7rCiWnI1r17siNVUd1
sp+Xb1z57/v5eNkpLeMFTM3Xme3iz7CWrGd9t0cr9YdzXoiCDe0msl96XaH1ApvU
9uT2ZY66lPkdoC4x+7LZQx1k8x5IDlKe1LRR+aYTdNJJyaJ2JJ/V1uNa7p0Qw8Lt
w8nCF+0vYAwvYtCdhS5xS4JncMeONWuCvkDzMnUKfAry13borMfOMc0BfYx16lRT
J1oc1jQSsIX1QOUSiGuAe+XNzfU03UGNzB/cWPBblnPkvFErRevecU5xMamQjA35
itxPfCxcCwIcAzuFU7fErgXC9h2LJnXyxbJQnsn4BKBxLZteYPxwsBNjjauM+0Cv
iCO7oWHYmSsAuXZ9fmjXFnXFdxRJrjKhubUjNkQVi23ZA+VY3aYO4vcB/zB4DGjG
a5J4E62vIOEJIb7pLhi/4R9oFW09r0HN5TT9SrMBlHvgc1vBg6YxLTQsb2tx0Qzo
wNcERiKObNip7VszkFDcgNYKUxK/X7UM+hFkYu3rWM5C9LNFLBGXVFjwO8NQggyc
8ZSz6SjIhq0A/gfXSHPnWJbYrcOOHqD6sgPqzaap8rH2SsijQ2IUf0EKcxIcDGay
BzVb//05kO2TIe4Ko+LSYg97LmEPUvFIPvaCg7qxa3O6+M3qTtCG5MM3PhtzVZ9E
PEbJzNVxbqBwYYKDwqPAMtMYhjGfZxNzFSsUwyAzYnVcxr8SUrdK+I4i1PorNQfx
Bhu1lxy60Cv/vlzJixJ8da4nUTKWJfYGn1eSLhZpJdwWiT9PBeCBfhL9bu/3YiEY
Aammb7WYgDeGaYKGo7wIBCErFIP7kZhCUBCfjQvP9sudlQaChAbSOQR27q3UNguj
P/qbt1UcoFFamwIeT2srZjfzq8/L3xktdAWId+E9SdbKb26hWwA96dPGaPUISP+V
9DHFnDsDAQRAXwa81kPrJp9VFjgjocQj2vU7Me8XFGOfuPOzUIoeUjhYUwQkhkJs
jocH6wErYPQj/no41MRqKbPgqHwsyM4wKlxXE1hE0H8An8UlQV+SdaHAQzDqfmNw
ohSd6cXT/tmp3e5MCTQ9y7sQS8HYnbt/ZiXgRnt+8ebdtT8NSQgjrTpxggM+S4+0
Z1PqTG+E+PxyS2iGv1fs2Y0MUkuPZu8chz2OC9iEak0D3WQ4zq/WBdjw1ZCt5HtX
yy+IMjfFct4CAVdCbDkVJtjsURqJEOJqXmM1eeBUoHhjdy5SQCMTGH4uLtcyKmdw
5cSc9lV/TFVqJWDypdXNjA0weLzJJqV1oie031DRvv7fFlabgNivrsy9h/GFg+nU
ifEYW3Kun4LAJB1LmhBmG//JtUQ94dAA/oFdnn0nUIixHqIOeRe026qml4eeoS0r
4AYpIplhC+j+TM4Z4jso6PWsskgZrm54le5aOnWn80716gb5n4KaSwwFYLtpTc/p
SxftbRwjSKLv7kIMckKT2CnCKYx9sDUCD+E1kd92xtNGkAh0eLT6drxiEyxEf2d/
gyAVppsYHG+1PzxJQXcZ8jH03O6/v3DUVKbsSOs7HnJbpLKNHgdw7T7qithYbJG+
Mb9pnjW5J7rLCyxJY3Dxdw2avhfLir+lGGPqEuh6AoDm9sNgQYQ7WH5RgwCL4GCn
3haXpR5OmUd89oNmrCfP9odPHQZ/b+9VlNi80pezrW12l8KC7fBfwp8uqr5BvMWd
b4k8o0yzL1BSOe8uCqjCgnN8+sA5BJ9qAwQS7V6aQBOr1iPhMs6Wrln5xjLXIQYK
LnPMyNXLwSXiyDGJM7D+nz/ntEva0KHlVHBUQRcdIxxsAYJYuqOCAyeZ5et929H7
4vVYYuXCyuEvlZ8yNlFb18FP5687DCmUdpvasQuIKXA0bVC0Uid8hRMCN00SFeYg
+dkgeQiUYUZZ8+A+vqdkNUuZdFL9zgAEzr6MVtpw02rFxHkUGdCQknpleBlepxpc
3C4QVTzdI2M0JIQoHnz1j2U298EEUg7O2twOBBYaNDBAtjaeXkFKCgcYoOLQbPnf
fnucxiYqQn7mXbtovLnSugNMGETuJw4HS5baY9DljckD3mv8lTkc06OPspDWcKyX
cxnCfVooQP1uUQvePTIAzxWOEtTkPAk0kSWbLDSh2M2woNYfsVOXGwLLS91dPGwU
mvH4DcyCTp58UfGU8+J8kzMdcTi4J09/ih3gUjyOkBeOUVSdmjQyTbqFoRBPPtAS
TLJaTGRzJGF5Bb4BkGDBb9kED7ZGWnYab4XHAU7DXlUrgKfTJq+F3uyzPVPQHFfL
5R5PRnJxx5+DcCSunuMLYRUT1aSxP8E8I5e/RVLDLdMiByirlkuosI64Vw4fqS2r
tD8vW0qtagsvFJ3p0epstshAhW092QBy6AFyiJ4Dir3zDFBZWlV1pEq7vhh6oE7m
eXG83/i+7nA6n63PCrdR7WJgRlVHvjFfJ6C3Et4xOYUNSO4m57iCexqHLNlAT51k
bkqdhI35dIEqjwne1vdOrNIdqjBwgQbKnrbjQmO9l17cWXK+9VQ5UyWMFE7ulz17
L4l+/rzv+XNOqHPTPdv0hoh7RcbQxE+Tjl5rZTxBoAVH7pnE1nYUQDwecYOD/jQ6
qTH3VrwGat1JlQX1N7gsXzDkvcCVRW+o3dCUe//ULJUQ0SrDu5K/YTk5blfe/J8f
cAW09+aSGlNi4+P3tBhp7bS311Cyisxuad5dx1TUMw2mgYbvBt2nstbq3gJBK54p
9e9kI76ikHH9sNgsh/hi7BgToYG5rHcKqEGPABabTW6bV6oUDdfXzPgKHczIiw36
ZkURymHdOPPihe6+2jXMseE9RwRYPHJdrEG1wiph27DGkaPPqVvO7WZgIm9tcdWo
FMyVDoGwh0E7aXTO3Jlajy2iXJ9nQ8iBhnCC6AGAdL9hjsAYWj8Q3crYpFdkqlKP
`protect END_PROTECTED
