`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cGbNNZPRSS9UxCenndZ6JfMFm43nnvHx7fGWR5wKz59aAmMAfv1r6Qlb3rC1GvYv
sGUyk4Rj0/PfJ6gQ+rKLFS1LME+uS7+6LuiK8YYe0d2n0jv1Gvl1i9JdNa8kA4Dt
gnyqL6U7pTWMFB7Wzw3/4//sMB1SLVMjUEF7dR+68tgi3ygTq4sTyGJx7IT1mcAn
eHkEwb+azy7BWnzhQjytJouiSL6enRfbLjrCHlAGmca6d8cYCjsBTY1TjUox/DuN
so7R+x8FogGW4maKCBwiQF7LOAYDUpzBJCJ66seSE80NTB8uzz3iyaTaZvaFvb7H
ehqAbB/i0cQSw1VeRPRwkeBfWdqdaVrlibqmf0q1QAG3nT9ot7bKoWqRGknOqPmA
5/uJ5sjg8ETte7t7IqnUi/zYPg2e8YAptWRpT0hY/XkUvTtLhWZuYXN0II9em5Hf
HPtuvbbpGgExBpra25Eil5cqkPCjUrEWB/M3hhplBxsh3+EeUnlzQfzggi3hw+el
GYIHW/M5RUKvnYF9I3c7Ty5PsE2SINgpcU05dkiv+g81tyxqZ67kD3xbfE/AkQlU
+3R/A9nb3950Q+QAiZAYjbdg6NAJistULAy4EdCtLQg=
`protect END_PROTECTED
