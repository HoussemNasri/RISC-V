`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pgu0TPISfK0deumuphqkiVY4IO8j5+fDZK8CLqYV3dwa5K3ccIPfDWR1a9JWLObb
hIpnYnRGOX2GW+POPFxt0JvNF3qBZNvGC6un7i2AJJREme1bWS8/kzGDEyLoazRP
zqnMxv0AFyE1IAQRbYYSlpaN5Go8V/cLK1Ka5+uh4IN15A6ZovVvkvuO/C0oIdad
aSM+iDf229ukshjKOpcnWG8gg36TrAcQwANiwvNs3sLTpMym9aWtqIjPmZ3KvogP
yvYVRwc0NtKFKMJQIyvkq1AvO+TDCSO5op5MsFj748g116xAt+3id50jVOAamiSg
4IdNkhAJQAxTTuxWZqbQM9gVbh2sKz9PKQemv82X8UdTw9GiXhnk0CDEQpZEzvDV
XcO7ZD7BoSPiXeEYgF/wDCAhUv5bq7IfzvmN4e876Ynkd6SH8UyuG2q3A300NlxF
qiJi42GyZ31MsKHakQGpiDr7ZE65c+IKNKwi3bLcVkjxd/YlZRtJTPEjaW/t7IgK
Nrl0A9Vt7OtPXLowus++BiAh80iP06MF9JGXy56WHO5ezAWfDbYLa2vE9m7i4u/e
+WiztImZWm7b3UiWTc/+BCXdFhZsObdQY2PLYgj2wVWTbCPv/eP12/A//0qBzDz6
R43o7990puu1ejPEAI3hzsTjNb58Qmsn5cNBhIuXzQtpx65pCaOMQINt4+0iqGp/
rsCg/AtAN6tPl3MVP1xTdOuby2T1MtzCtTRH+bN/2Fbth+RdQUPqWdtz7EXhzTnp
1zoRqD4b2aT3DJXHaSiuHzEVQ8ezl3+KTvDRJs8T2zdEVIxFNMwKyZSLThZd7Xvw
`protect END_PROTECTED
