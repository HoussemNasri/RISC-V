`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FUy2oEjNn01T1FYKe4b10Qse1qJnYGtm40NCTyKbo8vpleitmhzyCxdw1GlMWs2p
eB6I10tTEzuzuKlsN906xcK8o+4z6jFy9EjBrx5CkPwiYD/KmNZruiT24yHKVivT
se87d/tgNZep/hpGrY0nO3sXxku6TxOmeSlGDN+cht0WCzkf7mRo1kSRa0NXKnPK
C4/EErauEeGgHU/h7IFtndVtEeZoev4xs/dmB0Dk6gpy0buLZpujx4lMGVvtLULM
xPK89UzNvg27wbLbyvkx47HTsq4B1/oYBpau5/a8lrI9Xi66sGY1UiRMC5qhERGv
r2sLYpKxK5PAqzH3nLmoS/gjqY68AO6mm1aenf7iVYAzDUjBca87AnhxJkk5ZyxU
yo3MVlY4/VYpubvOq23/wxlz+5xAwtaQkjZxBiCfbLDDE0TJ2CVO+dI5ZUOHCUe9
9q/mPPJZ4bIw4Qwu0ZzWAlCLvVrnIe98m0GLlcNpoaBYJ//l1cJ4kSQttOY0eZbw
I+Jn4UIUQ5g+i0Y/7UoiDcxTPG3l/G1GfEJjA147u3k3r9GLwcwy8mROz5qj7AkW
f//eZs8C4njgCg7bw6QuMtRZvGjnDK8xAp6lqyvsyTPLu4loIHTUaZ0lfJeq6bll
DJZuPrLDsnavOHNAFKE+q0m6c45P+hsFf9GZqQiNt/4h5fBp0UIL0uigtLiWnLn/
nlMv/ZZClb1MaOOeqWfLaajXvmfsk4+vl35aNJKiFJEvQ7WW1CvbXLi/sQAApSDE
+ODToqmZEJPW8cNzgU0uYD1A4CIyY5d1sW3HMMAUfokr0qZKLd60/TvNUFUzD+vW
IbaDBfI0o22zqbIJAmDFV8xoYHNrhFwR2s4as+KT9S9agIZL+Bb6fOKpGAcX09gf
c5cACPjb67J8kIEV4gd+MouEiJWbyHGTEmrXGQ+nP9uJkcAiCkSRbwCwVzBX9gKT
aU4YGfTCuPgea3UagD7myhc/yoN5sFGiaLFNOJwyq5tK+rFFjW2jDS0/HqKNpciD
V0loJU2cHuVhWCCsA/pFmkigOxfZgEdbQLlB4jMy4WmQe05UJXDHGXFahIdIMUOR
bzdTIFuvcszdr35cGq7zjSwFK+Icz94dPwZjbeUG3OlRaorfHo7Quxm53x3bOZAF
5OCrqjxAFMMqo0wLa4kjS/0Vx/JssK3BjNVF6dGtJq9WVPGvKCfPusWmGBZzNqaB
Xst3HjaNXSMvgKe5CGRMdzn0wi8K4gF6w/P1W6SByEIOFUi9TNO2uCly450gDWjV
VbjHzOXX6xT9r/Zt5x1lEHEho5x89VEpjX0yI+z8a8NGh79o3OKQkan2QnodST7G
743EORSdOXod5UhG6Y4Cfjv8Vuk8+EVtnVPC8vtP8T14YzPkbiqTqHjZPvjxlOSw
CbDZMS2uInqn/NCaOxG563yk/dTxA0VY3v/EyzBIEVolT46o5I+Uu0R55WeV5FtU
GPpooyGOAnjRehOo5nxfNZWsRg2aX5VqKibQNXZP97/lH3WdFyFw5ToDB2vQRFDJ
5GaeYAzMrQQ/8L3hz9KB60Ad2CzGjrBhCTU08hvZUgZeeP2aTtWweJhMDju2ckc7
1S/pAcgYIR5FEHSN2EsFNkUDnl2bv/SfWh2a9hQJE68duFeJG9iSAOQBUIJ3ZQLs
ndDoDjMBrhTjbk73ULNWixQM9EBpaFVVhty336CynybmktoMp8Se1lAHL6hf+h1u
rod28i6tWVKGOX4TxrvRCxCDTciQXksnZyCN/qZkVwzQSHqZUCmKFKbJdm8TuPdj
qkDnhqqhFi5Z0ayugpd4Q2u+Qg2pagffwVJd4l7aZ//cyh0CSFgUPEDZzD2+J3ZC
pFuvd1oC2uDosPYmWnNbZunV9qA6XYm5L4B1bT29jdxnNmsmPATDjdaVWFkKn8J0
HYOmxf5U61aVwC4jxj87zrpawz8AMnb1YV2FPRPNnIdaeDXqJw/CC07b1J/sn9Uq
SDzMctpoaIZIEudOndUwOBFItTzrA9x+QTkBaRo1dEl0JzSK0xMb8YLUp8oLaKi2
HKr6f9MruZAhMmAlMtIBlwHAha/Nm86IUF5filnZ9DVDZIcb+utPtSlKvFCHhWv1
ijWryWneng2lLkJpFv75oKzUu/aV5C6ZUqTzJRINi3RdDm/0G8+6dW5H3vwAgc9U
MnwJx9GgtC0TvvUH7R3ODmTvV58mDkzgoSlQIWlQEgtFi1Pym6lY9DVpUrMW9OMd
p0GjmajkPFyUBXjomb5U8BldiMzhGidKXZWC6zGrG6kFDsdRZ0leCqO80HtUQ60c
ivHKQiVG8162NO/qJic2zAWO5wvTqeTh5tbBKrvSTX7uHOxtCGXUYngz7sMoGcbX
bf4fDmEp29UY5/v8vwaYpSwfAdbTt8Ori/P4YXzIUqlRvJditqxbMEgoUuZ2OfB8
EbYQJT0A7x+i4CF7HGy8iUVkqBy2dNeKZc4uabumDdPXIpdU3cVrW0swYwC+2gVY
5NdkSzDknABo7Fq2q9dQ1qIzGL4uQ8UFX3uwWjEnTnqQfp9wb3/3YRoTl7b+NWuK
Fo9ZXcTCLt4+UvsqC45ONwhtE/oLwXbPow4M3CObghaoz88TLNCwpjzuSrSLSxEJ
P2H/qQNIhukR2W4rFhYDNAgW/BsIU5hxsyK7D+Cpmk+U1l1FhueEJR6hT+gk6cHC
hRf/0mcjstC6py2oMgfu5VkMzg0w2O2oSJY3DYyq3ZLjF3JxacPkQi/18kyxEpDB
fLfSJrYqKYknFYGfoDxzm0G7bMA3EgMTDLDh5XDF1UB6jM1FmQr0bpaxGT8+nNMx
nbABNGVOjaGYzZfEgK2lPZtMduXhh9RCl4gyGwRVKVHAuu68QK0pSQwH+F7R2/Ri
hvttZo397RsiC7wnvJog7dmGYGpxenfJcHcxl7i99xe6X0PBM1vLLBT/w/w2jGF7
UsbD96p/KdJsFQf0akLEE2CYMeRNogTBBJsvwbP74ROSmPYVcjccEGOJis4Ec4d8
uCOzOMNWY+MWfhIWSVh7PTOgmT7Fpx9x69e8Gw2mUvL0845R3e6qrGpnN4XTLGCk
i210ylybrb1mgd5Y6gO+HoHDQ2MyN7OWl2WxISHG8oRVgrnBFZNu1AbASFwoJp6q
PGSZYeE7ejzYz98CcUhDvxYPkK2yc7mjSUcxFjJiCjN9EE0EemesEzu5jF67ZqJ7
E7x8PydLUz9kj9IbabG4Kp6JT1yqRQ+Ek5xh4LAx73ES2gxUOPAI/y1l9oBAltUW
XI61Nf+Sd0YSDbA640E338Tl4QzWZnkPekN0OJyGVOPCrBMTwMI7xBkjVf3ECEt2
rqhByEFouSTVxe69pmgDtec2aPiosfox5GQ0/qpdgMeKui8QpUELayXlyVJQM/N2
QeFArWjdIucTLHbWFWVaXIaSUiA20q8M/RNVpvAgagR6Ewk5G4mB5PsJWg+n8euv
MsFq8mfxZ3vU49d5Ma8TDelGMIc8v6d8O3MuInSgNsg5RGDhrhMzKTvwuUZE/dX8
3mJ8JCCVs/X/jbp03G6eFqsL04Imn8wpN1xkKHHsXLbLBLDvVwK/lPORZ+7/7tKq
kQUGg26nS3kSVMnWAKkfD0SyenNpWyNkuF1fCoxD1C6mVuQ0778DrDodAzk7Wp37
Dk7sRantPBnlYOtLP5FPon/tUrWYJOI/qjdKHnYDegx8haRVjAPGKaaO7i1bbFc/
owHuU9enk4XwYvi3833ycrc5oSATeUOSH1kpXUZQ3mpfxTs/5ZLilqJ8NagUzFdP
J3M7AwV44f0Ewb6HRIiGOcN9L2rK2Ur6028h4uC9mGyzt2IWfEZIjXT2qDTaN+1R
Zrf1NQb1MaRSVZakdZC/oEei7U2aQvUtaxbHlH2hsL0xPzCetPLSqf99KRXVSZpL
/HtXyqT2mZFCY+Lwy3i2s73qBScaGbPuFMXm4HWX1vLyEZvrkdZxLuAhffewAU3x
G/nqgjOCLlP4fp5sL1YKIs06nqUZwwOIdM3DD5o5ot1q5fIBISOy6wqZLc+JGU3z
QMlnNI+PQOCIENoHMoeeiSMkwNtb5zNZBW3jBdf0zwbGiKKEPMEUsw1jnpMHZih4
/Z6v23CR+WMSORJmUQyP1hMASCrjUj5iMii2U5jYRzOClfSRr28bPx7uf6+LP9RM
WJ2K3AinPRQhqwiHszHOZF9kDKTvO6u19AicZTYKw7BGP03BSBRM43QZdkeVPpqY
ukL49NAH82EjDymnXgkUHTsNG4eAB3n7kH1YTUcjrcYspXngg7Tw3t9CIjcVtYPV
jWHhz+opPESNUfXEg6VhpgHFy/nBXR+bdf+yb+ZO+iUrxjphlJLfkOsnfvJZgbSg
T3SSKtv2RbrLi5D2E/1ysNiKPV7hzuAXi/tahHTwXYk06nuiK+8oHR1gcMDeAWY/
dMyXYOuKVPghwngUlDUvyQSd5+70h7O0GUfdpPBrYgJgMajS4ZHudQJsstfjT81s
JAdM9/zuMVfPg4Zp0knv+CdE5pGooa2iKwrZ7AqlzNo2CJ8ukVvYAoKMDx3/prOe
fHP9+mh9SQbz5q17ypNDquEj5CvYmcFk3KD4twbeiuM7DWK1LQfNCkFL5AaHAjWV
A05KBmEs95vRb9vq2VDvesHF4669PMptj1WPaTveG4Y3qDaclcqSZ8EhBTNDm+ml
x4bmgio/hIPa/DwFJ8Hfe6X8WPeg1JsptVA7/8cak3RU50JGXrootp9mx6Ja+YB7
8/9B0gkzM2Te36kU9YNb00KUgoLnp9sDCfZeCFq7NNshJFFc/v4ZJ/URSQTdPS5L
qGv/9CfQOCDibfiH/9z+GqDSyC8LAMW4XqI9HwbVXYMFaq1x9BHHWrqoBeEI3Hsb
/YvNqQFvNhp9qG1stgsFejcnPnuGj+UqHZ9swrPFNJopJGatLXb7RaZdD3G8w8Kp
3Y2EBDJzD0QvAqAH21m6z1b1trpoRtnCwPL/++Pumw7jaQg8FFlv9vIH9srB2rnW
x3sTFEjlWzbGZQ7pfJt3EbwUrnSRpYVHlOVJ3ApyqGE9adKnk01TqJ4TOOFowGW+
31etivXuu1F6j1hNA/44yPbv4KrJj50L1lZptLoA0xTECkIOUUHzx0pjcJrB0iI7
EtJG92uEncsJc2PQ3YH/p/c25/dnAzuTHW7Vts42ncjrjbOpXxI+abwcbJnOSIDq
BCp/37zU8p27GOlEEVEZhlO8UhRQzu+oGiAwikrTMeA2FUuh5P314wxuHxjIUnO5
pgqyT/nR+T401UBRKzy9R4txHbwyHHmDdiPbln5lTFZnEjhWsISuh88K76OVyWpr
3f2/D4Caf6eSIypm5yiBVi7385SgFY6dYiIOYvEQW8CZgIXVsWhLOSi8Rn52PSP7
SBJjUzaEPIXBRaYMWRURSzzdzXkqsm/Yza2vyJ3cLPOA4UlLfFceZCLNpOieUtT1
8SKdUoFJtjd8wOXUiuKWgc7mc5Ijm79BK+dBFNWlih/5E9y2547iSG13J0Lkr4UU
xeUTcMkomuLC1cNi7JoaHbhaJI5RUaobIsDECP62eeM0GPiXgEQOmEJhAoJ09ET2
LX3R+Y0cGBsT1A7MVwYIDaVcYzNcMiWn/NqM4BZx1CglQNc1DhF+ta+bvXg7CBpI
6Jq61ilqKs1C04cS4QxpGJKJLlxEr3X4thozzUwIqbPtre7UvJGuAeQ7E2NJy838
Axr4MN3PwiiBcF6o+vP/v7AVogGKRTQfaV4gYRbnAgIUT/y2C0AwStu5bY0H9OXS
UDPmhBQaaVNed/wejxF9dAgQ5WFnxcEX5i97MoNWvSOtu6pgv8RXxBFoKilVL0Na
kD1knQLH7KYMc9ZN9Fyk9wqUAm+HM9mOEQ/v38XRZMdNZuM2zPoDybbxsjoi2MUl
QW/VbhBvqkevfjkI3HaTM+9XXxfNxWg5Pr4fDy5fAeg3PZASEONrc5ir0WoAPNza
63zjP6G2JqcvdU/nZTqHfJppUwbZk9RlApHR3JeYPcjfVbBLXZQVuYzk81DcSofr
WcnGRVebkSM1tTRZFCeGw7Z0wBwI3ek3DLO8NvU/aZBfEPhV1VFPFN/JRhoINujL
mppVcvovYsXKbE5A4aFVYJsXIhqpyBhilXCdSjTGOsCH/imujrTaCq13F97Nmk0q
bNJsr2iv80Ww/j4f5O8WUqj4KGpuqJTJE4e0t2eSLso2PVWqFey1fj4jLwjuobYp
fio6sRGl2RZ69cB/og5uAbE5zFgw5D6PR9hvBSIbxZhOe8nIxlPtyVZ0JLNP8CmG
eFMQt7GenCNkVJoaxD1omw6TWm807dQKnEqMoiVIrjgY2r1nN5UFNVXGEYEQgsqC
mJQCP8tvE22Gn8JPxt2YkwnwQ6vLiXM0ZIwULbV0eu7szp5PUwS3tH78bqU4ojoT
iYoXaEI2DEwiC/nY5ved1zbQDBxOZSH8wYyXnN3zcLKZMtMUqBn9Igl8u/B2N91x
fqTUMYBSYlNNK6LsueX6eWpqHgKSpfp6gYVWoEPFLQYBfsdp0qfWHl67/TqzIkxW
jAWgLWXNwSPaxk4PVrkABPG97gcldBEKvw99ZqwQLT5pH98P35InYZjFmyJ3crPn
JWnXX/7ehcWlT+CdPXKHkJahSjVwvF2yIqYcqEQGiRtKIIvrF6sgW1X4axVxQAid
BM1JAfOjB1PuDnpBlGniHf3xQIHEyEive+Q8uYehcGOdIweOt7q0JSopMypXjzog
WMTPw+A/OGMxKpJrncTVfuypV/8Tpe/54pA9/rlNfQm9F65tw9O8KEaLC0J4Fzst
L+J2OMTTVS0lWwf2IVe7vCSpXjSItlpUPRBQWXLsi4SPjcZOGO732sF3I7ryw6So
mRMCAv1WIaYYvyV92j6+cHbTbDFn0pv7viSUhl4sP0FzJBQ6gL6BbVfOEv/1G07Q
Dr9/W9olQ2Qiyv37uU18Tbdnpq4jsfY/NRAJUKPsx54TDYmlumbG4o3R2mg9HeRn
LeCRpEXEWT81y+dA65sFqgZOuLTxnO2UBdXR2a17QsQurlJxOwq6vEQKPoqSo/Nx
th1/Ko7r/ZQ+vE+C8x8JM2KcphGOf5pzfpnL8BRwkBZB6Co+/Vi9ZVtPYU4OqyLP
5iKQncmPrlIhWeGF1IMUvxxs56FwGeEECiufq9gvz7KotcIfEgkloFZCV/lNpLsn
K9Qil8tgm1l/lE+Sg62/w77SMcplmxuIxq9TgkBUJy/mJqTHBjE6blIlJIwIsPje
Ma/m4BfERHBK7mFo3vaU9ijC6EwequczOT5ypM0WjcGesyxEjISyuM7+Zkipqiaa
ZuKnxppBAcGOEed4oBwdGb27klkmE3+HaP2kddKhTzSfV2c8vrqEwVTO8eKSSaFA
DK/mD+tRqqhcpp38tW+zvPudeo7EJsysoStGywHuDUyL5JlViwyxOCcpJ+mt2O0a
t8swtwIGDLHbNq0r6xWBOVkuXhTyqTUEbWGxCan9xPb4qLiyJAVmYsGRY1VrzGsR
nwyvZowEaNWz0SWzgC1YxJM8XvZzVCJtKlwWhxkvMOCYAuu7HN6dnC8S0st9YNVu
jq7uVBntGfkPjgahh5vXZ1o/1g3swRUc4Fx9mo2urozhbHM5o/TkojXOA6ik96Sg
SG03Q0VqJVg357JeFUfPkpHK9Do0pTGIRleDdvKmnnBPu3VVa8/JuPvOTa+Vb4SG
Lxy0tb6lj+TOh+V7gSID9nbaZckwJLGMHfM8jsCKmCQgH/YjsxSIUMi9fWPJywj/
uaix45DxgnuqmFwxYyFsJwaSs4Nfk9nqaVbPPfjRPqR2cmNGvMGN81f8bL9VnvU9
p66Z4Cpz5FIzLyh0uDt6tZIOigDUsxJKUmiqCjGUSX/r4tRmczBzJkaevsiA9r9k
/LyJaj1eKycjMvSa+87qi6Q7z9+r8mJaJEejjOvNuY4N/3HlXYuPChILt8+Az7Lh
8lqEIyGwO5Q/xJxsEMVTtfZqHpqWeT0D0iqpkwZvY0Jvgb+FEokQHWh8Pfa5IF+y
QZFFqPreCOSlLCsqwnpIa51gwBAIZAU8Y6juQQkIqgoi/qwJ0eSbgLdbTqzC3z9p
Ztyc6Uh2Sjm1dgSfPvwIebzQwe3Uu+E0mSy533bor6jQBzT1sXiNe6fwW6Ttqnpn
3LJxKNeAYhLsZ+BVsVq8oNyrt4m1x2aOoXXWeAZcKQhE3+1TrRixbGUG5BIpY5we
HVyQbiMZ820WMK8Et4rlmLfjS3fsGv38PrjwxIBcRFpMGZhrq7qd0Ae88Xv+q3n1
wDobLzL6xSrFbN6Ux4+PSbeyHMmU6hU5W3DvOkWmfYYSm7bAzo67w1/6doJ79/8H
2SmcQlZq5kRxN1D9oyHZGn3fbiOmZJ9vvZcnSvCK+Vk4Rr82ZrVDaS2PZJ3IH1Kg
iB9Le8oBDGOmiNidgMzwcNSt3V9R92alx1Q742QfDsOLzvkpKxNJKLmhv7glFC2A
ZWAOvKmHP16fnifBQZExvT2yMXLLpr+vkhyhUf9X4wstfQNhQvjGSzv9E/4CYJhw
vmFIQINgPp/j/WvENVmYRxWCVEvDEmI8YMnwajnFxZTlfh1oIpxIJOOvy3DRdGni
rWRcaDlL479ETJjdZmmVHcdofE1Vn2iLtljCyuZEA8F++C5YhGb0xmsf7tLSKXAJ
7Uoj4aEgEH7ewXWReutbeSzGWlTcheydQDqSzNbK+tMWDbpj2WQiWxVQPQBRobpA
VY4a2/t4Ad9ydVgCs7XSnpUCmqpSS25fJ9+KAE1PMwc0cT1rPh39+CoblOqNfpHd
DtRKOwOeuHFerDfRuZJEl8JJhtH4jKa3Ay2y/xJLb2gt+bGXFdUV/eUtycmeyOYT
N5oFE6toBKlq2Qtt+xbpU/okyHRXuW5ELPBftMch5h/XqLlZpU541TIRav/A1Qw7
ioQ7SGealqM96t4YpIe4Ac7KJWGrCYa59pBTYQBKRQ+k9s8WDL0kS5lmbmJRWzme
jkGc7u8iyBjnuX4m352k40UY41Dhpmcx1txbrgHgFUfN907lQrzBJWE8xpVSQJYN
9ujVJAkKybvAb7K9u4Oc4RbVZ67tuoavBw2O9P/gr9URyx70eIl3WF5qOMYQHC6v
xA9J+MYSAd9CSWRyXd8LqUEg3rxGjrodECvSbKf6yAeB4hcF14erXhJaMDLirCQD
zlF/V2lNVv+jzf99V0SZUK+BbdcAJtXYeEVoQPGR8bVura6U6NiwH3xNWfCi94ov
x0QSrnXqDhWQ/Rcg7ErF2ZgEFEPT3BRmmNJCUoAcD2srFgvhftn/17tdXwv3V794
c8U5Ow9OZEapjV4XRuWJ1N7G/oxSQ/bgqY3GJi1elXiQio5Lu+Z88X4nEg4UnBPA
oueoGzqn2yxzzzC/Tl9sAjeyCMF+tIPGgx65A2Y7V9sJ4jFV94VS3EtWU9Dz20q5
rigFtdRItJ9IIVOUMBlvX8j1aep0L9LNCih7Yh1Q3nVPYx5fVSdyF6a2V1daiLmO
uYsOdrsJlmHCSQTJCfe1wmA6Os+msdzNBzpFVZIqUL5j08wqODpQ80Nq7By9A/zB
ayd1Um+OM7Gr4nBBz/du8RAUlxVtAFDkYFCu9dOTVl9COC2iiTqnij+QBl3iP1ay
Bnei9EDHbkoFTosqIPDhOxS+M5AcZin/o0HP6b6ag3R2QeXHfsk9LH0J2BfnwKAE
OpbZBBK7ski22aUZd5g5Huym6HRwn10agGURIaQykOBkubEQTqzwqtQBS15/gzvh
AHxUh0MVpRQTw4jXAJ50jlZVBZ8EIduyoW9dCGKXVR4mFaTcdu+vvU2jDHrHTlP9
K9LB22GEMRtvp3Ngjuepn1kJbgUPRdlWJiqIgGQZLyqGCOApVdwL1J4w3z8jfkQe
feWvj0I3cV+V3WxNqYFGBhZavVX3yZi3I7lgJ7aBwfOiAMV3V8lPmUbOydb2nW7t
GhUDD2erh8jP/gjvPs/L3XnnDhMav6UH+YqdlBkPRu5UFLSVpQgPRQilO4gxd1fW
acs/Nd7NZLXFs+vJsvajzLvzy/4rTvBxQ/gNtbSj4ngt1enCtWJMjyZVIW42vhhO
lYZzqwni3OCkfGsiiKNoT09kh595mTodYVmFtcvl2ZoFyQWlQz0tgq+qPRl0RDGN
1LxXgQmbntLfmLnKqOomiD8qUmO36Lj9ZzSwvkrNBpHWMQdngeET274vV2/KMHpX
f2opiX0dky46XH1K4L1/M/5JxYz2Vn4kIJLK2lBEsuQYBhhU7hIHEWGA/Q72Nz41
so6QXZNsT2WVSb07pN7e6oP1GiOTpaIRiYOvnEF8aqQ35JOBh4zRMwufi5NJi8G1
b3lOYa7VJVM+dDkeClfe/yyXKveyl7zcYYj3MTdJr/EiZ+Ej2Z/+SARdc6Ka0OPH
tQgUglZTo6Oh1oDFgu8ZLSyTikXO5Fm28oX29q9sXkBru8vBvJ98zbBvfoaHmi2G
jPAG+S/QwBVmsaFVtkWaHMFOGjtJWx6jPtL6SEIS2URU3p4IX2sBo2wMfmp98SiI
san5Ar1lT5MPlZf1kOEhc/xbN0D12sGke2QAhYgpVlVIcnhw7SLku+SpD0DtlXPN
1Y+bSBIAbTViS9EgggMKJZqdxhKgwTknKJABVKgGP9xqacy/zad2AdoFezckUs+g
NdO2m8kDV2ub7WiBYRIBDrcbSopO+hHw3RKncNPtLRnw4xNpe7qBAM5YPSKVufu/
Tc2Fs2T4a81bK6A5hbW0HGwzLrWsUMSvfD5R01QEfLhVSiDo2Ka01Iu7ajLtrhtI
tTyYwsIkiaj/xP7da+bYGMymOxHO99mPSCObSFkOnZ2vHP0E8dpZMKtHUZnpwyy3
AKew4PNkeMX1DwkeVY8M/fvPz6gA44AM2U8JGjvNhN7ZCacMbgVccX1VtJJYAv5b
PvMaqE88b8nX3dbpH4d2+TyPrQiXfJX3BKXFVDmQNaIJDq16wkGl2mnXDnvbrDOI
wEVoLTLXXAFy694Bk/f/c1iJo2JgiMNGgai/QzswbiE81rh/cFG/XfvRMBIoClXi
xMcLNazYA7Cn/wRIbSfIH+g0sGOMrePs5i+VYHsSbrWxPyCreJND1x91OyPGNVqD
V/8NOaXk62bxY7jmqxm8YuHl4igPdYmZ2kdmtfG/gBCwK1bhCe7VHSgAC6mpNXjG
XShMYMMdRdlfNcSkvmPj1/dBuDgilX0PP6ooXPBmMEBhz0Psb0ewrLHEI5WEXTlz
6jvjQKl1hS3OBmS3g4DaWtMrxFYf37dW/FDBLlLBJvwhm7fD9YgFXXzaeJaH+xht
jTgZw2t77XO3WQLElpEIRNbHb/SMcmqmFHgyuKeTktyq24hNVNSvWWSChzC/A8Ua
5vdHW2x3kpF8jSSqiXp6XTjNeIxbqIVNAH2+mPtZMuI4XGx+yfa7CzCK7nDzR1OR
JoWK57ccdohasqjyoP7Pib3kU1hMkYpt/dvPPspGSeKyIZnVIrMeF4Ews0b+ELDn
jmQUMHGR0LsTEAUPFLDKiOe9XIO07HL6hhkX0gNEJtKMSxgNqc7wI9YSE+Hw/rVY
JRbnI65inJt3cK1jC58zml0y2qp2PYmldcqc722lROvAFhFCJvlpukjylgJuILHv
np2grKM/IulK2TAFRnHpJdHtUQRnfR9ocslQ5OVfjb38FOtpV3xp+VPVOONlYxrg
PKufJ1HuEfCOjNGYqQV5jnqWAfOjMFQcGkHiF3A3DDCfHgDle3qSZ7mLNbIRiGOR
SLr3wLJ7CPG7oS99qP3XV/kG0Hg2/bXbIWizyiGLFXHkLpdqVuHOY/yEb2EjiSw4
aWrAVTflO4svdHqgftljd1yigKf+PjmXsNnJ8if0Z410X0nYHzcgx8+DbE93Mjct
18O3a+0j1BCmjCxQVcptuMd5wlLXagAqAJ+q/oKH/VLIH/wsmy2WFeUPCb81pZ2S
zYD4HoXSFabg7O3jr9JHK46fZKzBaN4RmDpuwJW0PqJPSlKOoY6dbcZR6+bQ/J5f
OXzGr6g4QFPzBdMmwbE158mSQrnVOnoQM3YwozSzAE+aJ8MHeIeELJkjvhfVHAht
rRqWZdT7qSp4pHn7SJJaCIYxa8MQ0z5ZCuAuFy/hER+Lnc7TGP+Wz7rnVRuw/t2M
4l++qULy1cc5PoS0IEPk2gu6lLRBGe8M+lYqgzDM1ZUpuLEjpkVwhTVcUGu71wqs
Ts+mT6IyXLerxiRAkQPeydqVWSgQGWWXnvvrIZgwL05K1qWeF1h2UYCfA1lsumjp
lNyP7uWHlmzXcJThfi+MA28tAEIZ4c42xmSU00bGdualK9ZCdQHm5dj7dY2ZOtgY
joyFtyC8RfOUN4zrJ9muS9XasjYZZmEV/XAXkNujBhJJTcU25hknpsufzLpRaZ5k
BFD8RlSzlchLzJZ79bHFW4LxrZGL4qftn9HQTu0wIiIzDQzu0dQUrLbuO9DV7lUN
dD/80YtOWf2eFfkCRaYAvoIfLzNNdnG9gLnZq9zRTMEWdNR6JkgNosw6tcE4NSI3
u2xHplGdoQirUajInMTQIs8wdUmF5yj10Zs7kQXkVjIy9Hz7xad6fiyp81e+icOH
Nh1EXhs8WO3ZiB5YBjlFGmKH9E1O+/JJlRN5B3CAul5RmnDTYhVu7IgEwQFrbwnt
VgyKevw6eq+mwSMwkypNJ93wfYR1fBlmCeHlTLJZmIXbe6JtaC5ganM2uU+4Rp/i
QMGxUEyZCcXZZeRVAHUjlnEexhxqyBZVYD4QcPPjBHVF9wT7HqSc8JmhFycL9q+z
OqUI3O9rfN1oW2hpfvgZ6q53bAwtbMuox42uJRUeRWwoIdUxAewunUBImx6sd9py
z5F53l7ZLhp5iEt3yJtid+FmUXA4FfbhIqTyfTZhLJUAh2AcO/Dv6jdp4ab9qMLi
JRczP8cssbZtmui/JnsJH0a8ImUiSHcgFJyH3423SK8KG/t3aWrVU3ike0SRcEnv
vVfNfKfDkD5pP12J8iLFDkLPCO95DqGdtk9+pbv1tKLHwErhRgjU1OYlEhqhlbrh
jaoRJ6V2tsvT+/c9p4HhWsA/319fcChYj+sLiq+Tupv6afNiQTawakq1zsVx+37K
O3WqLzJTRow/L5HFcxCQxWVeA9A7YC/6+ppreCnZGZwGiCHHUZsuL7wV++fLMYuv
WoeK2qNzPID04VhGpxa706q2bTM2Ow8UzhrGyVsjsBHaFdO3MZun8Pu6NXfposp5
iLdLZh4NJXfdCbQWkPcSUbyjSDXXaHGMkj0PnKnI4lL+UVmqH30YgzscAwGkl757
5MA/fmXZfr11dx4q7ZSIP/cdPmneOKoXo7btF1pdg47IM6XufWiug+1oCZDkdqZc
+R1QrGDxavBfSEL8k3Zcgg==
`protect END_PROTECTED
