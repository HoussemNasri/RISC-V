`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9TIs8c+gP5wMFAdNDSV9H3RMAtgPG2UYNA8pzRczUdY+tm9yWQZVBSdHBZwnf98U
IUi0qEeIlhHbhHd+MCqNHIwvUTTQlIk8ntpPXpFIdDHfZTud8JAag3BfN0l46UJ0
+J8qHTEKnLHJB+dT9Ga5pExeigQ8jjp7gbTwNmwjrhgYhbLxgeR3a5xKrmiS/TrG
J9Bfc5sB2wXd7xB/KkmSs5FzLSxBWir3viE7RN7YEVz+BnjPAegqieCJVrm9tOI1
1+m/52UU5ViMwc2OpfXSeCoOLCZevXaKpbS3TC0ALYQBxwj30uNUSCXMTuWaKMUd
9gBVtAJ2DTs7tWXlsaOwb7ZpnM5PbvDmaKN+F5wu/j5qwZJ12qmmqimfxnim/ANb
nvrbRssAn3sLuBmEBE76q/oj6Kwas81/vaIGBDK/F73MBjmuLZwWjH3L3X0Gu2aM
RnHvh+ce4l1IJ11X5by/aLwhcEI40dnQbZQ0hyAZViLskjc15G7YIneFXBoWJ6G1
s6dOXEKVcZ8CrDPPapZ46yuyLoRsb5bmIH9+bQAKLLt1j4CrH/YSNK5J+qdQR+J3
/JNIXm17SBVS5Znv92dHZB/whenHqWUilmsMHhM+RCqOiPohu3NXJH6Q/hVYBKz7
xhy10QqIXOwlEQXQ7LAVpkX5TfDO7ZkjkdBluRqhTXvKKIcNpsYkWGGsQmsG1M1H
+fgr717SrbTHES1MQ4lRaMeAgi1y3u7Vm5ShXYttK+WK6qX3bMC1Jx4AGwnsRDgc
ltLl7cSepghtcXHp80EeDSfiggeCZRdgT5qP2jMHJ4/NYkOGXqcEf5YeuaV1oAcu
6xe1ZBbH+IQtHoGRsSwP20gbT61F3IbSnfGNpXSa7+K1iubf+wmF4QvJ50OvSNkX
k35w2TN3rQdF2GznXlIn5SyDSbZj3JV7qqjRzIVJLxgUaW/MJSlWa6qs3kIoJmLF
5hV95SGrZdhJ988oGTFXdL965+qs4GQDCJfpL+445lJjp+WYj7ZeRtVxmKL3p5yk
9efvUEaC57+xjX466Sk8nLkGPUsAMs6uE5br7wXDjEbViCpOk2pXaE0RedASFYpI
YfeSzS5jBOhohcEtKMt/4Mi6VDL4xYt3g5EGjHK2Rgw4zVofSivpXlCpx8g69Ga6
0ANpSDuHAxv/5l4+feFlRUA/3zKFXz6NvSKPTvIdGO6rj8MOKRU1hXQbWFEKudgW
9BG5uc9RQnOfxJJ7Wpr1QNrPq4N4aTUAUnz/ZjOXaIHPsxoQ4QykR1+OfJfpWkNi
CDaTmeW0PLXHhnfiSdiQwfwYTHNsR9FsVINZakWLvNHbxDBCBSOcNWtwLRRC4+ln
bz7cJyT/zOIgMwkZp9OiUSpxrqBdu1/1hELfGGkjc9NKJGHmHxuPfJ/zN60YtWic
Bfw2VpnOFqHb7Z1tIu2KR3p8CBSZwCB0YdDMP+xrBI7gXWA8hGTGSFhTU+wUWpYI
OKAR6h3bFgOxN1y+zufGzkzspPgmZCdpWWSixEiEysPVbaf3DuwQ5SW1q8gZz7Ld
4Kyve2vS6b98869iASgINw==
`protect END_PROTECTED
