`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neNRPg3RIifBQ/cREB+Sy7ReyKAyUPoBJpu/vyxT00inFGkBGMl72J+NjmgFD6Pe
mTv+3tKq5Dt7iwyd8vAQy+UqXDDcH3LfoFHZS7Ye6ieZM6KaKPl+ZFpx7SWZTx+n
l35cU5K5ifVZQNbBH9a3B3JRgFezh29/c6X9YJRED6kiw9vzE7L8GxMmkOaDFtu+
zMJ1XYPa+AzAaJznTgrn8VrCCkeoBfhA1Tr0jd4IMKYNTljNnTPYnpGN6dDEqUsU
FLx4bvfkse+xBqX1jXvQyg29rlKPDafgDmMtYh2z+xbCUyrwnyLHfPxTjBMZ85qY
qDrI5PtjVVrAJ1pgMAlG96aw3IiJgVa7oNcxy3bItzzsZ6/36jtaxpv18RF9PCXo
luoxq6V41+wjxI1N8bNYsu77V7R3rwXb7kt5IazsI4FDUvRVzp9t3snbQbcwjUXm
iw2VK9fQIuonY85PKlToK8ocPnMQm9q49EJBS/z1EgEtFSYl8ie2YCBurjoGPLSM
3Tby7Ff+VwgaQZiqGEN2G+RRz2x23q3w0xVT5p9bXhSUnn7tTumrcMhpCuIO+x/n
HAmEz1RvCPP/SjpZdS7SQNw926q0vCiJgwvdv0u+4fpJij14JtCdtbCQbwh9LS+r
7MZf8mMrkCIzBknvFDptlKIOLYaC63DaXZexRV71V6hWr8FxZ7APV3wvvzPQzFvp
Ak2GZ3mHzrNNVRMaKbrVIsQQA6lk5glp/yu8QaHHhmM9xNuLzFk+JyjXk9hTzXun
V+VosELO4F/WsAt36l/lwkGF54ZqRGRXUBg0OL0T98x0ZwhWVM515a5mcFG8/z2b
1BcTa8oST8cfeKYLhmFibWAMxSBAx5HQP7VIEDdOaZxE1OBHyDOU3T3zk3KRDWgN
SvrEVxx9xm8fOq3DnsrJmYH+BSRiENtljRnLvVeVlTwm1/GtBxVFMhZaNpIqS97Y
ZHYtElQ36lCQFf6ulargtcmk8jdAMg13bOQUl8ejohklFefJuDIl7MOoH1jRom9k
/AmhyBTc5y1ubKX/BwKm1yu5Vu6nd0nB1nsAB4eoCSj0e6wUMyS3hKe7zrU8vURF
CpIgQzFRh4dMiymdnwKn8wn0NBnhvPLTJY8kuXGwzoZxUDabGS0cKwCy9NH9jIfu
gSMenYuv6k5uQt9WcltJKBKOyNXTSgj2it71wFchZVyXNUb0BBvpoYs4qhw8CoAB
16hQOYVZf0SrYaVtZ1NYJkQIMg5YHTPFAlwBeIrwkduiQQOSdNHFujTfzDc9+9Lb
w3DzfsMVrHhM41eP2n5CurnTxZe4k1LdXbDPkDMG6r61ueBWpifT2ruQLzLUa6yR
q/qeB4EW5T4HmpeKuT9pWoLyKyhEsjQ45lGTn8A0ylYNRtjHE/qkCbKw/e1nLRhM
UHzslo71iz+Z/V7Dpy01BY+Kyx8cmvZS9253F/nGrhWA6b8d8Iv0klR60q3fskLl
TTM+PLU2TtLIUMP4fjChOF2X4LR+7MWJEjfX1DJP5x/TnGrJG1GlSYaLSi74RVDr
d9hfF/+QNUSh4jvU877BLStHqHKo2SwjWfff1ibBJz4fE/TXyydDxQ0qTNl2fK96
gmuGB5C5ZJBzm0TcB1dcokJAS+hE6YnbfT0JIVVr9Mw5E5F4b1+o/m8Wkfp38pmv
gqylA0d0bLbFf9er/l2rjoeJznW58xtdUp/bxElILis58QPMlo9Lh8PV86yWor8E
Zg0mUw/Mnatr+ZxUWIdcW4Z8Fk6k30ohdSHr+6I6P1h0XHWTZEfcsHbeV6A5/Hcq
rIGbffk7nwugNaMJDqjBAYFsAU9nOZJqAUgaWYgQ6ctzWGIakPMHdDHIDy/H1ZPv
Jb/UyWbwkB8HIGLBlyVqzCDHvi8kqEa5WcMSgzGWm1rGecwfE0JfQ1bzWpb391l7
5BpczdW3P9s0qlZrikkFJA==
`protect END_PROTECTED
