`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+BPLl39S9AJcicOHe8s5mlOp6Zdxf8hHloKoJePXOSZqA1ffhQFXr9951+TWs23
Sn5MeeDlKgmwlD/ZW3T+p9SKe2ilDEUlcKO9LJWHUeE8DeCsySuVosfaDTdU8hxd
zwnVaF6kY1JvKokC/7FJd4rDrX7SFvDCM3sepMF3HqmWwX1ok89cB2GZ2X3fuCC5
ixyEgovYQakxbjqoiaNCdtqU9Lgb8Y94M6AVoNzYequOGctJZbjvhl3gGot9risq
kcvuFcRuylDw4hc99EmtkNGAhToncjRjLSVBZMXtHjerfMXLwiecA4wjNftwrJum
J0BHiIIQpmu+SEATeURTPjjdKZCkDUNm06vumqfgVLiNHHmpfHWMqKkgZlmRUna9
ab24TYRy5Y+zguQAPKs6fMpnIm9Y+B+8309e699c1vIAvqrihADZW9y4NwY8xV3u
VB1qxD2Pkon/ythS3LQOhTSJyP7CqNnznDAgGb8gGbnRHJsH7kndwUuNz3OqKY0J
rDQGPWjIKdEY450yBZCwlaO3PTgbllmwyZSehr7Ax9iIj/48W26LJiMkYEFEm1CI
cFjVH1q7dxQgX1aWWGa2AO1XsbrDnTV99d4NpWoUJNp2QJ2mJcqAlN8DTQLIE+Pd
jOl8vmdOTpaWMpgKBncodUqEBmfMkvd8XvHr2rA02IEyreIzx//V6jQImhAqHjci
EWrXYA3rIgLGnWhDdIN2s4NH2kIFhtLWRZBagMq8UseHU26+0nOKVdIgULX4sHCI
k6B9ySib4pz6/l+dmIoX4ffMKZNDkThQPYt2nODxTSOW/7eYkln8aTUN8/dL0QT/
liYibQ3huoJ8lQ7dPfkUGS37E4ezHM9X2eLgw2P32X5udG2dCfXDxvrwXvNvBMOm
XgYHTU+7IeMOhl1gAZx5HKirD19Orwqo+uOiOzgc3gF7As14/2BXZWt8zmLx3AV5
CwQmbAqPrJCaGU5ONHlC6X2pNkEfIxk8dYtjPAPrVp8cSvtmR0eCZ3If2OWbHh7L
+jIwniOb45uUTN5W7V4o1VJBFcIIMeLgqhKUzk9rwNKQtceVzs3+65XURwJwUgKc
3dezseoDw1g1PNUiRFuNuQiSo9DldpXiPsOxUalvpLktLC1PvSk7LKeOZlUA3jXW
xmciDUy7171zNfVyamIl1irajBJityzbQa6kNAxgdKSpGOvcS/YPZUX9Ty12vtRM
jjlMpGWfW3roUg4r4OagDUK0qffsQmp2h6Usp9p/hqMvmv7BN2hlsswB42084asJ
jZg+lgTCiKtAbrsjsiNiWX+d+O1pkNapuj/x5fcATlLpdM9qXS8N2RXEyFaZ1Sab
YA2f3okJa8E5BRs1UuM9wEuQTRbBt/woBIHNAUJlntozp2aMPPegrjEPl3JmRjY3
+4CQbwhc64m+I/OfunNpKx+MyiQgnNWvYzVJzsSrsRB5efSRjhj4tIDlql2Tk8Ey
vVELV9ZYpiRMH/qBcPmM2IzCjJubOaLQzbuVuv6oFYXQ7XjHVbID4svTSBYl3OoL
JWXCHqFSNQhUwRentvbB40mil0O8dtNRyrBf7q6cosZGzm2TnND7g3692lDS45JC
EbTD8MHW9OhpqeUt6NiKUGIM9vQCWyTcdweL2sUJd9SwjUYvIbSrp6tQAQ1N6Kn/
oC8qVkj4bHHpIarSBWiOQa5+eA1rEBjrVwGK3lAE5W8yX9gxN1K1wb6+zEgUwN0I
QJj9hLB9buPqRMjD4+/jCsdSk4V8iNxuAIPwqhNSMyKpFAWvzhA4ndv8ywi0Rw8Q
kDpJZ7HYMNyemtpF2Ase4axGMPlPsnv5Wesxlso9ROk82iSvULP04ex/kppZyYBH
7U5GHeglt9EzqbkL1zGmGVPmpbvBIbE7V110GSgN6wkXF4Cqa9ZA8iXJq2tADdIP
TScQpzOugsrG1angGuBWTTZZuWsn70jXX1qpdHsdCcnD35zeMxI9jpsDtSKZ12hF
x4izpoCU3jw03i0CG2iNmdlS7R8biYhIu5kru6zG5J39wKyvpxQKIxafYoSgqAcj
eB0c+WII73ptfM0Vne39xeIsxyCdWILAp8Z13olLvG8vzl+E+0uFwpCpA0NV0M6U
8oqB5E1w5SY7FKqlPoIy/6LdPbLvsiToDrVwE18md8WCsQxzDWyTmG6lBeDljRoR
IayqW4O3QVpiKQQn5lZ9Vm5m1od7lclFFhB59YoljVP/ZsGMr0bVsGYGt0kLp6WS
MG5gb2SLwZaH2PNFrDvEdkJR0F9x9BniyxuFOJlVkw2qfOmGJY30ESfv6aVAD0tS
yq/0keJLPpCN/nSLOjdjtLI3PzGRS8vZmr1+lGFvzw+N5Vu9feMwnKnlC0AGliyn
wqhH93nMIv1ZjLbakqUSexoj1BLhHb1RcMRC5789W4EKeZOgSYt/S6AFfMx+5xQv
dAy3yMLlnda3wsi+jmjGmu3hvzlq1djjy/QI70HGAcVlprqA6sBluKzH7lAScHF1
3LS8OazeCbNtSrMHnHG+0IuhgFDyMIk7Sm+1w8nWFBHhDnICkEPS+z5TYhEiky9F
hrqqDQSGRBMHpNgBVnrKcLgCkiawYJA0TGMDnJFLZJ4Y7O+7R3q+BtYH38dXfWx2
kiN7e33j9FyJgHf4euvUYrp58pxYm4ZCka0mWofalhNZ35tFixKPmu6HzimcqY1v
EyNrJ5Rxz0IDQSABjq9Oa9XtAa6bOZ9pfbrbUa1ib0kCQNtz/YwxfkjDHZWFtjjt
rnZygd7dsBfzqUFT71TffV5S1VfUKg4WbHtyuSpiGY3iOixZ5/rxsczF5aIHIPkg
Gw5G2KwlZJthLNa/RCZrrpywr8JzNgXbaERbN3i5KPFEh5sjAgCBRBT9zqWmINSS
fLG2FHEEr4N93whCyLmCMBLGRJEujdLTZiZEIOubGB8H/nb+9seMl9X/5o2KVMuK
uY6qcPY38sIMuVL4QZbz6GwC94ZR2KM7OHEzTYAPHT43jIHn4t74NU4KirZkSOTU
EqWD8LD0y4SSi59MkdheUR9RbE7YHy+QBuUAiq82VEzIFz3pQbg+eotU3LY83eD1
VZYYj3tekLIIRjTIZa8Sn8Bm+kmeFiutp0SMpZuwCg339E0UxtiNHT7YhMgnYzg5
E3rrMWn2C/bsG2wUWRfsAz/yZOqXrCn+h94BrXqku74EiS6KTLPDYal+RMrhgrem
jgNfSPfX+oW4sPtV3rv8hHuR1Rw+F+DABDwzv27r2KEczY2CKxO1h++L1HZNG8Mi
RHtTsB3Dh36+51GD3dlFhErQcbIjsH/9V/0m0CeB69pm7vlxTJj86XrGQvV9JINt
BvMYwQbf01nQkOxPcsEanAQh+jGJRyFzoGLgpIH+P643KXkDX7UTMw/StioXPUc5
Irtmh/3odkUgguVuIBtRB0uXPVMiDyY3xOsWheDN3yY+BzO0F6Dgvvt8q6rhg6B1
r6wTYuApjeOKQwWG8xeHGZs2TMryEFBHnDFk9/taFVyB0AYnfpf9P4VrT5AeKDJQ
XqID2nP5S/JX239USWMBMOZRgivLCjkXQBG2eCCM2z2My7Dh7eGraa81lMyEUj5C
JWmtHNNnLXLcdB+SAU+3F7wKKWilOTrLSS0ZQr/YccaXFKmCdpcUK15bhPLlFAzk
eJi5iZpLqCc11nD6EeSNWuB1+riPvg9vDdkJmkedyRMMVuKtvQf9Chixa4S1A9ck
OLe8zSMUt7rIgvWZaeU2AmY21tOkeWZQmw0UpgrR1Yki0wUu5V6FlQXws74tobl1
O83EAJDBZenqfQqOZ/dvN8ZOyf2MfShq13+DgLkRFMo+gZpAEpTSOoFzgZv8q/Ik
VDgqtlpd25d98V56yoGFiFy2/xHTGuASnSytmUc2F+HX70DMH5wXlKohycqropMO
AxRfLftcfHEC6+e5AZGd11tZm+MH8p+3Qvmeh5uPV3rubF4rPNbJI5XoM9uMf/k/
wOdKE7qNyoPQYQ6K4q6lNS9mpzDN80TXqV20dxue/b+u3K/9Qa2VeaZ4p7Elbok4
2IXp8mCFE+fkTPhPSotVhv5Qmut5/qQNmkz9yTsgVnUHKtx3QIj2NO/LNCLRQfW/
YsrlPgRuhrvqxruaOdK3rFZ0QH2PPNgDokpWS9M5zSc3plFD3FN6hiR9nA1siZvR
c7HeNVRTBDBTlUwVq1tS2xfplU93zhmQ3xi6ujTdX6IgyA8V9cjOyv4s822kJrfB
2j2Mnf2PFLDT0vB2qRguETp/XZohP6/gUqe/ZHLJvwgPh8kmkud9sm/SuIPUJdPt
b63ulJN+n1tVgZtK/I1pZlvcHdjYP0s5w2TcJPZDPNQ5NSOsRbCbYEwAk4CRZF96
YzW34xBjPDBzWqFXXlASD5SoZh68EQNOP6MO9YhyolS1lG9+9KDEAyO/uKOaqoIo
aZDKGbiMcUmTi6Fanc1bjCikn7ofcF+2GRgVMd2T5t18AUYGsvoFfLfZNayMANy0
2Og0hDK/UShbN7TUXCIndMFdWjOKaEmMEzP8rSj3PaE3vV9TIpLIYhH3tA3d6IzX
mnUfnfJb1nauv+nlWqmkSxYYWhi+17U9zd+s5UgJe4wuB5k6PoTpHB5idCI2Io3S
0orJbyGV3/rrDpERP9u5YRWqFrRYKgnUbhcoEoxmahgQRLYpCDxRbmXzI+XPXj7y
THUqiilkxvhux1YQifhrKgkUIF3rkKGRfgZOOGyE9Fu/r7okzS+Fsia3ZT/s05pw
BTWDtt/cBJgmcw8sOfkYPq+LUUSMVNWEVr6k9oCHB4jDNKcCgHAOKyvOhk0fY6/V
uN4CzwsxNJCvcFGv3qYs+6oAbJONA4vkQd60BfGnlCPtGKJFGDYgp/+D7TCLsDG2
2GwDiQbWda/pLn25EUFv1aY+exs7a/vg+A+kA3ry4iFKd0M2Xt1BQhslHXQVLBLv
/ivygvZ3LYi+nsL5mrL0cBxCR6+nEM1p6taUlddfeJrCrinJXgRBVb4G4NZgjKf9
Afh7WtyKph8LGko9JY5q/IJsz3hoI2iiH5I1xPjqTse4YvVKyFT4RSve1k1zipyh
N5btcxK8t6XUfFtGN7gg6TQ7+8MXOXNcGpZlEqlmsg818SvlrUO7S8pcCtrLav3q
RSknYek6ZWEzUZ9syuu8eBjK9qKp4wTp5TxiVyZi1VcNcmrR6gBPDRSaKBkwzULy
Ozj3fs4Me1mDRPpgRcSMk7WkIInIJDF/SXZhzl8NGyiDB+iJMf1oxhZWnMZF3ppt
hGQGjKy9jOnk1L0mKUjUDVd5IYXesivdJ2NKYdpworDw9DgNHQXnGQ/CS0f0jtJc
mbHPGUOUcxZeYiLUQXVJa9vS0Hpy9gK8zq3Wr8Jn5q8DHJoDU3NHrmZMaJrrol/3
S3i05/3eMeb36D1yfWv/SxfOAfvD+wbvDNQ+wfVvfiXRKEM0pBfiNnfm90ypRw7E
69W7sy71dXkoHXasTEESPn7dEvXF8/iYdrf1faQDS/FM8MNouNCEA5rThTsHOho7
1AQ16HkTS+sk/AvuIZP6VsGGEOJVNIyFT/RBLPPmFW1OdvE8hxhO77y/zKidPHa3
hVVz8LpzhIhwemQiYbZyVvzz+UwcMb67bNR4zew8FkDeAXV/29FLrLuANfArZ28Q
uEMO/GsqERtVhM3sv/fAxk6DJ8rNtvg39Day9ZcK576rLqFKkbeecRJK3QbxsALI
scrc5Nu/F8GqmTl8M7NEtGgPJzY+KhA5W8n+2hZIBdYOoFVOuCXNwp+0w+/6gewG
xHQSOcsXmHdpeHdAcCw0fPqc+7dmrf4N14DXdvHPnzdRgYV3uLeuJ+8+I2NRxZ+u
s+YE5AdfzJ4a/f4sxW3SIePsdgQJKplWVCzmRW2PZfkwhSClmE76/EfKo26L4Hsw
yUVUsD5AQXgL4EbuB4DGP4keoQVze3qAwbAqLaQWo4/1/n4ZBK3KS9tAvlXgiknN
8qta00D3M+bNEqXXvJjhi7plpHDsqCC7RULgcEcHdoyL+47G3VyrdymXCt2XCDtG
AXErQgad2QyiAWM3wB42v80+E8lC8Lbt+uJHEpxrm+tFxEM+dSE856NU2BT7LZ/b
V+XvawVBLu5TyGQYoN5xOzULZxJJ95ebmPbszefEkwOhU3eeiDC+JB9zRZjyVHQi
fNriaFAy9XXPlaaCyZc0+9yvW/8GdBv4USQOulP/Nf/zmVMEn715obSHlkKL9bqT
2X1+0l66Wr/ixvN4XTSklv5tRMekg8Ifz60TxYO9m2IAuTCmShx9m1yUqEWToJFz
3PVi3QLOzpLLqxKbS/ICfq65v1kPHNixcFztrdTNgNG8+pzVcbIgCuK4EHA+Rs+Z
HtL9ECMcYdLuboBEOD0k3T3sjPK5DdRd0N8OKMlbcher4YMpgToHQ0Pb39QNXqAx
Lq2LCdsD+/SRyujHiimNga95SMzupC8IYOV6PjFNu5JHtQ004mIyb163qtiEUZYD
w51poJW/rrpnkRWFR4Q4DuVgQBg6Q8RMtCqTJnv4WkfJ+r2jOq96OxVoVAy4LWpe
TVmsu6yIHwhB/iGxJx5pYQnBCPlQ5Hm/2EWdy/vwzFanh9cEn/ypQv2FKVOINZPX
O2kxFP+1TEGNRmYSb59xfNnquI48cvx223csNHthqDmpnOwkH4usIa+ed8zf5sJ2
Ex/rkYDhnt2jv3XjmbItoEBH7YjuwgeTVwZFOZgkEGHzcuB1L3F8S/lqDha4+Ndn
GDW8MDY4YMrxT1TQPuXnTIcL2df9EE4nZjomzNcmYvZ4OGkyoIo1ZJSZnR/rRCeC
yQKYEWJ8Y18QjVH7QJuyz3V0ZlDJOlVF59hDoyhmTv9mGI7SZ9pV/oNRq8BkcVWu
ZnXmvWQ59vqZ6wno9uSp//u6Z9hs0Ks+4DNahg8FtIPIGnWRd+r80q1gWr5SlSJ3
5N3ex55ipnFIbH1TVxCYOuHmApgfJcpp2PBUlZc9RFYsi1Kx7IZewAq036mNmBDn
xKr1HyTCdBEMYzJeGsjgCGBNKXxG+8kqiYIFy1HE8F7Wr04Ax8mLZdAX+8E/LPcb
rCizeXdxddGCUa5Bh8wIklqiVZ6Q2DaLCO+nSyiN+GcbgrxfO2/eu2qJIzr4HKk1
dwajJHsXgF3Z40ZoOWt7LR8JpbGMETaDOYLaO2UqvO4k3swpjVjRtbYLAVgWhjHU
dbQHd11AVr1U8jYJuMyBLthu6RscfRt0oksbbQD2zy3FZr5XBJmc18uoaBiWm97p
fTCPNHGtaiQx+NgjcEA7NsD5J7N+7cxpNBiXCOZJ5FIBGt9isZKNFtA46vaTcYYC
cQ/k+bHqD7Z0zu04xhxRpcS4JwEh5GLeyV7mBzqcOgy6WHoIICXObWfWZFnfolpK
MSMD84VfstNakB+nilOqppMvJSEOl4N35Mi52QGLFZLLfDdHCve/g3RQJY0itu9s
iq9rHPjcA50jBHVU+YwoDdcwaWSjNGkXBx6uPE87ihdqHTNzU+I+fwxQqhOluGvJ
priXTGETESPaX73aeuN9xxXyGcwwr4AxH9bkeuZC/s9MsRO8uAv0m+9Z8IbzRnru
POZR4JF2XATVpta/AVSEeNk3uTxU85ldDAxvEzQXgD9zRQfBMSXDsfVcIDe8Ung2
Cp8qHb+U32NyNpqWIgilqDqTVIlHTUMFjoE8cvhw9RySHJG24dveQcy/VGmj++PK
b3wW732tC0YueNco+HvjJL/jgMETeMunUytYQzF6uJdflDA08VFkYhlg+Orn8hZ4
xIC31WS5WMtk3722A3Wy7bDx/ilp+gT77fOBFEup8zE99TOYNZOMOhWnWPX2W3gw
IAkD/QS1jB8lz0rMvgXrm2tq/br0T/Gw2Cvhm/exGgbDtWRe950oCV64SQv6aJsc
dZMML3BCCAS71JTrPuoBu0Lcy6yZheera+E6trEbdiWkfw7cKlo0E64tybuhlGOM
rnxnPjzgfv6lj4SJmnKG4X7ZN/Rj3csUP2/PJ6nj7+8deWtnkEEFYvWmzQFgkXwk
GcJsh/jQHs1GjW3y0gn2sDXdevacBdARLwUZ6N0u+a2smWwv1V3Z4dtLWbKf8mB6
UBAX+XmkVzmP9Q+M4rcZtQsTcehLFijl++gktwttiz3a5wlLC9jmzqdw6ILPnPIe
42IqqTnfXRaVsiDrijVBnCnB7FhMGIVPTcgoxcjMvdrc+TExWFp9bs4U4tO2zkm3
pv9PjAX2AKgvLHftHz0fnp0boTkBStEWxnzNxI/6nnoO4qoydI/mb1Df8A+bkP4I
wJGAgIKGJG8ydapQvvoFCceYqyqIEMJCM4yUxj1zrQxUlLC/iEn7OEhqDt4szYlO
uh6Mmsx0EqlHEPJowSkaEXlhHZcnQ5CweU2pllxzR6GXU/f8yymZlt1aRftGi+q1
hyrJIWjcgD4F9Et0eYCqRkSBQ2ByxgSLl4sS0vpG78ItX3lwgaBkIjDi6C7JEvQD
WiUAyhRsTXeCIOT5Oyq/V/R7EpmR5tweKjeynUNioNP/+LZJfzOW8dROMX9QcVLz
dIG6gDNo/Y3rqTy4JWDs+NJB4FHLFWwxRBTcAq4LhErAFStfqktIXDnzqOH3gbWE
P5Z0Fa9S+ZRhY6HaOX8CyR1PoT/4mp+lbuJuPFshsiMI+AApysBK7BfRyKEUHxOW
/1+kyCnc9/LyUVf8LGQ8xwHu25DllpvQBidFcMz5CEY008cI9vw7lF9WZM/a4DxK
26iHH8aTN62dWtqL9s5OWP8mwCeDxQT4osScJFOKtMc6yDgeq1Yhw8KoltUbWcNm
7e7bCP1AffnxVorXtHZzn0Dajmz0BDxx93Y4WnDbwRlR6K7UEdH0Cu6fhzvL/dzO
oDIhj0HOnXgomXF8/mooOKmwv1QQSJQ1GqywT0rhkn5p0KYDadXZKlC5/dqcYZ2r
VthUHW29Wljt1AfW+JVWP/Jfack+pNGRo46g00bxfKkbo6BlnymsFjb+9RWYXhJA
3t4DkKqTGuBhhr88AC1foZP6esH3MSU1nwj4fOLzOqKMusHjbaUQxt2qKrEfC2Sm
2IYJCSBaKCUF3Ac13vDCmqWkG7DyC5p4RA3hKRiWAkKXPuf29n6VZcVZOy6lIv1m
gHydLXvl0EEBoNEUjYosBMR099dwb9GFEsN7h0kG8rVh2FuQIEE2dvK+msRm9Agh
QFeteWFn3NJW1ryhBrjsbOadxOAqoyeqGQgyN/w1y4+0H3V1qovfPG1tv6G1y/za
2GdAU6go+ew9ePwFLG2M4XObrLYk6pNLXRKYD4gtw1Bbjcvjd7xZxJSp3iOEgxL/
zM5gXR6UuVhhgads2o0CJ3FGJHq6ogvlK80NIoa6rIAdZwD7eTtCbb7OV+cIJ4DK
S3Bmc1ZOI+ynR1HQJhH4pybvyV0BKD1wZFtLFm+CUlAtJyaUD6CZk16+zHtuRUvg
wUkVcx6XQzOKhW2jWjT6LWToqsPXGDqq+upvu1dSjkqEpxS/30km5eDWsSxju7nk
LEvQo3IQ1fkK0MTUHjsCyAhJEspA/+/DDSZJprBzdkJplu0pgjS0aci8fS7FBrUw
jR6hWHbG/3NJdtk2GLxcj/doU5ZrPWL0kHHCDHioip0f++YiQkKudDFFWlRyNYA8
v7WLGhUDulR9Rb6yJnVGvO8LgDqJz6/e6O5wd4m+AZxNC4atVKlbe04TTOGM1wCC
3TVrGO8pDwHZqRVTDYzZrPqxJtXlBJG3VEqJej37xOT4SVChhAhpVY3yn+frV2WG
PEI5WD8GadIlWOVwr80JqC0MeNATZJAk5ZzZGb9BMWDLLqBe9Cs8Whb/GJ33cR8z
bZSwA3v+NOWxsLxkOrXR/5yvwqmr3jJN3VvGhP+z3pjLQ5n1eURsN1An2Qz/tli3
KFtgBdtsPHQ4tddR24DO1O6IdmpSkpHbG93/yJSKzFguH0LrH0uu/iRvWwbnyunm
uZVmTFKChNDj3LDAXxhEj4ld8cmDm57vZV8IgXWC4YsGKs6eBSGRGYFzxCxiPOgX
jXxdVJQlDhZshcgrLX63NAkvuJrlQLPR7eVgWmIs+Mn5jUr2J4Ln9paryKMQP9KK
sNZf/hsbgXoEaUJ1rnnxTwCwvZ/z4XrOOEPCnTsb1h8DR6TZcJqgoYp6N3ODTEJ+
Y274OEMwEqMQ/dSbeUXAfqfUe1hzHSsj9AY8lpTxDReVAfYSEcpnkEvYZ+DhKyq9
IyV2x+8kh8GpmzTkX1dEY6gJc7bEOEhNuzFi0IbY8yWGAOr7Dn8bs6YIVpc0TQHj
odsUjk3RU6y7+ssUiJXZ9chRwLJhOONaJEx2CykNFIP8qX99EZrQYyJ4lD4rka6r
tlRjgf2btRHWmFaTTMmTkbw9LM0sYvNnwE4G7bgU6vYbuFcNonvb5YXOXSthMrTO
gsqA1fUqYr/wSi3U5RHpxT3PBCfeau/jSqghy+5JNSIgjvTcHu0/t7Ag8inFEMRj
eQRQC/Dov58vdQ1y1vHfMgUxBcEgfQ9gIxKguizEGDCKWLIdCQv+uQgpPWZpeGkE
nWLDx5J/nw+/mzPUJVPZ7ELYfFTmVthtgr08i5yz0JhMr2Nvusno6ygKWADQZh/r
qql2wNZrngJ0VoR6trpfKxjPOG+2zx/owU6RHyms3oecnHX7vWQ8/XdOjZY6paQl
9pFvxEqvbokUWtq9ddnmZ3SX1G7Qe+k4ZQtBQXeHg020+01RlyvDeElO61fogTCn
Jsi6d5l2D493MCa+HvimMQ/15U9K/edmc3xNlyPlv+Bfz885IsIKd/JMs6gI1OJO
UuqL7wTc/Bmwi74zXDZdsTG1guQdz07s0K7oUKEk3D+1ex2nYFzFrSW+P4V36mFq
PVkIwpUAsJcgHu8yONTKSkTedplBUL+FeoirtLBd9ML/J7R8Eft2YV2xVtjROJU9
47wo22Lk1t4WRGkXec8tALtcA88+xzU+XYBTFrao3XZ3MCyO4/Ix+FDFb0NOaxW5
zK21YvPWOtLTzQbOBhEDNF+YyWKemLsIXYp2VSRGB93pWbrftW815JEyuqECpKyZ
68OU9tCCpzvVYGDsfmCagcIAQM1hKOD6/C4v6Ht7bXCECnA5KdHaYd7RxuOV5l2F
jO+UFNKecCeh9J6TAP3RbNVwVG3WTa9wyU6xa+w13QR2InrT8U3POs8wXojBtsAD
kyi6Ex5tWS/IIiZXTaNbfZqu2C0MP4HW8Ur8+NtUkAEjkb8h1LsIJah1NKOOhMiM
9+JDtvuQJzKGqQOVu0p/UDuQxqlZl9R+Uu5YPhuxVjm6+WC/uCT4KrzbmkEvZAoT
NGrp22r3pdJfa8ZQQau2BxE1OIMMbDq5sgmENT7yuawfMLVY/n9uVPZci7PmEvXh
rHspjbrHhZrNFGTMao8/Xdwo578o9FjxvPrlp8x8eJTRSgmbMiVo2d2zTYc9Zg3y
KEaDHZK332X59DJgMBdM6+vz1LY5HPSAEF9qOd8hVQv0krXo4QgdlqoOcsEWiOom
GUm7bZwXt8Ah/vanqfayxXG2BJXHv3Z+RT+AEhAEdVzqaYMuhKrSwnDFHpcU8d8h
vK9vJ01wnh5n5LBNZkEk1i4v+gs0mGWqFg5/jvBtBqsDUs4FPX7GFHdVQ3Ufz5/z
MTghRHSOXZoCAn2otFJ3p7HbLjLnEyFH8VkX2oEcpWRNUT1Aq6+6L+WNhFmHf+Rw
3D46AE99YabUIYtAUwyOp/5QLNUsKYL6qquFb6fQF/Xq/ImHRVNz29WnvwJtO1Pm
z+2jz+zCxVM3Hk+UKe1PPk8wnP/60uMIVag/4komEBQ6+Zxqp0nvk/7UHy+Fz5Io
doEbIGB+OVkdzAoyKovpbTsXU/+bjjJ/+iXBHgPQ6l6usu6OnqzGdjAa5aDa7irX
tMQ4sfMcsw7D/HyAn1qV6/r1qo8qc3yAIbPokd8wrZo6wbEqf3QNhewQ8/yGJ+F+
Sh86DZWdEss2nqVAGSwvFoum+odbu/cDKf7wz1+KAgtQE4cT+WTI+laJjhhO4OZy
NJejETVaBc1Jfzf5G0n/7G+yQWeNKHPX6+pvXHiR2Sm5cRSGvgmlMG/oHqMCqw+C
TmOQQI94Nr4tPpM+ZzGT0NNIN7DIsQJvRXlvL54+w4HYBWU8Tt0fHvd+Xy1Yq00V
Q21tN6YvXP8QusNwvJnyu7j6ZvTQW/jWB703uCXX0Z57H+joqS/0m2ORbu9YisXg
2F+ilSJdSqFv8+zwSht1D4w0sb7rr3D/esryzdZqADyFeN5AJEec6BVHVk8uAbrF
BmgJN53Io/cgzUJiVG8RFe4PqcVKZskkShIQLTtgrmNrbe7Kqndx0iUxlEKl/ixK
raIZCie8zdgy7sU0QEa6qXO7aJeOXUKQA2varbX6usZfxqKtzfG7jHuWT/9sGPvB
FLvcb52OuK5qZRMC1PUVaYMxeKEva3CIXZDyVbdpBE0PNArXYlCwqpqZpoeJxFef
ndE4Rh8JBLVDL8QRnZevTl3m+kQhfAJFJYG6fpDufOo4+W1uH5MEgf8bWOHPioYB
nO7ZFPD86Ecy6t9ReEhTxtyYfERHVmQqh8p17zue4KECp5/T+FUpNzfEvuhHKKkm
mGS9rNnSBY5PNnHcewV1qd2V99bwseabSJHPmyjn0Hx78MsIn/ujEz3tlXsvAnzG
L6wEpUYp5TBPpnFupDo5M8uLTggCVtS/7ADwvFWxShFra13ZsWaIoiMrq7cD3gNd
lYbpqRbD1Zyd382Tmlnh+//qDFtRczyVN6laAHW1mlvVc7oU3DQqVxavO9Gz4zjX
ozq18MiwNAyWA99/VpAay9PuGFL1kO4goYL1DdygLExB/lyre2IQ+n1NpYK0m7NR
DlhVXzattIcF+oCOmcnxL0JSQ7qtmx5oaVkR0/NpQ63b4muJsW2YFnXG3ThH7fAB
QoyNY8UBzvYBzqdIww3Rgxft5xzU1j8PeqxHorUv37sNnk5hx4kAdQ1zHTAgKjYU
vdHOyPyw0vLYpIyHTOCKbyDfEsufvhVxYbfKCpMnLf0n7jExf3Jyfmkte2l0928U
AZzVFisvLPxCOYi76qCMiQZRIkNMvf2wPY2W4qxD6y1m73gXD4j/cHQsbFYkvQIm
D9pyDXsfxxrSvkG/Uba9XMXvqS0XQQJGE7BowIfGvwsMq8sOOwsJ85zgLs3LX98V
wTFkDaKtsc6H9unhME5y63Ii3y4NCPtjeiUOJST8dNSPaSPVEksHuOsMtv8gP2DU
nMJTM+0Cbe2Tep1Jnm+fmGgsxBU6lX7H9UFVdk/xjBy4lRzwv0dzO5gx7vRxlAQB
`protect END_PROTECTED
