`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MWC0iE3j6dvtQTt4wGxIxX80QJVVQb+FClE/8eMm14GdBbSy6ALM/0BlOS/KbPa
mAA5SXoksW02AdhTBuo85uD/eZ/5MHCumgP2cQpyv4ZLu/OefiOuCaiLcUN7dG+H
cZUomWugxHHKWV24YyzakPDx5jkPQ6i+zRkFg6yOHSTidbqqogLeFtVcQ6eEeMHC
qDqBLEIE1r6C23FSgntOGCn+cW9ZUmvdQdM1EyPtwvIEQ+mFYHghs7697K7t9v1C
tq8r6kkBvyPdG+xttvaDQdoaPgfLM2+DS09qqIcqg3j6nzlPjhZdpeF7dEJk+B22
/8otrNkTwQ/tHLzKwUx4Treydy6w9uQFk/CuQfhN613EGEkuJZ3OsnmUlVb/Vk89
A6+OF2aQs0ehSCDILFjd0HtkTBjeZns5GD1D8gFo60Xzz3ijMIfdwYiTf9YuAgY7
fgYFlQUgGjyfw7HUk28Cw3/u+r/Fs6cW0XMjHZne6P6PIOMOk0UEJiPbNL7AmKDA
lAlF1KxElPvsplnFbCxuRU3EjsefKvX986ozSZsh9DagML3bXsEyzVjltTP6A9MT
1+MJknYgpcphX2kyF4A/NYDxUfYWrTUzzQ+ObLtNGIaqsQETe5hTWXQ2le0BdHGw
l9KfYvjWUXHIcejBKQ11k7h2vJQrBqauHdM8XZNAFB7qJ67Y1EgAx2DDm6A56lyG
rHyM4KQrZ55Q5dPRi3jovLv0//II9wU5WU5fQ/FubZ4pM51BIZc2+d+KL9loWh9o
1Rew83yk8rx9tyz9zMnEGfOojQ/W5Raq4dqilJC8NHrLBeMrX6mdnI21K6GJvZbc
zUWynpPqFRRZ/SfQixOl1+MSipsMsoS9+rHToxzXmBqAu3CtG4sZi6g0HBAXETbB
DDQ6EF2XIDTs0MQp0FNfgCPXP/sBLK8aMFi8RDVQ1NhIb3bPNZfyxem9bRrN0dwO
bY5PjmxaWOQfUBEk/jeD7ecBE2Mo/E32/nwtv73fLjeG40lSBiLZj8gUpZWr3xGJ
Y2AQ+Gs6+Il+T3BDYZRYQJ+H9iYNVAXwqJl70fMOjM8d26wpoDwwtRMKD2Ujhw/U
ExbGepv2ieLEBevdMSWNYsRCVxP4tSXAmb+fc09bnXRxt8xMrnzLYkKFjC+mFOVd
v8nuvwYOqUqOIqOUgffD+uo/MiPLBHjmbX752QaRYKVebe6Zb1DVqE+66CbeL+y0
2KFfce/YvrxBSXQuaC085wycpS5gBy61eRPQgTO6uXtTezUUrwspVPUix+kDueu1
hUkYhrGt6V3plmDdWQfG2p2CbCZ5k1qGM4U8dTkjSN+w+psbv9PEMNzsQWI9qnTP
WvRweNNubbhtBel4PIMH2J+9zZAKtBOcNpxmDUDdTw5MsUHWFBnHvQ2vf5IPoxa8
rU6SVwQH3mZhE/zjv+wcKVtJfn326KVcSJA8WUG/ei1bX65u2798s6281dFHGQC8
mBvAQ9VsX2SZGS2G64lmpFMZE/BLP2zP/dFU9r0delyLmYPdn39QZpLY+kZxtd9P
reTdVnvxgmdIBP+BkF4jnxXbrqnFFsOCaNvzwQjEUAIMd/jc3oKB4uW+S1UJlBmd
8x6eHYHTaSKa1M/AORAN+Xl0NMrbEp5OPkVMZj3Vva1N2hCD/T8AjkgUOhgOZ1D4
+Mn/P4581/7vPQWNZHJWsP+H9izn/4KpGsSmB3PQzpnM1ygsIoH3c5yxnNUPxQi/
ai+tOI56VOi90TyNO7j5jQg473EcatLtdR27CzJ+5Nrd6rHwxt1AT3/n2/keiObO
/cVY5VxAYXFcQOnzm7VkSHcUyj4xAVolCfcSU5vD92QZ+s/Q9JEh3M+H5l8zq7tO
EZcb02UP0RfVzpNGGuiWssAUEuYQ6odqKGri7rSls2/05F8WdToGLSXgsFOHHsru
NpJg11rewm46lG4PIINzdixYrEHGWN87g/01fZ79ya+jatCz4q036fTlADE5Y0SV
GlbtvgWx9MIN8tKi0wbbf51kQmK0ILY8bmsCPDwC/jtAGNZd0EesX5mjbeuadmt3
BDcF8YzspDjRY4aviFWyJk1ZPF6NTsNumEvgt+FwIOZDcoUV1MMXxchxX8ts7/Xs
SqYxAeXIc5YAchsQU0yDq3RE6QzyjStUWezROnKPy/wnoobvZGvpxlFjKjYXxRiG
i6w6IoP8fcqZfj1qhG63Rx7G3hW+26AzSo6AH5+3R3PxdY+DDBbJnhGwUJ+IkI3Z
RqWL6O6XyRkMQN7Ob7hBFZHBQQ7Yhli2ooKdmfHlsKmkxoZHFG9EiXpY2vmupDTU
nJ8ioikI8gyLtyqv0CiFaYXZZdYrgCb7kwbTUORwXc5y1JABiYiGJZBz+zaxhMuN
T2Xt5cdJPjwNrY5Igp6YiOywyHY0rO0wmyEeg0gA0ZpdjoAdb7NaLHNGeyD8Pw5S
CjAjutjbhFG932SbYazMKoP2bSf1VcyvSxCEPbDj2EU97O8bvmLRamQ7ZmSDFaWd
cUSW/w/e8e7cce6boJZBOmA7hHgCsxv+uwoVETYoZjTihHXkU+2grPzhDvZx9UfK
/TkafN1e8mNRSQyMeDkDdKG9Bro3clWpn6I6UOIjzdwjRJTTXNIV591AdvkmJZxc
kLiR765vkziXoSiZTHW2KxUCvc0j05LsyzslYVTI/8KLdw6hyji2g5F0P8qbUrPr
sBqZ/y5YBbPpTEO6j/HH9Rq9u/kKIB+gMqq0uXOYNPIpfhT8Ii/tWYDLgrJc4CYk
oXcqJ3TLceLiw2aGGSHJDIIjEcXt9pczyIn1FA+UrMSX9XHnSaiLp/x/sWSkZXl1
ji8R+wuEMBu1w8gDQiuEXGpKC+szGaqmH5J5AVjVIlW2W90reZFM5jzNiMNjwZNy
SULxRf96BKdcyn4nHArCYxr07FwepYsZWVzQAYrQaxqybC4Kk3DBWr9Kmdrlcq0j
+FeDqjP2KGcWmUSYRpiPdfeTH7q8e6wuVEend7dzC/uaxt1IK4KMStbdRYBSROiN
//Ihz1hhQBrxRR+jabsT6bhRqxUoU9S1dUrJZWcBRxcW3RF76UfWfzLoklblzzBq
hvkOs5U7u1BjtjsAuQKHS22SkdFiU93HM8q7PwuOQqxix23DWV2n8jSL7Xghh939
XVMcMsB5aozv/6bqXPVyCqdkrjivOWMMkgblwfP1pAVsjcSCd1MAQ5cylHktEXJB
Ysrf2sVXQd7/i3jpOOQywtOg0uBxdqFeRxQLamiExqRddkxWO5mlXAFNfTty4dwf
j0FtqASxJWAydQ95Fe/hC43ja8KQccj9tM8sx94VJ7QbV7qvjRTns2LpPqGtBCUr
JC1RQ0nnpor6hhAu5LeVxL5jX1iMv9k87HGw8yLS3sWwVpQ2L4rP1497JmacpMSt
31Mo/T8L0FGizUiDk/F7Ow6bv2FumhaSJWdyFy7+02sbDxw0fTGH/TX5Isqd1bXO
t5gedqdD3usT3Y90BGZXh6RvkOdZAcz9H1OTGgfWx/fXT5dvsDPtcEswmY1kcpOR
9D/lkMoT5m8mixaBTdCmRmunx0maHC82n97T9xPPYs2iqS+kpx0FnQsn6WGFk6oo
ky21CSt8MCPFQ+jXDf3Tqng5oqQBvgXOeYR936263gH+Z1oQ07hUaiQ0D5Ro4PR7
vHaMR2zql7syoyEcmGSJTTXCyQBzzQEuc5p6BY4v5JRQVbhHeuOFxRLFNJ/JINkO
+Tb2hpWVOMD0wJDiVb/YuLauV+u5cdigJ8Efj0HUT2FGx4Fg2qiU3M4BYsEmCwDa
ftSeBFTgSU9fNZSPJOqQwleQr8JTOXcuO2Myy4I2tluRBx84WC4qa+yPg+roCh9a
B/ra3GwdiXnBZjqrQwX9ctSLpEYhUpBnKFpBMFVLPeeauyawmQ1Vq7GH/a+j7kIh
WKj3QKdU+Iwf7HtaIc2YMDtlm1kHf4xj2SGrGXiF9Wnd9z+7LjxHFjYhrLdoTfS4
aIjLgftR6pAaimqZxh0NJFkvETzCPzcM1Yopns5AXsdAnUqKEBkIQPxotRImMWwp
++HKSooybG70dT+D9hMVBA7Kq8ocDBAtT0oInYJooMmoRHSyHygxn79tgmMP1SEI
xumsxwgCSSEgetYdU+3GtyipYsFqwu/L/yYLP8LrHXJviBRiQKFR04MumBKk1P6C
ykI27lSHAsKEZGuHgs7y/xscSQ9FTDtcYLGpnukUefOsk6rcgznoCuMsNx1Pd1Qm
gq92IYJy1PYd98HP3oqpvuKZ+Yevo97MdeTHaHgU2lvvj+P4c8XatUvE7zYRyFvu
Jr5k4ZGumt1KGg0eVSK6ipHZBiJfuMfQBkL0PzUgN0EE3YMDAcyRDxoNEmEV4IYg
bBcDc4zSR3NHdVJVZ6aq4W8Z2SwmscX70OY1IiY5j//Ujsu25NDe2k388C557nG0
EFtjSxIIKY9ycucajaXRUfxbHE6+rolRChbwaOhBZGJVx25soSR7VDI2ImmzLllK
/nbx2pQOhTqSk2DFHS16fX17B43BziwLfkfAAdeqhuWDrY2BMHnkM6ETMvbLkGy3
XO3w7wpSpDQ4LylNyOWWlsrvlLmkWAFE47HcrbC66zvp39d2HDv0k3T1GyEhhCKi
KoaPEEdfFb0Nx7H3CrESsaA11xFxsHi+9xjKtTna4t8Zu1RPMK/ohriNh5gPTX6H
3WO2bniRDavAT8t806bLHtfA2dLlxwj4uHRnv5cIV7ZrzXyB8yUnNLrz+lXSzs3x
fMeYYicl2RZQQKcQ8LovG35AOvlS3uNBP0K6ekfWqw4ZmGcK+wTr0JRdH15qnssn
ALH0LEqK3uUholK8l4n/0DD8pfaZkPKXR03gIyak0r15sMsVbo4XICa7cxtMUe32
LDJ7Mv2PzcGYu2p6UbrKvSkWUQHrEHCfcm+nfbH6XXaXCYLvp7CLUOI0UZ/4opW0
xD1eeHFu3yyTkIPAZyOpWkyuzIf4RiC5+v2cuX1DqvWvCy/lAvimcfqaPA9aGFC0
BDj5KXi3Lk3tG4XjiWDfnW1E4rGrgq10zsbPv+HW5iE0rWpz45oIFW+Axuc68BOr
p32KeTVbprFYXrecBNg1kS9w2IJ+xP378xk9z0n9rzbv2zMcH5q2f1MUOObO53Ef
Dpzy+p+uOdkgG1/vUfK6r6YCYeR5iAG7GYDSSJoAj0fjUEvw1JHJxJgmv8NRzKuo
HQDv/ynWuhFGBYnHtAwKlxM55Z4OyxNbaK1Mc+2BTUtNyQicSxYe5ciyhKJJe4fm
UP42hLRI2QCZVmoqXaQ5GcoZKzoOD3T/2xKH0v/Q5nmgIuF8NyXRtG47irrpKbEH
zkRdjRP27OSKzNr5mi5roKKr+EWPzEpws8cjBsGXUo851bqHgtrTlsyBRrB+BjTh
HKmw2ctvMozWCJJbXCesf4yjAHTUIevQhOjXTtlYOJQTvhoYEwHnMlin5ABrHirv
6/UP1IR7yOQIsBpvzheJxerV4Vcz2DDy7/o+dtz7RDFqtTHdI9mLF8Bm/l2pUX8v
RDPGHFYOsbR3u1ThMLYOiSgbrCDZ7yp6uhUpdjWwjnzQcyLmplMMbJP59tr7Sf1N
y3jx6kpZI2B7ei7ySjTTJrBVATb89FQNTtG6xYb91BNeB2Ib30DSEheGBm19XYFv
S/xE510P/+difvNvKL+qryGIK6KYney4q5YEyF9sYsSfoMA5juBuZRtxpM/6M/UA
vEniVSiCPJ7Vrb0sbF/NeY2ZBf0K1W+fohHn28rkJfP0Ka3x5+edLJYYP2MayrJ6
jqp/BOV5eFNlCUIbSldw04E3v8Pn7gLNgSw7kCQJZNNP3JWTyw2fubvnIbMAKU8i
NGavsTTJE16SUK+4WIJkettZsyOIcgVI1RxbOW4y49ZqlgRVX67NGuYKhyt9BcSc
y9sXW/7aPsOGBpIxUttLHMOfrGRhgW/S5xlZsAd7B3d+HGAA6i0xtkdkO+sSFVWE
Jc5o3aoozkzCyScpsUjwSg2vbzhLNhckjwSG6idgLZSxOB6i9Z8uZsLWjvNk95RV
wbwWcmucvZiO2LdBmM2Tmy1ZgWbJGVeBx4xIWCridlWp2791iww+Fyq2j54kPEpg
c6qgYl81cRiS3CqPhis4VuZoOYoCeSiLpUyso9QG8qRnIyV/5uZOhCgYaXk73Ulz
T8HPG1WlUWuTqxxcENZBle/Ve6BDeAftkD1iqmcYXld2LR5Fa9qS9oKflihFuA+B
zdcdM5wZdZhOskyFxWXUBJ1L/evdw+GiiMggeRgN1HTqzYqUiTb2MhwYLQqw8AbO
ytS+tgznHxFFPeowRUfaip3pmIbGiXoFk8Qncz8maHC2cVNCM8try9oQjbpDEwbD
z327XAp/SUvFDFBv9dRZNUZV6fOLDTYQbi2KVm1zQjaT6YzG7ezp4VSWrBZQ/V/R
KAsBfNf+9OpWSvWIQ+fJGzmgd7SI3SekSS2DnrJAX+/y28dkKer8+xBBegQYMzp8
1275kk7asrM28xWkpAUysV5YoGbGsscIupVxhT5+K7kcn6Qe+9BgOIJIYoWqe8MS
yWZqM/spRZ+5ix+NBTpiEEc7Qp0kzFW/27DNcD6U+FI1D1Y2jHCIJvvs5dRCC5ep
OhiIkqWidBubyG5bT8B8ZhnU+VZTi7Bfs41yKY9G4UqwGyhS4gH1Fn65obhrqZKA
ggOt76cQ50VQnqraX0GP1C/fc7Xa3sCM7XA3FlkOePmafJTnM3uRllyt4UkWh/fb
ADKURyyWSW08YJs0NUbZzLG/mUBcPBuXo/ut2EpghS8ZxgT8CWmS7GsDhaIcM673
pkShNH7xcBEJx22Tru8SvsaoVUnWTusEeeH1M7QKzxNH+LVrQcBbjO41EapJQc+5
+Y077qsQc1kNYO1isGcFlkBubzvxm+1Zfj7G2SVLQR7Rg7Py/zaYhyKsSQSvT7JW
0vBsqQv6PGkQG8xzA/nf2CqN2LDPo0EhrXX9EqwGeTx3vo5O4disXDMhHjY9Cng/
+x3uPCqJwLKDAKptwqWBCKXYPNU0jHr5kIChI+BlBr2bCmBg9JlyeCp0C0Und2G6
uuOCZOTa5Kr+OHBn2z1ddbyUrQ98JOKS13QwysGZ6dOU1yCogcDUJh6XURrOgNsi
ckNdip6mZ1ObeZ3kxlBVUb7tefzN36Al/vjcbNNwJjUepK1mg9KlnN6duEkihy5t
vIizUVvVgQK2jZP/+54mw9GHO/2Plp1oIw3vu9AUois17otJU24fRkPWV0V/RHSN
K4joaRrQBinfo60ddMlj9dq0+651uJNU+q4UZsrB5fWOxu1uhkSUwS8LO1wE9QnK
BQvztOLkcGwzoLNPKDvDtwVGleM8zVldcyQLY+s3PlFs9YkPvOfGjV2DayHmT5aA
FTfUS+UuaQYzGSpLshyu1c7xUiMRBS76fiSl8wRAZiZ4J10y4knkId3nYAhc5Syz
iX74DRb4VnkUE43Tvek6MiHFQDYG481ib5jvKqik5kmo8/KwZzSQq2J7gcVdWdre
+AhDcHUUDVyCEvQaHL/gzneW0zuCin/LZiiBQpsSyMSoDahSJAKfe+2oAFxW4LTj
MR2Mh8kEqp9UJ33H2GkaPXmObTPrC7zYaXT528ycbB4auylBpmZmuQL8uOAAtrqf
1NMFXX4pkWr3TTEUkLEWiJ5G+eINCfPjM5GXhlqLAUMQIgnmiXP/KjtvaoNsTuE0
cSw9p9pvSCcmj3G0vWNullYJHcBa6iItrh/WsAAPb00XE1JEwXSPsbZ/3t2cbZBN
ksmCuuTQEw6vSmbnDLHGcEfF5gtUG10DqBh4qFz4lsOswt81rqR3LPPkuBrIZBJC
eFdl7urDjoeoq4GqcFksKFEB9Pijw1VNJjPDQ8IP+YtFKzjEDlKrvn43EJ3uvHs7
Gj4nBScL6ECs++njn/uZBYxnKUNjcF0UeQMhNK+8psjr15aDWzrNMoFJS5kmDqoY
s1cFTvoVhG25LfWbXkKgqb08aw+00XqJkLRCXOhf7j9AQtKr1qnEIiQSByp9NAN6
K85EdlehzRJLdNBX16mNN/vo8fXKjjkUyRQt3ldzLCsadXq2zXZW5k7GcEqU2VKp
Ur3gYm5abSu4pIsz2EWBs8PmmPyyOuUQqyB7Nn9clgFm5cqI6RcVKq3VQCCh4jbw
cI5+EY1TdkY6wECAAWVsYnMCtN6zHq5auCcDgzf/HF0fkCmGQsT6f8ox/XunJtJX
19OOIPl+dXtyG/YuTIEq7O8RrHxF3JpiXtxVypjBqLEiIm0JP0GBvx1O3bsEc8sL
WGdoqb0R0PgYP/ZjFq5qPJQr+aFoFwVl+fyM+QKPotQg6swUlh7aJ5KVMIn6oBNC
e8q0q3tVGpWWziekvarrpJLjhhOtOhU/lokviWl2Jy5yTPri7E15rP/fTvSSaGub
vNkG1Uo5p/Pbqx73khf4hgcTNQtFXerZWfgmuRUD1Bb9pzNimNKBZKy7dtJoHHQ0
nBvxXdHcJUc7t+YhWJSs8s7YS7qFnlt7eiPIhClFEgXxuUzH2S0uC1e2nV6T7Kji
QhcVtgvQTk1RzdQio8Yfmip4i0G7ZDPqXmgFAKfDNZ8bSdtBzSXARcUBirrGS7Bn
oCanC5XagWyQ+eW2UOTZRVrju/hjzSd6Lk8g9YOfG4XWs2mZ/68aWohLOS831xXS
CyE2LA19m83LafXva6hUhLvuzYivo9RPdmi+zMzyK57pi6fwtM5sy+8EE0HYbCEW
P67TwooqGvtSvcfrvrZUzF59IWhmhvuIb6UBELPtEnwFL/gmm9w3OMewXgU6JOTB
RjlnJ7gYz/78Rha3mxxMvdtuKAZQ8MU7SfVa1sWc9aR2YQkcpM7YctkDRtZadwql
z3xKCIcAu4QXDr1swdhMtcOVyd40mjyh6epqpbW0XNrcVzpD4Z0Bp3HuXj0o2Y5X
HJ+eoBrvgxjrqjzkAwLFiWKiNCFUG3inbLSvqqCp413xbCcqfcInLKUTyMHCIQqO
+BB3LZFPT8Rj0rFdyh7lT65AdwTYCIXvdNRqcWbb4GJZkhApZUe/GMduY2F+eLXz
5o9ihNpJBDJ3gQ9g4C5aNqNkCXk8GtDAuihqkdKqI66Xrn+MAXiiEZCiUBBua2yk
cC91YMsm5OirwUHtviOCYMKx5sBtwZBGxfg31jGHtVVzdz8dzUGTX3edmW57jFVp
wZrPPnp2FE+CcxUYs3IF5SC/V9pxkHzNy9dFhaIJxL8hoSfe8ue+EGXuGulj5bOn
uYcJNbByX6RY2Q7ULhhRuRnBut8Rwe8lq5kvrguLHsMSsXJ1Qx1AqVEU9ix9mzH0
witmnRB0jdYi2hf5iPIAbciJInG7VJijwX88Xaui2fnWdA1dbDlVKvsXPf9+yDGJ
uJbokeh6B77CN6UgdLy5W5Hkk59zBYHHsR2GrOZjenKxgF5acVsWwmr6ELf8W6eJ
gHxZMnJ99AdPf4ChEC5KKasYNPMaGNXjfy+QnOnSStVdw7dV/GQ0QMWb8DbEJipc
XW+gMAw+QG9ubFXt+bnQQBe9EWvkrNCSh8Ikdji7mJeRqpGJpBW6+rgrpR7K9arZ
mfIJ6aZ+lcEYA1d2uYIciZxlV2qhA6KZ0U9Cm9xN0My9cBL64GwELBqZJgjGNOtL
WtAi6LZYwG9DYjhNL/CUdtgZMH5JMudiGgd6ylH+rhb+wKS28RSE6UiiOaPdyajX
A6DsW4ah4mZInfjrY9yIZObAYtEiT0AmokWlpEyFnvLVrxLUGHbDgcGtZMF41QzH
mYCiiKt0uIWijW+gVKAhA9NTDDS8JyAt8UnoU/yLbCOPKh3ohvPG/ynk0FnhQ4XW
fsFPH3DVTODEyW0z/7Sj8lMpjt0MdbhW7Ge9x+9FppNHX6R/uaaHy4k9h+lMexUj
6uXA+PCcqb13RJ1BQBcPX/cyLkXDXRAyZ649FrBBHzNCYLzTRVIo0vRRG0qZ7kcZ
GXfWX9o90Kwyg9FgB815VEC7q9ELaEv48m6yssb9thRZKdLcXuyALMsOXdCa5FKg
5ENhjYhBcUC5au93bYcvFPuA3V1+v2ulFBJIOUIyQ+F8lb7t+1PDCQUKonGaCBSo
b0+3xSOtP7mA7oxNgqJDTTeYGgTvhVQ7/SbijSWb0pzBK9UW7YTa4FnBQxes7ZOz
IWSzQ2W9TLQ6TAguiokMkMlsU9fAKIs9IpGjOJpPbzfbWjA7LoJ44VRHQbu3S05b
e8G0IA36gTQ7t8j+Q4uO0/aK3WENmApnaypUHvFmCWfIpHHJ6c5VNVMw24c7vonH
xh2uPSDZczL88tIzm3ylj1FypvOVxrrxdmBB5AWZL6lqEL84xY7aZD/29Uc5I3aE
Gw+oDcMHLAXZgtDFwGoxt4b/EEh5j/UHil8s1NELHj+6i8+jQHIxXl3uoIHa4GFu
DFnYWoMXPtcEDSqI7Uei/pVR+MJgpJwOYEZZoQIovfHtzW8GM8sGY8MTWi1paPdm
CZVVZY9BJAHRI6kbPzrxE2cH3g1a6z+Uon3KVE1eABFOgu9OReyo09D6APh9uHL2
5mSKjMqhSi7zlIJ3Nre6p5rcWRkd4e23i+AKaPfnC7F4qxDPjCVlzntmkn4uUlLA
evQG8BU6YbOwVckYrvD6YHymxjITwwLLpFB7HVTQVZhf04hltGbA2A84hePiJ8pF
Cw4i67ia21D2n8huN2WLlxmtnEyh/bEO03XJhmgh9KqA8IyWQ2mS3xmCRIb4CkMy
uvpr2ZMSnNSyEwyrls+owax626xSKZz/TdJ1rPx4mJ2lhPmqnhLxBrtnASZIev0J
tRGSXIATu2nXvrs862Xl7LIz+1x85JAh44Z5ktAJzpn0qdNQipVmt/Y6TnrlCrmr
L9Bg+fNQuShifTEwn2jR0RtPy+P/G7lAxHcjxy2H72Ndh5iuKShj5fEhbJ7MHNt6
5uXZVEHDnkiuIR414x1G2ejDofB+HFZkXmKw4Y49x+0AGvyLtjVQiH64Pchfxj0u
nY3LLOdMmw1MP744DIkBwr8BcqodqvnXwyzn2oI1EyxlQXPUcZdGdD4E1PH4Vuna
aUc0V52ygo9jR/IAIqXuxk2n9y0QanXCmt1d7t6LLRFjhk8GuEWHbL+6IN/jitu6
qmiy7iVlqV1VP5dMFWPoP1/qlEfmLK4LRsWtLLMYpqLff/cIc+YEfTG2g+jz+vso
zW5pM/WTh+ETToavJlunvHz0po2UZUlSzPnmf5GltVDBhhNE2LTrnBjSA4Jg51ME
c2XR1MBg/md+V0VY3+uCiD0H5DW+uHarU123dvZL7D8b/tZn5B1afTQvXbYJWU6o
RMOk4/Hjsu/aYNsV6CgtwyjjIn9nXfCuPH/cyTFWoW3bV8MdzKhHrfAVR2yofChX
jfRyPCY9MtjC/+Dzm7Ma8Q+98ZaPCol2RcmmZM3IzRDNeFyA1OjyQINyqfJvF613
dFdnXA9Cmx9hw4pIQjbB46EUAtyaeu/V7eeOlh14G/zdnvTS9e9wGwxXMHIHIo38
w8Lt/JLmhTRYQam/6IfHUIwQhye4wv70Q4fyZQFkiW7u5L1r8WiXYSrO0iSykQ1G
rIJky2ZBNIX3FTIgb6BS4+De/1+lqaFruN/C41yTJRDh7AFP2lAdIP4VGzRpwE2F
DMRvPtWts7ODdpiM7bkEzFhFQUTUiSnp79uD5Rm2YRY4YgPWqzV5CiaPMnvcqmJX
VOpw6iS0jrcGTW9D3zsLSFNspWDI1zQHNj1/Z60A+z085E4lGVOJACu3VLe8gU5f
XiouIKmWKCOKMuVnLzZREbPBUczIWSL73RsYLeYgp/HcOicYkVWh7FyvPOjpPIs6
92UbQ21oTkN8cjKmQqLAAwtrjf8do3CUa/NR5ZxCZInFV1HyYLE3yvKE4eRK5tcR
f6gieWD0Ki51agpHFrXQ1v9zPuKjfgUKqF4CEUoKOk2wqriV76tQ6B5Oz5x/BjXe
StYbwM/lIiPxBhd+V5V1YZq2jF8R1oLwqXY163LMUsjQa5JS7RUrgMBDCI2ss6Dj
BWEc9r0j0+i5ZzJJgnLCarkaYoOQxj27N1MEO2YBphovw7dkSySphTj342Fdqz0u
DzwF/GpmjrVstyrYpO6IPsss1/YUwQpd8WPz9iv9Ugn2iDafr5+6M5XBVDyub9LT
VbpzYZHXOv5+V5yS+lXHMC4Ew67SASECS8j+u7BU2pqv/ur0WnPDgblZ0zeI6asx
TBYp19ONC49wXsPWH5dF1AwImoMfMFcFtCPwkxECfMnxt5qi4wSCJyB/lrmb109N
g1WapdZGNTwmpiU4gwlAJA2W0JUMOCf/JVeKbvKWQgUhtqHURB4lDeLxyQ3ain82
Ei0dSKOoK8spCnW95WV5LFWl7ExnKanjfzzW+Y0PXxdtJdwAwoi1LWHNZbVMkRpk
ZeKcObUH3LdD8G/xNDiIYObsNJ+Pw7lWn9P2Y700bdrlXUGMn4x+hoceaSEYm9LA
Li+f5vFzc+VIjI1V+wn08FzRKMELyF5+IjRaZRBuCePmAjGp1IoetBNYiBVmNs3D
Ejb90974mr6r6SNyhv++NDTr8iWYTQvANsSiUfg954gaxQtZIjKtZC2Zoi8Wx+/d
vcE90gXEg5BSGPfoLU3nJgHqqg9VCr1y/zlZgH40ORc1x7KqfIQ27WPUNQ9bdoFA
hov+K4eTdZ0uvdtK+mzVGt+zlDex+3as4jmYWt9F6ne4W5to/fyW9u/spxTaSqv1
e0lxVnVUI/oq66zOquFZFg==
`protect END_PROTECTED
