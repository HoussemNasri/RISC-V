`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1W5Q6xnsKX6JCh9Cfy+JoAZWwj+jxrFUV5A5wZRIIirDrRMK2l/RwI0nYKWmt+ee
lnGZD/f9S6gXXKRrVCLvJAOqgnqYvp4pDrbS6PoHgBWw/Xa1PxsrJXWu2ZTHZIfN
aYwbma7rl0M8VhPRlDCsEGlMsytEuri8hsr+mga54OV6wko0T47eUBz0c6TM3i8e
r7srVX6Lg8yV1Tl9lGbaS0w6ghAAUwiBEW2BMggShVnmQf4xIgSxnUzzdgJB1r88
zhkeP3ZCBF5AvPEyoEFT8zxd+j1+dnUgA1wHgq53wrFQy+iOY/hqgjMp3vb3Bih8
FnE3HiUMe2Z9yCSB7RfBS4A22b3O68tIO9fguneLwppvvWJJZNfhBrnnSIVe7ERG
lhtqmr0CpcqKwqe7ZXJGEQ+ZnboJdRbKWmw1Bq2O2Jg+ERJxFaHSwFg3gJkWowUb
`protect END_PROTECTED
