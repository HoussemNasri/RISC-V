`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1aLl9iIY1SX/HIE7zlYUW9LEQCmvuLSiIf6e8KAsv0lts1HQejiJeTdtLdsW0qJ
aBNUJl88E1vTR6dfy+5ldCyje+ZFenJYcWKp+tXQsnu9XJcDdG4gz1jUB74/by3p
l/3wUVA+pm2v5/c6UUFpE+GvWPP9W1JMDPnSG8N2F1cyBS6lsCHtWTRbNBjan9e2
GUbSF/5D6PAQf8GHnTTxubtwet5zCZwLDmv4YbjjIFFLFlXqAscKaRTMUXVE+iWU
7q8x/fmmZpURMN/2qzqeXYDEacpMr7ZA1TJ2EpaEsCR7x7OPgMjOa7dkc41etsYQ
N10VHgSGdzDb8Js92arqa84Z/lZclDSDmJgzp0P/CcUKp/aNu8LgeSouoM9MuJL4
rwzLJbRwKwmKiXmP0tWmukD5eds0I15oWvg4eKBuoO+9EV0BDRCyFpXwbkC1gjUC
2dICwF7CeRJFhRGm+R+szZXj8oe4LqcvrEoSrcst0+JKQFkuD6sEbaFi6OJ+MuAR
ftDKpDkDRnUowGGkIc/0LU5PK3Mopf+8cSivGO78/ddRNxx+ncOZufUPaEEEEzlU
swgJ3GV+Yk1lEGWy3c7wBiIQyp54AA79cXA+z4b9zhtBoVF+BvhVAR/OPJ9Fo+di
/juCSqAWRKIYD9xyFjQC2ADTpLaDRVrQrqWs9byWZrqlnCdt5DTMAP7Bk359H/No
u6izUA9UBIA8EtF9Ng9dkxqVf5yJAkwfpXWinrjRNAmOlvnwSDEQ5L5B/iKPgqwF
jISogN23dB1s82QDbJbjrL7r0USVcQB0ATDe7ZPR85FjGn99k369vIrsSIicUMWL
rdeCHrnwdBbD1jJClP+0V1RJB2aM6m74puxvR92+PmH0be2E0qqfl5eKq+rCTAav
kTbztrKyyM5zGtJhLTOX/582mFfQ2zsVOZPGfyMmxiznDZUcyJMUfJsFjWWo9Oyl
UcNYRgmvP+74/eu/jgCkTl77cy1OfveineU5FXYC/sFaKz5hFshJ6P95zj10OB6c
nH/VhP/uLsxICCJ11hOEoopIdFlQJx9HbxhcXxKXChKB10VsTwM7v+5PJLIJ0yBg
1XfdR83iQKaIpbyUmTJ1jPOm9+4BnzjeIa07KY4+I/OO1pBh0tYk34+8S2cnCCSd
rqE7YoRcEAgx1/TVdqNEF7uGgCuTtDHw+RuYWNS7g66Jk7JzWBaJsftABMkInYlj
k038zwrlEWqlMf1NOs7cVw1oO1t7NE8Uam0UJe1BecPHw5bXvwA5FPRHUbc8Qb1Z
jbbc7PtPflR/Hiz5Q4UZQ5DxiF3UeaQVTXpgHpWBBR9XzHhoQZtchy00kH4oKB3E
WyUSMg4ojdxEa13g5vw6cAHHtc1l+jq8r+TY2Y9cAobockZh00XiPbE8BjLGyYEF
FymgDEHZYZCvCQKuER62YgYkY5jtrMM955DADK0vnPdc0hFg8U3DXaKGVxNQL2ap
f3VBnA6axU3yOM/StkCKzUQRNoUYeABnMVwrpmAix7PVQ0CunYjK95gJhhwvWTp1
b1s4sJmWwJwgXdFXcrjDJfwXRRf/hLhzS6zRDtVE++Y=
`protect END_PROTECTED
