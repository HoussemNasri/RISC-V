`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Mi7dx34lDq9T8aBbFShRdbr+cD58+Ai8KWjnbd1XxGb97sB/L3fe3HpSLc0oDpW
GQqYon/ihYK8aBCoOHBHYnCeBoh1h1ZfysHrGmC36YMcxVOaaz4nRiMF5Hf6YqEG
N7cFf+8KpspKq1iLFxAecUGleMMGikatyvxFJg1bKu/V2CyYcrjQpN1GHiEJccP9
qTlwLFyhWIXqxMSdozn5rAkbJ0gJBsZTTMAPnjdAK7WwxutCFpBMx+PZnsy+9l18
7WsR7BYfJwf1VcSyXgUC4Y3PY269K5PvtTHTBZoAu/U3vwUA68tU93ey14TXLx17
RhH/k58ltNhxA+1gMyziKT6o4sygNmOJoC29NuV+1GQ7tPO1uG4HQmTKIMn4jm1R
PcZO2shJTOrbLm22oTkkD7bt+f76ou/9vIu2ABduZG89AcghUW2RX9wXceojAv+L
poVTX76FCEUT/Sj2v9JB3/6sizcd+uWpcY+4ZP9u3jizoRybCvoyFqWSo3GSeDpJ
RnhLV3oZLTT99JJZpBZAM1eHeVu7h2wrrLBmn2FC50UKE6jR7mFBB49ANV32+ySm
4QzrB7a2p5CsqhWUVITI5IoB0DDxBw/wmYVVFXJ8fiCG2wqqvyG+VKR59MZTqHRb
GOxHzMoibL/+XgRIgeB4xuJlscwp7mupXzOZ6+6ahVJjoJcABvJYqNrHvYW7Un0R
TCoMRT4zw9WEDg/k4XCoy6iudcD4JxA+lvI8v5nAJ0avfg1SLVuYF+sBGO7y5S/b
p6JZBZmrxwqIcAo6u5wSRHLj9f6PWAznoccFIuJ87FOey88CNo65Qau18aiA5HBk
lX2ACPo2PUpWvh4f3T0cqurlW7Ml96CLVKzYD51hlMy1c1q2qi/usQ4kvFwQ9htW
M1HZYTwrt0b5toChSElxEoYMG0dH2sGkIH4mIJ82UdMgjOG67NXc+aEYGEHsJq8/
sdku9YI2Qp6K4dzPInRWo6+/+s2XiDrCOqeWFwpBukqYczokcEH/pN20yeWO/nwQ
wW7XvgNnvuLXeCMq09UA0QG04RtU8VK5H358aO7U3K8JrZp1v4yEviAPekHwD/aU
ahN1BJLGiGGW14Y3Il/t6TB9WkI/ApKUHZt5tg9CsdTzXttjTA+jWMwQAGlckkE1
nJF5b9pUHVYLhutxYT9PXN/0LOgBdCJ3ZALn1d3vTyDzFFcXYOSn6WdEo4ZcT9Zx
k5HXLgWyN0fESPKt2Ohr1DpL2SPl/eH5uYtTh4fXNk38ewY9XJSInje0tbyWzMQH
pX0hXakY+zyNs7AgNyYCPOLiLcDgR/5mqo80wNf9YNjdvtzj4V2MRtKAoDwRC1mN
vk/UXf93FANt7hxvFV2SUW6UOHlbjlaufa97yBKHUcWQgjycERG0Z1WO1ZG+IA4p
UHSdbCIQhOH3JJ6CGT2tGmTyOvqfu0nJkP+27VV3JTtu1WxyMAJI6pzrWUpPBuTP
BZ/zcX+H4Yih/lwrEciIUJsLx6X8ENWHeDYpBKb+AFGFDTA74bszE7Ka+TZrg3/H
sxy0SIOSS+/+RmRTx6RHquhT6n7U99O+w+tbnepJKK667jBUjyNTX7kadicK3RXI
7oN3HVDWVx8QOK+IKz9eRioFe60xWARBvY8wsnewpZU9nJbpWULaI0xeCquntl4O
Z03K8P3UPq32LiVC/D1F+UobosJAAieNJ4mQzm+o4KrFP2IgFRnW6zLMf3Z1ikrw
BrQI/oLMfx5mHZoj9BxPD28rVJp2SjbD0TQlpngq/Mu3cKOhsQXOGNy3NbJ/wrgH
NMdoJl9D3XccK7xsVG8Bq4v7kyIRh23VAMeOADjdiQX4xgHGBkmaAHst2zZhI0wT
4MC3azZLd7fAN36JKJA9wEo/a0KEHLJWAwPODIM+j6oinzWrlZi2qf4IpoZsMssX
pVIQdCJOC/9t5o6Lsvnus1ILzcaSzHIrWi8UBK3UgSdkA2R17ekxh9Vq5d/RlsqM
fiWJGjROgql1hH6fdeC+0gMBdoMlUIgUPHrNcWgBUhv84GNiBC9PMQVj+kX6U/h6
1WSDzrZi+SyotETQCTZr/sRh3VRrb20ko/V71FgOkrFW6uKlzwNcB9T3wCP36sGh
rMbbRa5FvpWoq8HtRms0WFdm3sXjjeYvtQBRqn1ofwQtMH8yDh8zIZfyjSGtyJTB
KOsrwcMN9F1sr111ITASMAfT98l1ApPNue2kbMDapoGH2i2BhPaoxHCmjsg/rIpa
b4GDdND8aa7dmIpNI5CcnQVoSXIsSIuc42XhPkfVpKigLyjD56+1+kphPmHKcc73
OU3kAbE22Brrp4T9yIbSe9JNs5PJROhO8tHS2nAx0pxq6qDRk5mwfKVfvpOVCUag
yBG3Pe1f6OwTTSYET3VtnPK5bLTGJeeC8fRchZiYp42kkBSwKdAGCpL5BR+nwwJh
VZOIVK8dIDrK0MutRGTUUYcfco+pXakXNGjYnO7SBWKHW6HRrefjAz2GoG6QZyEj
cNme4c6JofQnCRZ7xRc03fYbM8aruaVCs7Q3FhSBi6tV6bDyWP+uIPhjoJX7qwZL
+UUTI+GTW6PeXx2o7g/SQahILLk9lRVNlqA76VDgLmhFcP05y1WSUrvzmv51KGGN
r9KwqGLy+UvIin09eHmBO6p0GnzF96X691taOGznsMZP4ZJoal9SRHp2iwx0t/ZQ
UNEdXmdbAJSzndnbMRpw9zc6MB9esug5d74/LiB4rXBUGRnFacMEv+Rjlh6hU6oO
v3bQdh+UEOp+YpynkfmCFQr2WyN8o5VklUHu7rghzlhhqnj82oneWBF4YpkMmvnE
e0FE3GmZMQOIwxMUO26kblbzLYfggU9AWyrni6aWE17LneIinTlxENIFaE+B5O1H
e9dk9CaOVCiT7QMZTNqin8b/0OOu+o3ZvXAuJYNHdcZHU7L09qIS8sIV6oq8i8pP
3o/VEWjzbxoXXJwkS0drJD2cbwaaFHByuJeLrpPMpqpmZtvBaXAHxaT559B8GoSo
IB3bPq3nRcPBy73AU03Ei/Umf0S9y0ley7ag4twcjdLlO3r/u4NDuK6krFV3pYdR
sFWWZN0UqhzyJcgthr68okCV01iQAAkuELj8Vkr8a0fvmCXdblgJCJbm5GGlssR+
zrQahqJ4t/9fJmO6OQadkb+qwTHRmAIyO+hvKQCpWsm3Hx7pZobTQIhxD7IlqDzs
oUsEvq4EFSOd8pGCn9ICb5+XuFpHcqVLi0+e4GZA61IO5D7MRoCki1q4dZ9UPhLP
LSa8WZ7N445w46AhH5MfJsiRJnP55dK4MAXhRy7zIR25ent7u5cFk4w9AW0fbKHv
FbuyTzbByqKYoMpNFVV55H37C7V8br9QT0Pzn0thK3+p/cHX/CPr6SoLuDREbyfJ
tc6MYCjoCsmZpGDhjeio1N7ip2+egExkWkCBYpG3nQYBcc908qhEpkMRWe+t3Cdp
ruvKM9DopR0qtYDVo2HI57y4N5adGGGgixeJoDyPZJCK6sXMr0EHkPIyBXGgkEQr
FHLFTGGKjU3jf4nH3DHrDMZV+X0q7VemaRShwDJdcXWZbZWFsU9rcw6ur4lkWSgu
Xiw33lffUZ5UexWtdwSzWw0gaRUHUQ6veKN9aDTI5MKR7VqNW6R7OsC+qzAgnQNK
pz6AB/HwGIGYMtFLzKc6DqJBOkeQruHY9TVRUurDtDZMNfIlPtAcQBL+lg0HdkPb
C435Ee5wTj/6iiRQN0iE5anCdzJcXTm7ffYDPBZMGIpsjT5ebrHIIQ7dmwJuFmGh
mWsB+MaQlzBW0XbRdAeJI7IcbM9I7+rfRL4k/YODQcPprS4p5ZLH5kr35rRpPtgA
yZswHZbtZDOLmQw8trLPcWOcwmjF1VKqXSD+FPrDbkyii4xTjXZpx7EmFLcUKg6h
1/zvEoo6wymi9N8T9vvZEot2p5HlZbLELEpBx18LPWTkLVgJPoDnlND4s69xyMiD
wcSBXd7kyX1GQmYOvJjZ7qSPJlct6g43G+7ElaQ3zE2i/H9qgRKc1i3hH5RD7aoJ
NMYOZewl+l5H8QVZMUVsx8RJN9wNT4xq9C+/YQ8K2HjZ4cN2daNe0BEFXk7jIktS
etYj2TTEtwH8MpRCLEMp7nas52JwtRsLmWS/ihTIbsMEiaZ1Nym5TxSJzAmiZ5ah
uLUuay6vqw9jwWVW9og0FlkssoMJdUS3JKnCWOVqrk+1U48MO9RBeekrB5umZMaW
QlF7zAewHBMCvmB7EKqAA6jNAlTx4voBOqAHULMtxzlKqmzvSEj5hKyRw9bJ3x0J
aBGHfQYHIPkwSHqEHMN0WA4in+9HWkHC+RRs0tCUE4wrMIqvGP0qEqXfMjcE21wD
yxUen/MHYkAhtlTn7lqMKu/sp/LVT7qggCjGoQHH3AaIpOcVVUxFKLFK94blHa6D
iH5A+isHhUVXmZh/cfvVZEBDQN+O3NoyF/jSnHI13hb/AT34oF3cNXEZRVkzxIwC
9LhKEBqOU/pQRBSaZFxzbogk4UI4HTNpkdHcMua7gaOSMwRGunJe1XaiFaeEdHzS
LWb22W5j6YbWlwJsA1lOvmGYbaWqsO7RvCqsM1jWzR+K7m+QMZMG8IuHOLmueRXJ
jrzb/e7sKlNpQijGTZglNkMU1uL59Ymavbz3pTIaHqxUTZuDudAZPyDbd5Y4SM6t
9TMnck3gjWZkfuC2yvokBeFIoQZdDxnN+yJRz4BgddbEsjA+bqVMT62ksWZkX5Xi
n9frqTMAKf9EZBp9Uj/iB34HVT9vCwAbVmS1aoTjDPunm25qWNoWU5PcwzKQ6ZcQ
085bWQJtVmHkUj1BHluL8PsCagn72BOL3Mnp0pu0cJBoskxqm5y993vzAXq1pFSd
Lu7sBRqQN4pXaE0IfG5N/uhWFLxPTEQNnh74ZbKPN/Fi1iVerSEZV+5kWNoKNk6k
GYnsSMkxkaiTTaqNA+3UD0gYaNpLaEc/EYth09AjTKxTqmUt/EP+Xr+dJ2ZSxTlH
F2ei7CXbg7TQBp4ElhHHyiDCyp+cC5yLghUxwy+r9uilVbxs6GtAADegoUqOO0jt
UXxDK9kL5GsNzknJzR8d8P5suoRKvWyau/Oc4oW5Lhz1knR3h12vwuK+abFZiUOB
klFFoCVhujtpocYtYZlQ8Uj4paCrhL7gzuwzVPABwEVb4KyTnTMbnj73id0CgJ24
QzW2NsrLYoZJi+NqPnowUTKH2aNLXH3QQjeJ7dCbkQJVw9/8G2F0N1gnYxmSdcuY
swzDIVW7WXYBPU1+1S2VKPRMPWaykNznw0vejfcjd9bwgKZ/QhwqyZf6arf2CozN
LPHXQKh+pXFonfls0ofJ2h/pXLoL5IQtnL3VHydp7OWCN0+KKgaPdiFD/L2KEm3j
7TIIhUEvePQVNNEicduLilfTcpZml9xQaYXqsra7lTOohrKvYkOZGuibj5r0kJ2K
X74OJS4Bv/z+UbUbKg9grhPufUVdpQmkkMaue2KJ6qtnOA9WuumyGU4Gti4Or/gY
mPey88DNNkR4p4sCEv+s5/G4FFBcDui+0D+Evuxmb5tmdQuoc3AcxiNydLsxHtb6
LdniPPDx6ulqjtU5oOO1a+xH3Tq7nvAQnfE99BhQTdRhV178fM6cHbZnx+bvyaP+
UqjyddgkpJKK3SmjYno2+ZckP9kjj+q7U1cyt3LTafL8g0osOILrpSLy2xfhk7W0
bDWGPgR5jhwtOgNRa0NeRm35/AExkQjWu2G0ZBU+0zly8JppYkvyYe4gJjZeYVOA
PGNlVVwU3RXN9wI0Sa5bxwJ+Jad3LPT4+zAaLW+wCtbFS4rtEUFXsghxZYG8/bwE
0oW9uCovR9zKJdQ6ObEvJSJ09Err4c6lx5QtDYicBN2L4LjzipBByHuDJODBUFOL
3qDUzaar93RLVRshOorUxsfc2TWmRZM/nHKudX4owSTJ6t/f/IdoNQa1mBX/WXpi
ofddTyuU6YMfWyMaKxoBgewtXjRdFs9xYmXvQ0ezLQMAMHfb7fm52fowhPx4PM2k
N7pZEiL0Mg+N9yb2xYxJH9/ziDpQHVgho1tMBNsWYbllU4lz6GZ8ImvMw9nzwV03
l+yAV8eXeds5YwS8FQvALjltiApjgvPl3+3HMNESag/rLBgu1F4dZUHUnRb8qV1p
Jva5rgimGXb9oLWK0txuToMNwcrZX01ecGbiSskQIYphQK7P5SZIjdJmAK96CHjq
BkeUpxsu7tnJEIFdV50UHOeEfuHR0ANup9oMCSSVrtnox/FrLx7UxXCC/X4RY35q
ccmNqW5Fl/IiuZrrD+6RAuwOC0ez/LkcKHCrCOYq+0xA8cigagC2Rc+mJSvNZn6t
UWI2fLbTCEIuxyUbtwHh+mBx4UQCJgq5VEmBJXp6DYNMuO+aWgm1TXjZ69kq2n/d
DlSKa5I//c9hU4AQE25YD8A3gdCtC49sJMu5dVBuFW4uF5tsbDZNaVLJVfGL1xUb
2OZZjXp8XfbF6t9jNbs3GxbiVAAVcqOodTqTyL8TwqUSQIun3aei8e8gaNn+ojIX
8KKpnxnq23TCEUQY1GCJMNGCeV41LBIjGXOZBuWzuVNecbmjje3cpb4VoExWLUf9
Oigen0chD7ZZS/OJeXPqIjV6Ay6BMN7RyfwJVNp5fXlm4nENG8Wr61yU773xseyR
2BnnmuukrvUQtK7a3EK+vFnwjwcB/CRxNccEbCu1mZSLXQRZ1YQU4pQJxTfvcdL3
63Mb5EU4XQS5FTsmVpNJ8u1if/747oM48TF3LflmjtsvTFcsGsgOIrf/7qBxuHph
JOXOgJ8jfapX+U/GrsFbHeJt7Jq85TvCnzvcUw5L7gWdBSjUJt3kcoYpw1/SYj6A
n+o74yErdljtwzp4ifvIJukZzJpCARn2mioOiKXhdeizQso1CPR+Bpzdsc1zRXk7
b4k+etARsAraID7VpGHTK2xX2qmybrJUKjMbeemdF8M4ZuQMU0gme02WfUDvLbhH
s2fRnydKTGQThf1wKuhkLF7jv0U7phhTvkjvOI2ijLDR4ZZzCk9aiAB/pUdJcl7Z
lPb6Uc9dnxdm8vrvPHt/A0OnEJmfIeDOT6hFOEZOBJC3H1u240xTzcBtTNES06qt
yp1zbFxePtOcjNC2UJ/l3WKEGHLz+tc/cQ8SNCGOmVA+t4F6wIu0ijpfkYq9Dg1L
LLXMZFUq5M+cH4SGZ09ZzIesi7iFHC+Z2AxTCk/+PkXlB0mNjXVBF1CmIUYNuZAB
T5JA94kCpumw7iZ9AOUA1Hi3yOmVc1fHzSHjPC+q/L2STBhg9iU32lbjFE46YY91
x0ZWAe42wK9WxIzejlIWVvTAnJ7g62UPmi0Xg/m7Cm9cBeV1dWe93rePc/VtUTrF
f99eAnw8dzzpfTe0y2UawxzxHTeKI3NMOKP3kjdRdFWwxNuSjLphA2MOzEhKe5k+
o/IkvTXVhttY9XbW5WcjA0sAHq9dujRFfSv089zSfziHZh7VBMSmld0Wn2V1gp0I
xNrkLUicdMCW5OtNO6F/A307oEC1alH8DzqSdda8JUHExcHZk5JVFFbTMWS37tJT
TDemCkaDp6VrseHQvBL7USSS+PlILKYyr/QK3WIq81U5RWcL0QNP8gcelLPdC9mq
N7RSwuklzYeeuHbtntaMgzLTV0RcwJ4sOkEmAF0YCFSTMbGUjoSS4MyapbqqIByo
xiynJ2Juloh3nrdUbewoVpkwjcwCUbhQjzwZRyPEhpPLTXqnoRFKYi6Hx5PtJPtL
ruVDiAqOpMDj3Fz8SGHPFib53im8T1OfcE96vZ8CPBMfMNYUUEQGQ4MF3KFAf9br
swP+3vcKEyUBXSvDIlewePq96h1Dz0fL5XveUplBKtXX2LkQYB9/nE7NMP82RGRe
EQrA5E9R/+Mvqx7THd4vGj2btYlwiCBc5ct3kdU8wbqKImZcZO1pXtHJhIgVqaij
EcjDw3652RJBf3coLs0b2fqf8lxaFD6KcRlwTV0jiMNe8Wl2islbWXMS4TehKJzE
QwMzDTVzcbcwddbO262nCfOP7tfXukJVFkSQfCiT+0YQOlpUE8oPqJBYDONJuui/
KGL3JYbulTZSSPgCoctv3b4NTJBSn4r8zSOXOIW5UltVtgyHcZPp9VR7jx9p7e5r
onHpGTyCkEKQUFcqvjSeD+xB0YcgS3QnNzlpchlcqRU665eiVWABv2XsS8NZJKhA
kFo0qQZTSU/ybNNFBYcO5x5vh8gp28oC2kZn+FLCzaDU2pypIS886b1FDemasz5B
pauhjvmxjRfONvHj5/D9MRy9k45GLv7nCxea8vNFmTxip0oYm0nEqdkIeStcQFzH
ixgZeVH+q/4fx3qzQTA9HqnBZbSqZYo0xCtMmw1wgcAogJABcC7eNDBG2xBSzXs9
g/vWGsHrt5BaO3FtDBAxwSC9/ecUOdHHJjd2i/WzpJw3Kz6zSItxi39gN+B0geYf
w4T5LMov1ZI1Nemu+8UvCUcZv/b5IxTk4QO5lVeYDPd0k6U4QEij73WJekVN+sGS
9RcZ3RW9Zbzr3BL/KLSMIBfI7Sr26GwF15V3IO4l51grN/gha8JiYy6509ZUy2T3
udrveVkAk7EoV2sx+TOKGHBPHhaFI9nwKmSY7EabAcWJmuo9N3YL78ZFKnKnfxOM
QL7Aq22Yo2+KOpqAYfzAUjOKdsCVaNsW9gsefE/phGszCcC9SEcE1fzD6KlMHJ4A
vRfRgN1FHRC1Z9RmlzHTn9Z7igUMnnGRAprd8C8snqtUWrn8e6xIGX4umIcbxlrA
+02IGGtSj6O89KFd4WcCdYIZ73qWjzkwJJklQ55ktRp+yQ1WZ706YCiAh43wKhZQ
FdZRzZ77yQhb57ei3CqBTzjsbidgzr9RHbmOYsfe1ofDAxchNO+k6h6wZiHqbdmu
i8+MovbF+lrEmuyc0immkSx4Lm2Fnu0EZkcoNkYwboG2H7KOURwquydFstqwc7gr
z9v+oTi5UzFg4Q+MhbMnL1wdZR9qmfas+/24IZxsZCZ8+/sFo0coyu72IB3D4Ax3
XH3xqAF+FZl6eHFksa39jrLNbZf7RoTZP9POBUxhDlfCIVtUW1RlfBXnZY3L5bCC
6+5YBNg/g1TZjfaKueYRJI6I1+Pe71OTIzBZ91xfI+GH6JrOajI/sH57a+2ul/V+
7V3+DfMsWKeNYNFCwZeSqNCEPUPw+z9PasMjichZYcKamqHHnZDLj+CBwreuRz6B
1IGP22I8o8I8+9/dft3cQpYUBEmVG6SO7vsTp3nl2vsau9Iq3gXdZlnGwdZFiZJn
z/lZ6nQ85AWg93WoOOND/jJcrriq5t2vfriTimaeMPye4YTu3/BDQFdO1D+vpgHD
Lw1gur/DBF8mF+fEVARYeiurNQ7mcrr7m/Fr6zImDw57sjHupc2UfJ04a7q5WVgG
HyKR/4SkkQvpp5vrQS3CDh52G0o0rZSExbSGII71kxLx1XfbwStW5KkILbaaJvFA
5Os6uob+M3Aoc8u6sWSgovs/lJ8wfi/BnLrKYZ6fR8XBnnXbfqcCR6ZRRpfSzdtX
Bq4FqzbIwMJML4bbrZUaAmNzrz/0f4YzDBsAPM7qXUqi3iEpME1F9/BiHzazR7m5
UQRySFRf10L8J24sVc1UUuIwSsnogvfQgD6UsillMFQVcRTqtjxpaVngMH2NneDp
8hT7Cg3oEaBtTUf13gXnG5fZLkayNh9x24zIVmaXpgDxRdZLJji6StHirNSbC9kO
IAV7DmJthMlIT0bds0gurTdMLweCQhS7PTcB/cnXJAmfxLl68E9iawmSA0A52m7K
gZcrAkvHDshsZqgNPoaA9sz8c/GS1xeYKYv8BxjdnoZu1IHsM9RST0j+wA9zULZg
+DXF7D6Dp+PHj0obexgZrRfuyAQVXplLQmq6VXGa/nH+X+d78CwEpr7q7wRdj8P4
aKxxsyatugAm2zx+plhOpE7mUUqK+RwdwRD2g+fMf0mmlOSgKpGesLtT0hQ4Fe+x
2xWN7lEkthAj5D4ZZw61ILb1Y+ajkayQIXqT9Muo3c+LR8fgoMCbQaf7UPIlT2CZ
q1+EzpG4Y67O1xgR2gBXG5GlZU4kRuHq2jUXkAmjdfRKVsCoO2Rapf4ZtFFUYHPr
3/YZ1Go7nxcFnf5aJakRvZOL2tldDBkrLwdZAo/4n2SbibKYVP136WzMLavrQCFX
bS6HNwuBoGHFclf8Hb8nZS91lmvlPke0+YSk9zfCIJ+adggA2aS0QTqdBmdPwqVU
76iKFUpnDNSiskn5Lge8i3VEENEAB56m/3kz1oHjLUMSMLk2bthildQivDOCN7ZA
V3TqAGFhBKw2Rc2t6GgkRp2xxEq5UHt3jJJzBfKp7jIdvTXmhsvH2/1NBIw0pJ7/
luSgG5G7jKLw/sRkVoGYV5F3dnXTRTifkexojkBUa93fWk0lmaiyXiqjFfaGzy2P
K5TfIUEJ5OuNr52mPkRQCskNlTawe7tMBX/uTgcvK0Kq7lqqFax4uv1sGfDQGdUe
uZB0CJwQBF4H+IPYHRq2CavrCIWuXB7G8PBDmzxBlKkFC+8nRQCG2SSdU7ZPB0vd
2WrIZFuTrHK+x2bwZ9Bd8FY5dhJbK/hLfF7HATa55wMwwSpBFtZcE0oK8G1x3dz3
fPO+Vb4wz33qha+pGbj4hhCkWJCSVX+MMDYu9rbDWy73oOf2SgcU5RJVUEj12z7e
6yaSe4KO7Zz+xWBcqwl/GvGufJvoXDT7jyFQoC9RDSLjqW+zZd661IPBWv+FdiML
4sgLEnsfBRPp7yf+TOq8C2NvMQBkdvcJcc034oq+9L+O4Y0RQDik1W3XevkYzdi/
shzVH5tPUdRlpbpix8mtqwvnMdFf8tYgdbv80m93XNSfVF4vG56yJ8FYKycv2pZ2
rK8DDWBLa19CRxMmNZSeo3cJS3ow+7jfUbArQu6p2MmlJ1XKCqTlbAVXc0WRVudc
gK3A6O07r7ScfCFmR6SXk0KhpLUWvP6I44ZsuHtmOyBkLrUE18gzetLX8IfXHAW7
s4609a6ybXruxdl4YQa/cFBRK6LBHMAOOgYslPtbkUsILa0Ws8WWleXys38FU/Nt
/95Ca0D4fkROx7AXMpyWVTo3k+YAcwYL8rDvUXSgNAwb9QiHKXIYn1ypJktlZMM/
a9BqBBWBHHoiDQ8xXbKMC51nkZm2sOJFri5QFOXBe0udZPsEi1yGdmSCNrqZRvvS
rdMceoIwQBYJ/CIjWkRLcHxaYxjAz+2ovkZg+MFVB5kwRTcr/NDPLMTlRZhntunp
x8qDL0BJALQTAv2e03BkkYTCsDaszE0WbFbZk0C9mi3Zgig2oJytPMRyeCI03w+e
VRvP++EhqEOwsRt1BcG6MSFvjEUDUt/ELgBgkxb3sDXlLkw6lzB0L5SD4x2+o0D9
LKlINpJPu0SLBJuIx6s5sTIqvQiiAmOGu50lATUJ8M5y7fkLg/lIAhKIfen0A+SF
wF/oyOnD5Bn7qsSTaQ8s036ED37cd6mGZsJcCPBEqIHoTnpKwmCCxhbtGEYGIXPw
Q6MuBsSGlFvNs2D+rzX1dAOvTJKngtVzFliwUMfmJ0Ng6R3+G1BzM4fR1e70umsT
VeQJ28qFXjBLGBkmKYwSkaOgwmo3ZKJ5lmNH9oKL5uCCTUff995dZqImd0rhGs4o
ayjy3vZL89EZOkUfb+OkX9JhlgeJL7XCoXDGNgzJfztYXmwlJYL7f+aYppLIRGRG
Dpin7mx95mtiqqK8ehpq1pdHMQ4I7cNGolP5AzNkWAQV+pvOmlHfYB0AWo7VclmS
KPDfSLxZYQZ3GFlXpn4c6BsvSitMfPD1NE/uVSbw4zvmsA7sa6f6L9zStaEBLlT3
VqOWC9Llpk9Wa6LdPiBHR3zw9NSceHuWx47sgg5/gA6k9pp/k14ymLNXHfJmIUV7
cnSi8UHXOBl52kpcA47BaEOCKMUvzlTewaZGyEBpcso9lmod6SDi7slq1OSS6pj7
3PdPlg238Kw7BYijw2Q/ewXP90oTqTgtv3SwGTgTrEvr9L/K7PiRsxyzvGj2tpP1
4Uyrv1+ruJ4vUMmrwCy7pTLEu5UAr4/rek+ydXmmh/sJBs48ZE1+F0Mq8/kK7rJg
UDGkoM27c08zkwxojn2GKy/gdlUkp8P6l4A7+9bzFsDbQ8w9iwc5cZ62LbeoDNMW
heMH7p/SKL279pM0qbKoSuaVPBCRrTBjEcWCCb6uktSQmNKSgjXKuGcG8A0jxmSH
IzR4s0v9NSVMYPbxU7Of0xhiaR5h9j/P4T4L3xbb+50ZhFUlx8vpD1VcHCDCI9yC
v2HUx2l3/9i9G8qnxR64Wj80YYRMqJ0F5n0/92kKOCFkIxP3oqBmvzy67zn33reC
jlIy1o54hFtAEqKpPitGkuK7eS/QfdqitY2l9oyMGrMpofXPuV39q2/aXx2JczuA
Nym6UQRKeU7DDCAcQiw+lokYTyXek2ve6VyxmTQUNFamOyravNk2JmA1CDaZV4Z8
o4InBaOAckz4gjPC/HMHePnn/4Djv7aNz7Dt8ezxX+WSCX8E7lrMnz+KEjTH9qZ4
NZOrp/f8+ETWdL/Ru+wT83t0Gy7D0yYldUVMIcT+0SFSB/qIBvEYOLwJc1G7q/xC
rH6kWxL8EAGdGdpUKku7+AyP1zPS+a7G3Nv5mSypts96vVXGeMYswKISnf521WUN
lzF213nIY3sMgw/COzqxxkgYjvHnPc4YERijln5rlp3wkcA/12g9FPrpWE2KxkA5
xw4taq7HM5JNGX5oMUb3SYJ0PRLKuqMiMNSNJkXL2OSwOkDukeHrUpS/zhNxDpSK
xZLzL2sw1l9OOzX5XpshikkbUQXEQ9RaKHe2zeKoFY4EYSCLKLJ9lJ4Kc1m3iOTb
87n5FURoosrY7lngxYBPVIRtIVvz2NjElDEXOlUjIhNAGchtUkZ4nPxwpa00xdzC
MdHw8iAHhbeUqm/FxO45dtAEvozM4qJvsgQcrE6CCxg/acQBoRomlW9dER96cs0r
ZPCNZI/anp6ootUPscVwpmKi+P8fBJil5NCuRXEKd13dBCYvq74DCrwSANMvrEHk
4HYsIz/KQrlucB9XJ7INWZweFzIfORBaQC/4PtxaC/YXRfC+W1wHsuq+lhaAuMeK
eiTztdmzyXSUFSn2LE2S5P62g5MJcSyf49cM3i858KhRWrrBgi7B2/okyIxTCEnF
rSLeg/rOKdmjvS0qUBzNdJ0Zc3ppAoeydp1OYDELd9qGN5iXp2BfDyHdqPZ5iBp9
yj9OyRs3t/1LZRkHv7zBZRQnhvSLnrnFexupth1b7JFyugxq9vpNRnyehijYtGg4
OrLveH4d/0Nyeuc2sNQdkYsDEXeC4doxt/Hz6/ZOpULX7Ro+d1c2gMqIC/IrGiJI
uPvii1Q5v8lJ8g08apb3M5vhmcUKu+ALZjGxaHfI3cytHoIHv5AjNV2cKFFyPRqs
VLBuHioBCD8fhgnA6CaKMO9kotsrsGG3GZI/Uv50k3ZTU1PLBqEOnifLnfT9XHP5
/ASeNnf/YpccsF2KUA9fxnEY5OkyyjXwmiuwfkxw3AVM9oYHyVwkM54DUIxmqnCv
k56abOkuejW3HZc/ODnPBsB7knLL6CR/Lfes46eBhrCNqKPyTmwIDUJtU7q79ltC
hj9DmsEmqIyMib9fg1iuqN1CkLyg1AZVDcYfq8xOcuY5ADIRtmuh+LJNMluibcAc
2a8ScAJ5TRKrhAtJIUqRmnXtdwf/fUHqwtKvxTbgGbjDLPshdduUcypJEt80qRVn
nKUv6qsTCU74BZkvn4p4nWaFDBGigUit46q9vAwDtPl3oUeMvp8u83sbsCPKfkDH
mUKNE+EjJ9vmt12L5MpJnVbXobMUdu/k9QEr6xjqIKsxBM793hm+XGPZSrc3iCU9
g/6rCn18Zc5Zm4rPOfGiKr2q4PO6tAdId5r3gKy7/UMEU3nJZ+8+D8WB830+dpFz
gU7E3UC0/KKBMZQLDWZiu0vNTyekK5IRZAL5sf8E34OhcM7ZIXR7aq8wuUPAClq5
6wAsKVPVoa1OrnRiQdL/XaMTiJGB76Ewt3ZIpoxb3gQYuvYIXJoJC/7KtKIbR7XS
sXGPWtOZQcBejNcXONPGJKJDuOpuJCdqcGqA+6PsKFnw0o3YL6uASsqyToSdl34x
IbcNfovXK4KPUbq+jIkFUfc1MzKitswNssi1H0x7UeW8rgmnSbkxXyoHvk0sqFPS
RdK9qWEEDsAZbgc261Q0FerPRdeuvX4tGWDcKKSF8rDXYCCgXc1RCVbX6k5Hd3qU
sGvzGV+fbAwoJ2qEeybzCEV472c3r7Ebyswz697oSCf3y/ymo+Qmdq2iOGvIsAYm
a+YAaC8l9JwxquadGPQJlct6/Euqbu2R9jHxDSdouNSBL3iR3vGOQgol2+R2aWZ4
xJbaXBelPvVis316CxkSGhh2NRKzF8GXz088RZx0PRkV19nGk08tCrgiG2bbEJ19
3GKY8rfuNizlHJB6c/R5TsTMq4y33eJeIlCi2qh/A349YL7VC6Y5GORQImaUliok
cOiAoLhwHRn5viISNPOEcXfZE4DbQk7w98b7gyKEpUttKBMKOeKdx9FNYgPjVVFD
bdYPUqYPNwgG5pGSrLpMrgSdiwEW986+ba/0Jn7Px3UjTVQOTjJyXoYcPJcqeJMX
wolcfhHWkx6I8sjljkzFsE1vdZ8kb7oNPB4ZmP0vTCM7lzK2Pcz8PmPmWrlMmO0I
NG55o8nk1Go9TVeqtSKYFnECfnq6roMwoDAlYV9EiQnrnp1pGx9cb64eDqIQglBk
zodnKotAKk5dqQSP83SoN74NlM7wBoscQpTkHmx764RTbsxjCqsRstEBe7t/FVOH
AaWw58wtjJ6sefqY24jCpGSIikj19Dmu0SVua10JEyjsSV1EFfpYXUXRWKHmgrnf
NbVU3lLJb1ua8fUiNVmaRwiGo1ETk7yvch+pmV4LSmiljHC7EFcsJTq0ePop6Oj3
eXN4XWwjyARa06eCf/cEQGQP6kevJi+AWwtDCrsoxBjdLbJ4prRSAaqfipq3Mf9L
EaGdu17zZAT3OrOLKr2Un56LDBIfZLdve1IKDBgzCzXW75rLQmf9IpdlnVhVmQB3
snkmQuuPm607cYePqzbLNGdOYEducjnhtvXF4b6AqadEWAQam362YQZI70ULYYBD
NppN9zdLpKD+ZNlTXEra+9jcgH74/iINILK/AkHj1B47U4LK3NrdTv/QzS0yQkH9
i8EnK/SPqLSz44b0RPY0dURq/zEwR9NcOoSjkHKZWGBhoAEQlPaxEQsNMCorL6lk
/YaJ4V2QZJaVgoNkpmhmkK95QVLDyY6G2nUE4nOhY0a3/LRiZIETVjU9L9NEMg+Y
8BmpsQOap5zjM6/rSwqx+soXkZeGoVdC4cqC3UfABfFiLJkDBSTVDgrG6Uo1bQWV
5qc0ZQr7HVOEmzmgope/oenjVQ4ChFKi5i/Ss8GGS6cv95t6t7o/+LvyJvQnaGNj
XgbrepGpDDtxFy3nZ6ZLafEQH8doDZFz6G2Ts+diSgkKsXhJXQ+2m5zZKdxQMKOP
8dk23/n7fyhW/+25LDAFJrqUMiqXNBoefJVZgsk8usyQg7oNwbzr1hEFpHgBjVGf
OX6PTF05SlgZbRCJlAilOENKXwuJEsnhRP9co1mrGFZkhXBx6v/ILrwKH3KXFXZc
w0q7AHvAz2qrXznlrgeRh8agOpJQxy8i6o+b9uJbLvof3ybqyqoSerMWzivhJs2p
3ibyjANdbCO7G/hl7TaibV64S5QIcyFL5FKIlghCjLPmHpMLNHax+QxEgouUc9uK
38XN4GFtCe4fKzat5pvyexTReyk1EtEVRXWLuRsiMzpWXos+aZ+Yt8YVsLXwsuyC
u+BdBGscjgyiXKFVGJCOwCBOeZsnwXqIzBG2Zai7MPX2GAghGRrcwZ7xcWeuQ8SD
WVvzQV9DcYrDuNOYxw8r1B1kVoTCMKMUhCXV7UlewONUk98fv28JIiIeansUCOzF
ArzHY2FOGZQ7OP2vOFfhXp91gLFjV1oueKl85aTumiB2ehsQpS4KL3bvezGoT+4g
2dUKxYUNEGSp9d54tSw13wQKXki5SPaiGik7jpNckrwK1cJ99HQgtSfgxpZqnHCQ
g4ead6UTDMC3F1CZUD0TA+VQgI3ijKrY0pQBpl6x55Y8roZNOMwyh+3AWD4qcqts
gnA2g38h1g0JgG4jbP3wkiJCERk/KHAooHIrRYFJ5xtRckLmOuFCJ5FZqodIqS6z
ZFTrbF+jyRiZwY008Wf+m6e4TdYhTcJdG01fe4Sic7alTrP0rfu6b0JgGv86yO5x
Rq7zvqDBaWJj0tk0uioo9H8jDRuafxndCBoihCltXkpTxOyARvJQyDMVd4brBpIv
1Ub+rMKncBVLzJl3C8OBDGRRz9l7i1K3+ga0wy59iC1SlBW25fnFw7T2F9GXmVDx
XgRL+DnF+8BxjHdjf1jwhU0/RYBYrvByLAZaQrLBE2monT14HZyUel++6+Xcz5k6
Octs/704/1UWbpmhNS+ZEMqBoM9qe3LkluSgEb26VZ5XKiM2/YWc3+KN5zanLFHi
av095XOZOgz8DpkQId7LR32ImRFohawdBH3HTiVILo1IxBMo17E9eXJgA6eDHXAD
11ZvYgjink4zbUBSZJ4fuFB6X9HfjUU2Kna6fae93Tvv4LwoUKlNNE0tPOSlvZ7o
+jOuwDvNQ+szLvSCChXlyP3IZXqqZXHet56vWxAVk1YK6rNXfeMrfIiYFM5mACnK
NeJ9ZwMGAjdfEtIIjngSSevQvTDZq0/n0JNspAHdXbBInEENIIV1nHFQrSaciZp3
eot3yv7nMv+eLj7owMSIGtdMq62iSAsi/o5HewXOlwA3x1cwjkVXhd/4bc+R7tEV
8jSZSEcbtl45BpWg3aAKystbdLnZ2NgGf0a9w87XFfqTVWv3xLuK3efhjcAEwBhk
OybrCevR8VrFaKNBmRFiUUTBr75kqAJdwBcOJ0O3RsN7K6gWocdNJ/qL1SKmKVwr
A94sOS1UNzigpuPXJoxfEcUsbD/1rx8rm+0CgIvHguRQPAsE+J9lGcIdem77xzw0
oprnyEvqD4eTP9H6UnuriUNgSKLdZpK/IfFVWe+m7hNsg8G9VfRIObBAQLi5dESt
k6QTQdtHwRIGOOmnuHOpbxncSAxWeSBnqS0z3POPpR5Vk8wq4tIu2p5S5PGXgqHa
8wNJUBH7xrcnINnZs4OwQbrMbqGXptit9F7ENvMJzDDIoVVw2AMx11P4QJCWOMaH
GzYEAU9KPsMiGnstTjoM0DBK+JAvCGVt9fmykSYnvqgQ7BHBz5yA6kCGEdr1Tg/F
3tS6Phtmyeff4wXEz0qm/4b1x3O8A9aWT48cZkHQf2t5AKPrRSS9cqyNwxGj5ZUP
ZKvpZj9lnl0AJ1de1P+Xb8PwvCtbFeBaAV0SDE2ItDjJSFi0V/whtR8KyLlpwhnU
MB7+ex/ug2/yuvd6RyGgbS7VNX8M4idwqt2cWW7PHpEsL/Jih/eBDGY1PLY/3cXk
3dmUxkml6HqHZFtFW7R40Ty4ryp9h6ZRxP8YeoQMsC8z1iVUgUQBlmFkEADD6lJP
HW0+bnvgBcr0+o/RW7CNWUdV4L6QLHc7G/H9RwoW8JIRRa/Or8UzPqoG83nQrtYz
K34VmRfm4tHaq7ZZj0/YhreZIS/5DlhTf7t9q9PMs/DxdAC2fWzHV4xh/n8k5aT1
fE+ufAmgiwL/xj3jCJ4qCBDRPSrQXtofQ0m8HQJNAMzWQHar8PqdiQR1jXYyg6wp
AYzqSehMlDnMGTo4Gy0NFupOFM9WN3jmZ+uLS8FzHKeATvVd0GQqKy3OETGuMy50
U90Il4HbqVNbWIw7lZ0Y6ZcbTeAWrTzDlBD4ssAkeRfgfLFvdSrjy9BEuhFiWO2o
9fuZZ9uS6WFg6xc0qQ5TeVqlyL77rRgKfb93eCpIq6cby8bn2a0ktCiyz3V/sqix
vlTLUWuY3o1FnUWYDn+Qvv1+CPtus9Nv8YBeA4mJFpKGdsoswwx5qZaf/T6kGGnW
Y22rXV52IIXzeEOnQbztphVWiE9jYyLlFshiU/DlBi3MUOsuTzf3q6dpvewdvKYe
3mBqiwBrnmKT/8CJqcsYTg92otHFy1LrY/sy4gxUfv4Mj/HZI2CGWEaxqu86ofYl
m/cmaTxYZrvqkJl38T8McXD3SpFkPS8fF90WOhez9vC3wa+tZrLOUOB3RR7JVCJN
TvuIwA0x+fGcztFb0Rg1Aq5QcvJPPC6LuikvkkQtBbrF88V0A79bkOP8FZ7QO+rZ
ybmuldCYuxVTaWEjOQOYADZVlSnZNh1l5FbvohiG8Y8MrVOd37t1PiMYIX7XyeBW
ZJug8CKw3yYMKc9WhuQ23lYwc5p3hzfDyQsIoOzQ8NUEuAjqcCkVXjJBe4X5kP0B
mgBnCIRLKOusayvTdSe1ArDxRdMpGGwFSHbUGCvI2LuzNXZq328eYir9J0PUT91q
/eHRUdNExIPST1nUTO4W1/3oyffm+XPVmOsnw9PXOQJl1+t4OLoxgklYiIP5kNYQ
uNVhyXRD5L1nKB7XJ4BoJG8fh29PQvc8iWZfsY2XFazNq+7U6genLz2BVpzX+q5p
liip25gpjQugJtZEiNsW2EfasouPQxOKEnJPk3SChiuad7/5rlD9UT5BcRPdxrWK
LmOSV3MiFfINYAZuVapWNy+Iy9VlQonMw8NE5diOnVkOFNe2t3FefqooQ7mNuehc
k9weWE2ADZVNjzSjMZlze3n8z1ucU72lFNrAZiYs31G/4pm8gZGsAapea0ujB7sM
WUZh2kPCBeA1OxJDs++ocr2DuzW07VsmDezy5+PskWHbE9RlZ22+gQWvzr55UPlj
xq8sXN8n7F4cNArzEEcE1ksJ92dQpslElxZXL13Tv01OwVhu6D+YHDFS5tJyBTkp
YdwpouJTqrhIZ6K8U0d7P9ky1l6ppkAsUuzkOgDKv0dzuTnHOhJdyWpxurDyWHAB
8PcuQDBT2N50V3u2BMmkrzF3FAqXsHD9djxrknPayZZQApTOmt2h+0fk/L54L39G
NwB1RUiTMbi57IUj50adeDMb0Mxk94XH0KiLwRjKoyn5uVIYhRT8tKtsS7GQFo9+
JmZSmN7KWW1ouQalhx4+vfftnCLV0674u56Dq3A2WgywDbkePt+/C4TNKHa3cTFD
asJoCNVkkpzbuB5KUg8ukjSCQEbV3eQNj0r6CqAOlfDDcEH2/7PRzsTRi7bkxE3L
2kp4Tb0dlwR9+wvXLNNGGLF4wwcQHaswMX719ajxgsA6/D4nVE1s+YS3pH666Ish
jRlEFR0z8STJv02ZGCjCEp6qRNvIvjjM18UU44i4NgPITxJ51hog1GTzp7VJ18MH
hmbZMwK6xqmZg8C/etGHRA9o3XKAyNKH/h9lA2O+TcuQHyVJu6yEqMRcc9834z0E
Ajt1xBMOToX9JKrZEQlZaPfq7NftDjf5UZqe5M2TiIoIAvP+UvpBCVR+TWEO1XUs
Y+X1tjCpEpoSqpVk4k4PNRH0RE308grILePvy0BGdlwm/9lkEh7TxKrvACKAT4H0
ygmBUsUErBmsUThLC/rPD5wy5IyTqLialivcrcVpZv3dRttWrmLwW792Vl2JyyC+
eVnabUBarvEcOP1DSmmW8vwOOlByYipdCDBEI/JbZcq32wHGK7sJT5c6ZLt6Cqp8
YEJJEFfznvDvo8Dez73FgpfjkVWJzCBUKdimCwlcC5QfkbBXkYAeJKZ+nOhxoDNp
pwspiFRodcqYGEHfsxZro/UMMRNmLLL4/969elXC6EK7xCW2WJcovq98cNefqu3O
/Q4xBvFWhCQ+OxmaCwTnpsddwL+wQSHCSWlcCMOqXMJanpGSzCBCs1U54bRRDJso
tNJB4uJTXp8/QAdTfWocwtje1kQ5e69p3XI88u2Rgd505qingMk7zz+LZVUgyGvF
7QY9u6QjCwPWDzNknzkrpQzeZJfUO18OAXt73c6enjH3fFzFkwPo36ZuKilDavpf
mCdWcWdkuNrgG0bBu9oWX53+Nm2es/mzTz3BDXF7yF1qVokLZY8VD1yBSaMYEKpJ
kSt63odh/+Dj95iOceqUl1h+SDOLY2hPkhuqHTq3BQgftqZKoc2+WxIUCvKiPh29
0SCwAf+506bSkCg/OgVuH6BTEPpkUc7cRI4Bq07pfoaAps2UlkJ1z3M7GeBGfAyA
JEs97VftULpf3vIH2nk/P6yv858r8U+cpAAUCfsOxhObIRJ1GiK+klYLiTitSjvp
xzpD17lZUgeqNfGo2VO1wtId59oXBirm4Aqr044/LsoTjoW8MlEgDrAli6sThhtt
VGNZKGwHTOX6J8b3KufdDEIe7R23o8ioRntYlOU9YMk2+00QIaFkwAORzpsJF4MV
hXBkMWRXfDlPjW+6uxvY4kmRs/63HZ/QlFCgXEblLmzeZ0i9ZrVRaMlAebjYyaMm
Q7S6/nEULJSp/tNczq+7LpDKmTQ7c0HUyhcJJykfQ7dqWpZynxwuU8u/CDIeaTgc
Cl/VZEixEua46RCFs2W4dog11DOFk6yJgdYzHFLkggp/Z1jEzOeLmvFZsFNPMJXw
bzDdqntBSqEAYi6S577jhSYnuWEIWlcdNmeSQSpnOFa9eb1S/IEzBJmoSycl+VHh
VUteRQLXZ/WTkX1ZQDJN0Q8ean7nlHC3ivFRLJ9W1lS/0aLqyajnOMpTfuS04O74
7nQyyqukkGbvHshfQetnlSghMxclsJL1hQmsu4z+h8Awi7Z9ihBXGzqzMGfsb6de
ephR4hrRUmbPHaGOOAIxbNPcjcx3qBFS5EG7dTN1UAoHoMBWlAjWan57+G4pNRkp
tFVjsjeX7KFUh3ajk/lVesa+0zIzNoOgW2ZDblTXZE+raKy5M+QRoZzRs+8evdRi
EBJby6ReAsskPFk2F3j+898tNykohHHnPphciFWXDql/SoVhwgza5vDACJEPdZoU
A7gfM2zQL0djJ5IQpMN8aoygHseNBZB16Q4yQTbEMF0eGbgCHxTFgY0iXSvgJZMp
LvXk0/19WwTlat7HTV/84faniR1IXp0xP1CB8Xs+fFpu5GE9YixUoYM+G8elHZMH
vVa3vQGEc7Qc3KuO0VCyqgGu2wTD737nq2/ZrpArp8tfeVK5ZyO3m43/PrGOngRv
aG2dJYeyAF75X1O9SDA5OJ/pgQuKlEkuBDWXnzfcyAmGmf+lg/lWjazGcrcbfXO3
yFhFLMwYGVwuskxKW3Suo7lcVtmYcrveANhteP/T4O9UbR8od0upMRdZZ2yRxND+
g7/hIPgnj+ZuUc0CKCzwGBE83OmwIg7dccSBxryhTQnxKE6d7JncXWKLlJj7eli7
oWP7KFf2ELS8AIQK9FQgXtfZ0jazmlow+BsJLJRmUPQQ7h75+XtDgB4fXaSWhpB0
/eYTrE+QTPFUprag4c6zOrNmEvl+Nn5c4htcr03g/VNdaFgX+wZFN7J5v9FyIVxB
87ytWcjQz3GrfPPDCWGVBB6j4DL2CtBKOGKE9wIkNO4Vmmg4GPMQrpe1g+mLYEkv
h9GwyEqv3ua/0+UFPyw3W5zmuPmYpwsQxm0NiD5KACy3rGwD2tkN6vOun7Xw45yj
VNf8+LrmjVVu/xWCn+6zLVlxTw+e4OYTkrAIhiYDUr3Yqqjf4eCeE5OyHqHG6atQ
sWRhxNFbtaU7qenpHB02K+tGIZnbcrXiuFqO4GbgjkilkiOOxjkuS9Y0QzFet0d3
KI8a+2Kr+T5YBDw/MoYb7pEyc/LA1MZsz9yG4LTvQLa8qM1GtXWXky3CJvUDXqrM
y5/B1KL1iEKQm6cQLSh0sN6/MUaBX1WYXSunkelCpo4KZJt5nsC3e4ommlAJ9Vxs
YX3zKHVJdG7C2NfgMRVC/3Vw4GGyFyBi1/DzeVahsluXiZkwyL7Hmx+PG/O44fII
vPqMAOjxrmVYqycb+h/tT8aSXPH2PZl+d3merriX45PjZvQx7wfqmVqMVkGxx1Mj
Pp7vZdrcGU4H/UJX+ZbjtU6LdE4sBPuwYqK2nTSE7JkHvFxZjY74yJVDPz3bC/L9
VKX4ixX0lhEzRkqLv9WxVNKsswXfZjJJ/8Cy/7E4iQSBz1AIdDLCOVRivBSVEA7A
JLbEJ/wfv/NOjaPbPXUpBVhlHSLzGQm7PJgj53lasQilEwVaJtnpJts0csBUoads
KkzSrWNeduoN/FA2Uc6fopPAp2efsoP2sRsZ5w9dmucCVEbClOcGtOpkNNApCNdB
iOWjSafZPFnst6Q0eEG8hamX/rChZ24VJZ7Ce7s5Qbjr0WfdtllUcQ6P/VpwGgiY
n0i4OkdPJ1C9Hh0LCcsXdSE0XpAopIYbA/8egHYIOBComaiwUqMDk7PyqcAOMqF3
ioqJtToJDJ4O6sHu8g25VcTnEEbXAc/NfFxyVzWcQP10wCp4j63wt4uKGbQzE7Nv
htQbcNT9v6iEU/uXEzd7NSPWY/eUE6hM86SjdONtsACiXItwSs44bS4dbXcwxMNe
EwlspNYsAszuiSB9u0b+hcYQ3dYkCTXn1G6pJ5ZBiDNR6W58wk1hjiYkGNqzd4BG
RRqqBg6o840RJAOzhQ8WLzvBv1999pwtSTuXT6L17dmFISnRxrAbn3VGx+soqyOD
i771jGJNjHqJQGzkxboun+kchfmLgSNaDTdG9OKtJOcw86bV7RedXIkilpepMLXM
0URQC0A6rxm4XvpXBb4SSgk6nMETpSW+a/E2odfrz/ta0HPmzoB3nR9yaxjx8chP
T+qBFL6nvDDErw1NPKJ5HcaMEwtOLev0Wgtd3Dl8ypiUStGbO2DXZJiiOv4sWU9u
vPY+etmfVUPdOclsJmkDH5oQyR06lYBCzzHgQhXV6F7vJFK8gKhxRUbJE5LX7ivQ
LbSS3Lx+DXWRF0+gbbu0zbgSchw4ma1kaiXUusFz4M1TuY3ZygFZx/xon+sAFFkV
Xgrcuf3eRuDqsi1VzuUBpuzCMsUF7C/0qQIrpxK+uxpcwoDtHtzahYiw5rEExGv8
rJEshCHVgy2REJCH3uiwGGJBCrEfTYwiuUlgJxJEzcXVu+3aagdjHm81xjDO0wP9
u3mDri6Ot63QwMu61uRlsvyR6fK2ACM54STjeU6SNyX56R96cn06bjiZ4GZRleil
yyb8XwU34fxl65nt0+pFcyQ3WFCsedofvECr52XzW+Bs9vlHTA4/8CGadqMq+IXH
YV+nIF97jve1fq7RaWJZ0zVQiMH6NODrN7yDny0UZtbaDFEThRbl34XHipSTvuMx
GqQmumRU167DcVRTRvsYKUU1WXlLHFwDEaFRci91kumY4RRxRdUMci/FQ+OJaG+S
0fg4xoGRBuhMppAR5l7Lj/SKgs2XHjSFBlaqbN6LUPWQ6PlzwO9+nOXczUh9r0tV
QpZh6vWLiU4n8eei8SgdbSJr+vchUD3i2Mr7sEHsrLvlobqkmVhN1VAVYOKCv7to
bb0w9nVEmt+cg0gm7OS+0RS4XfAwfy+MwX6TC4eF/iDRlrUDFzraZioZ94/vEK7E
u7cpM09279R8vbzGZHryevjhhNVJTUqVnsczLBiWOyS2B46879j2ZARHOANrGXh8
4Mmmy0/0UTccMliG8+zx1yzGWPjL/U+f+aitENtRBjTHUmHbjy4KoCl+2uosU220
TLhmJFukFQPGct/zDra0imO4Ck8e+KX5BRkA4D13jGlzM+b1ERuZJvnVyE1BetbU
KBx71p5kxyCGCnye+8awSw6NqSe4MlP84vuTb69Re+Jf0+xt1HD/1TXsG8oGrPb+
mspUWR/tzQH0oa72aW7FItOqOv7jIRBIxNcaB6BD75hglHrMhH8+xqV1eiR0vi7V
ciaRk+XFN+fep7NUxkzJ5DSfQCF2yzSosCBTrLVzV2M8wYTu7d1MTsQp03PevReO
tCQA5NlwKLhPxNnC/YhfVB+7BzR4+nv5M6qP8hD5v5DaVjH+7synl2Pb7lcxKMM/
lUWlnRv5dypofA+n3UI3WxHuK6MpPpdzd1SQaqpUuKKcJY7Oc6zcHZMFAXX3C/d3
CQJ0ZEo8PIp0XK9vBnKTjvLuiZoffPfBG7H7IozUmCOhsWkOW11osVTsYkF03MZ2
HlEyeLkrvYVDd4/RHpqI2zrivTw87q571Qaymlhe9Asglru3v5X9/j2YCLP3L16m
plc5sPQmwiG1rVWpvdllEQc1iHn/5PvUwJWJAI8EsK5sALljkM0V+x9PFFbL0lTH
Pa+56uAhs9C5UIb9izodlLAY8FQd9fhFC2JC3U7DM2Wk6uX1yzOUJSt9vkX2SUSd
80sBOgdnQR3uVCjF2910dM8tHCH/V3a73wi5GFWciTL70HduAysrKKk0Ni8H76hJ
2ywDAoOFp3dpgJuy2aSYIoP0v/H01SR4cTRMMbKktSARgh+6D1v+VdK6YliClxnP
mI8hhGoQ+kgDEs2SxPJJeJoRkQp82huxxUczD67jNly7OeeR7aUBP4YGOqtEYtT/
cgAQ9zPlRzEHpeotHdde6tbT1r8SBeYtTVQVc30NryRCqKxtY1+FdnKYHjKAnKdb
gjMavzamu7R0T6B7SH83xiUA82kcDA5Ws6FAx4P2EoLTuu8tiThKCVUFyh4waYes
+wAcA0Qa9L8D7Q9k/PmrDbkwNy6jh2sHM4cRk4/deOeXwaIJGgD46mzcplHkiURk
VZ/9FXJkKIf/L6zBFHlgjrQkeAz38kWEt0kVufTk+QnroQAGia9ahmcdGRkKB9QY
AdaIIMbRKr+llqqKBNhyxyRlCXQdxk2I/NMZhJCBUpcO/X27qWVptfrYGkGLXjuW
KjT82R2LAU0J6SasLaz85EzGoe2XWOhbLeLIuSMy7SqjED8ZYvG2UkPRdIwBg5Dc
a++Vyne5rEd3FGVRCrDo2L4/TrHaVPTzLlEmDB5HFlUh+ZHHLZ5a1hfiPSPcUZ4R
XAfBFucILjaXw2s78O8h3x88F9+t3+2FiRfe7vFU1QsGOiGQSwBy+yr0tOHoI36M
xTI/BB65R2DqCplfnTeYFKj5tTaZp9HXfcJZRhqbr24OpDEYfiJgJWus90n+SQQq
C+IHQ590PKWc+uToEdtSsuYBnF3ozgroDAS4unqcsBfFCIATn4qLrKPGSRYy3Lzy
3e6ttn13QHDUfO+g21RGShNbYjxaZRRkyoNVpUlfIJ4IatbhLzOWLRjGI1ERrv4U
OOiAh1LAglm31VJWYlIvunJ5ox5OC31ho1ik734qsrcNg2ovUQj6W9MKnpb3dEa3
wFQS9oU9LfQzjVKpLLbZRN8Ei29/Ouzh6V8Q356W5SJPYyslzrD4hPlWkw2zokVe
SYypKXVJriHgdHJHCegEZ6lXtPoWfMsZQMSEGBOHK7SmjWH2OHeHQilPVzFScpIP
Xb3+wIhTBUUFPXZKTU0yW7WqSrfGU5ONC0YJ7Ggb5W7U4xPDImptv/iuiEdJp1Ny
EoCkcLYA0h/DA7twlIGA9ZkrVFaQzdtQTDmfCGUFM43C0fJNZbRBVjex/XqqYNou
9R2gBGqszkjs6FucNgNPmfXyYIajulMEINlLqWVOeVC1ZWP6d6bpv8aIPW4OvfnU
rLE0DLHo/Qxz+CCMPuXEf1uiHiLLv+vc+/QFra87B542w2RO2QOVN+KZFAVKfwZR
4QzEiDsgdQW+jlPBlxz2+zcMSTRnsxGqu1o1H9KRPJIIwa41pSRnNzclE8wcFdxN
eliCDvFfp0qHtgW6Ftpj4Oxq2JmK4uuhZ7bi/EF3BzSDwz/wdQ7eR8YQJuUxL2xV
GPVz/S8kXs77GT7gZmjeXNpUpU62e1pyBu0lM5HkEoJma1tCdVYXTLarzcmUWEYk
fOdUPKJIXifm6KEe9sas76UpVfHUD4sqYVtp1Fzx2DEm6nwLegTndD3i4ACQjNGk
S5jEiW18UaiFRH67SR9hVbeR18dmVCWjcKNm2RWNsmniGgYvL3ZOroabdcBfnGYJ
khFojK1kfsbGHIFJ0RP+hVSAY5pxVjh+e5/4a+IMBIxlLkqiXEyVfilD3s8qG0GE
AtUeVi6fY6IFV0ZqqyoCaIMCB248lZ/rv9N1W1RcThPgacA0Axdf1SI5Dcfk/crV
GN6G/lhTaFGUzQZUo/nYQiW18PDolXeXHE/AYaLoAAuRWqNUldzjDyrmBQxcIrL4
tfLYGBbHz0+6aZKP9lTPLkPyahRjlgV6yC2eFNGrsViRf1tH2MVMVDagfrIBdN/T
ujTQHkG77XhEUQc8ienVrToCnti7IJ8bIndmVoV3qW2+SlykVXclR43fpr2IMzLw
Rc7bhy0+Vh9kemlId6laIWTYhHdSwWD9/XAttNHbD0i/wKlOWRxfEmiEpiVIxbsY
7M3fpnU1PmzH9yecxzYsWB9cAxna7UV5SYYATniHgKSN5YDlg6E1pHf+NzDsE5rP
J79GGB78VOhLUi59LgQxI6ZkXU2IFODm9hYjK3b5x4/yydLA3lsHXLnaKwiSR1t7
1V//S4RtXyb1EU31IiFs+FAw8ftGhXTGww+X+K+8X/Iywwsb2F3gMsRE/+fB+yg1
7XopcgYbx8frzMt29NNDZhn4Mrj1ImCt2QnP2U0Z2hgCcqwZ2Oh8umrkrR8L/cy3
6QV3/hOuHjoC1dyhHBU3hHMxRmtAa7s7VAOeluZu1Vxr/4QJOXtooK+Dj9wg+AYE
IbkdFgP2GeyCFgr75xpOEECOXRSzsioiokQwtIZcXK7Onw6eVilRzK2I0v0bE5PE
wZhJP5oQER7bQRT8XXBELwT9k+BUrISq7zH5j42DWh3TCxv3PE+7e5TDbzFqsTbt
0GDgXYRf9d0B2VThoL/NPNMMa2SZbl9o8CdkmoA9GDdNKd/CYPd9AaNPhBQmtepf
ZH/7F6wuDoLitPknXTtHkbJxhIDssOz7Fa+fv0d6P7Sm4iPi2V8yS9fF2OK5lOAn
hcGFd/60iIfoqGI86yu1lZUS+2PLM2ZMTBgoY2SDJ5gqo9U97dCDjcZI+3vxKqjY
fkXO86lHn8Ge8QA0191Gbu0Id883OqRMPRfkcSSnmXIUtpo5tjsoDkC3ZEM/ilOu
6UetPbbxaCC206GY7FjbFA6nVBPw35XoEPK/XlqUgcKixeaplbVbhrrn/39K7lTx
pbxyo6qcAxqbzFWTIpkcRCn1442x00KN8U1xNrjd6Rc/JNbgr95EpW5zNFum2M4X
JoWaiYgQ+HJziHWohZYlcTWfEDJpPCQCiCInfMclaeO1pe0KXwPwnf44EzMNe9ET
WOncr6ixDOpJVYxzAHrxAqWzoO8ejnY778s90DRIZU4M2g9Dd+ySMw2xxsvo5xye
iW9lUVqJfbVxQTmEyUms33zAmkaJRxZUl25Lydd+ZHDNOdZsPUhj9Ng+aKydPp+b
zZqf0eK4ix66UiY6xLZMggsNqVVvug9YV+wK0/xsRnINx1nNWjSgfdQ5bBjod77/
x1YDBVGHgOpIpWXRK1WmidQkhJ1xS8dQ9f7fSXXyROhUokZERj5N5bxHLSo7rtFq
OvdFsa7XjKHQcyqv9QEwJr6p0XxLUJv3+iIRysgV88ryQe2ENXqRVSGB+skqy2lb
d47RvKes+wkpxw2+WjqnBy5xBwDvpMct9QanomV+bykwB9dzNcryhFDG4m6cduO3
NoGIBME7eV55zfI9uqtodyL7PIr00eKSj0L7jKkmqnj4oj55/UkHwwIPjnEhZUdv
UApRyBt1KYnOjvrXgruCPUyNTq1TncrAKH1mfZu5Wp3pwP2qJE1pvzw59UgSOdny
41LLkIDS1EWfKa1XFTdDBfMkfa5rqN2N0+/ii2sXKipPceMXdmNuMpitFikbHtuC
9zv5kZsBeqvCtVEHthN95/nxGogdFWGgoqjXrkr4Q69NTcL0th7fGPrTEOGQxOcb
Cl0b/j1tKBpP1ZCM49XMKYOYEllHa5ovxhTZ+PLf3whCdDeGAHf2kOxrdzgVTpFe
wQDHSWlleRT1J1QcnD0x52meo3s/frEaMw1WiVIWrruQ9GajJmM0HrUCZYmHyJdj
lOnQ+y2zBROteqGWpJPr0rnlCdq31VQ4xTw9sLVTdNVaIjcnHcojbalqLmBzoSjm
jHkLKpD4aw9NxFNRQvw5a02egEOz36HR5SJgTQu4qQTrSy1MhsLGFXdAS0z1uyKz
gkKhYS7Inn+X3h7s1DwUu/fMkmD6PQKnXIq8Jh/NdhubOcjQtEc2b5PoysQ6UTDJ
lckrlUnuw82NGvUamFFaoG2IQkdeT6ZE+IS9SHwlXnlO8/bvwIMo+oNm1yqMTIf9
KXRT6hUoY7G6629R4YH+3hXy2FXpiaTW4x9pFDx5sYue9PtwAB7R8i9A0aNVGg5W
FTnE74MNJL+ZcmmkYcZOAGvFC0f70onzYjG808o74u/5SWnMyQ//HET4N5WPD6pm
dqxP5X1HZoLnX6SlWtYgjwCfiDWvDPq4nP4ABmqsfSPFLaRsG6OQ5WbVyla6ryCZ
/ZCdZeFQWYYeYjB2JoIvllAcMG7lJgUenF6nr9qdbRw9UgB/zL6A96Or6Lvtpuk6
3k5RSa3QrMc5ydT00yziIkeZIs13atTTpjtVvNWlKfJrASXe9AkftrcF1CkJpQ8h
rJ/6RCsGzxKrseOe72om1zclxEOWTxavZGuJVUcCnzbQ3CGDB+mnJwQU1HYy6Bbc
Ev3GL9QyCajB69modmGfwvRlk3Z0qXwZM0B7lS/Odmu6TkcNRVpZrJn9wT7EXgdq
sjEopYpTUZqukiozLyAdzDL7P2+soV5H3ZCNQCkfQyiFfrC55FuGNuVCiWXqai3T
1UVtit3oqnfEe/hloTADatrtRDDVciPfzDKMr6eJECFaEx4xp00mENzbOxkBSvod
+Ad/U64jpWNLXPCaDlJF1mPqabuxvq78LUZArytylz9+s1DKN4/0iXzSSK9PaEAg
lAU9+m7sNLsm+e/QFNZ9KONkFa1hlhyLILw/gXaoVQIwPeksj2cPaunfMsLlE9+Q
2O+uK/ctUmmkox0mep/W5c8CNqFrkvnwUV8s0RrmSzIQHVFij3r1ldSnQvqAcVHc
b4a/GKEGDpvhxDwIZB9jNBqxqnJoC6rjrd7noOF9sMxT5ZyVCHL/SUWt7o9ubkKa
9fe6sa3/Ec+lppLeoSjlihVxhfswQxYxJPfSfbCxlr//tFeF6lSpRD+hmBqQ4kUU
dQKOzoGOqeTj4Dk6K0HFEUgTN7cqqL0Z5ia6SDWisCFeXB0xrbMC/pzYzOtKh4dd
VdyAQA22OugIYjhR71HgGeSe/doYS+5l4ZjP00ksAuwigOZhKJ5vt1XrVxUnq+Eo
ipVC3ctVta0b1aZX7aWjsPkwNFNw+XBpkaCcz9SPATG3nmaLyYaEf4rIhY8P7Cbu
XqWcFu6NBS4ie0zNcO9Q2G2w5GJgzV8y6G6yiP1/vR89STZ6NgJo454r0FYH925h
Jv90qfHw0yN9IUIEM3U2NQM2aVn4FdrJnioTF9fyH1B81as8rhHVlb5RQfSRmL1C
anaNL7+QnQn6ziDwf6uUQoBlpzMeNmejwJ9RmY1BOe4enmL62oHjErGStee3iXc2
KuDIWTkZx8NPXVNisi2y3kCWV0FcvGIzS8LrvREuunRS1EuMnXogyBqMBaPUQGSJ
f1/P1bELZAnOTiWyZVLeAHm5HcPB+r+aqvGfiy39eGeDGGfnFVNMsnnpY/16m5Qw
XiBTRTLy+t1fUdWdYuPp9ZQabN94W4BCKOKIyrWUgk+Y+s3MVL2VQctOEUiMq6Ip
X5ApY8PLVloisUqTVm6rRH/Y7ConOhj9QU1G53hemDQektXKAhmlaTegkFtFRHnf
+73rWUmMNpN4pzZSiH0mc+Qyq25kc1IOkn/wP9qZNd6J5Nm/vsVg+flTWUS4o4z6
kbedmzlHQ1hNGUlwHRaFsX9NQBqJ2afQFPmTek5UFJTahpkxReim8wWQ/23BQndS
EKXqMdX0PCmVgRw5Yh4qtW6uecU7mXS5ZhUPMG+jPEw9C9YAPg3L74daGDcfUBpm
IYsM4zl6O5+A/v+9GmGjUg6fnbJ4ICIhOuoYIgY1VUZpAzQhtnGQcDT6p4mGdzr5
kj2atydfBSaNC/4QVHIl4UFo/PXNe77q9HCcgzauCWPV8T41IGgeUhIN4VVUDEFZ
w6cmWrOB2l79AH4Y2/MkfLvFhQIv0ugzPgMhTwkEi/7mqUf4FM6BQt8HLQZSbvcz
yM2DlxpNSVyW7o1SzfYZuYtnS3Sp8rakPQASl8IXPTAE3+vEOA8I9mwUyuOFJOJp
MrbbA9nXr4L931ajQTYSHa1SyhkQT0SW8bYo85JL0cZqK4S+EHSX2tMZAPkNht9D
NiH9NG/jR4DscryIIKFKLYkx7TCG+B6377yZf7iUKrPp2U9gIg3udNhTOCIMew3i
rqFcjkhaFXtCva7h723/aZzvHOxL89xQIfuRrenR8CX7BR1LEo50iVUZQNbYWO6x
qYt1RQsk2WiQYcaAuqURoPFFSUX3JhNoKXKDxT0vWbJT1B1Ii/NDUNevCfHnTiyb
wKPH0XKPhxtxHrzGjqIlZwOcVd1NF2otjkyPZOEdSqJEkf/tyyDdvOxnOQmAusDJ
JWNpuPKKWt8XZaRAtchxnh/xVAV/eN8MwvxxQTodLWjRiTkZ6KcNnPgTe4h6K0Wa
mtiNuQa6/A4NAx7VEloVjio2wzcUOYpyoM0Zlu2W+1ne8AILoqck8B2LD7kI9Y7R
JCVbWV8/th/yw+A0OPrnIKt4ZAdnu3KZjUGTMIdoMisjDvqT4V7G0JSKPJKzzvvW
AdUvLkHgLhAJ7fziCkknkrHgAhfFr/zcFLFoUTmqVFheHr56KkB0yBItiil0fE9T
0G5chdRP5URIvX8HXAC3x1uuetv18E30oCVC2Ymc+hpv/ako+J+WxNwoMJoE8Q1i
UCYqwxlYv+itgXHcGiinAySIt/OIzWwbU4Xf+J8SFeNYMkIMjoter+XDJFpXufgn
exsOHh20dYTJYJiwYuWCI7/9CzalATITE6+Dj3f3redspUuHAvbRv1/mVzdCKDo0
zxoE9VtTBtd+v/FQ60XWcaqfsBOgjCqg+rMAdJgJ4kVLvyZmkL9QbWoJ1/ygEbgG
JFe1FCEEV6PHaK794KejCjQg50HNj4lMfsSCBesCrars8RdNHJRkIzIeQ8ROEame
FKYbP+1l7aDc1t7/nM8L5oYLQ9VLJPWe47bZhqIcwdXK5ZB7UiyNzVG4I9NOR/nl
ZwxOmV5G1WVOFfdJDY1vUKvwUM7Fsz3HGfWiy26RCSSxytQ7ktKbhX9/4cp7lvhu
xNqv0u/x+Xk0XnOLzSRWtWHLj5vlX17o6a0csZdiqpBeSLM9MlQpTuqWXDjjKFGr
gNSDfP+PWgo0UB4/5yL7UdYAzt4TrilOrVvkxlEYiVV2d0+xUDm8ack+rM8c4GmU
6wYQuFCYgfKCLuuOg3t4P7jKNm0YYvllOpNr7gVo+SE1EpMFY5fJfJl+c7ybQv+2
nKzGve+PSXjBY9fbvp99n4/+SJOLArSZCRUFlQ5hQK5zrvvLuJV/hFTtf+CfE4EG
JbPn/SENHfDlPigBR+OaW1yTXpaweXmleDMqBebOujaQC512nPQDxQBqlet/I0FZ
URZG45ii82vwi+DbQVbvogEdeq83b+0bo/F8q+UbIWsQM69ousUtkOwJrWPa5C1v
ntyCXLX7y2skKlY4QszuIEcUb+iKFp3cCKOkYCZnVFMbJulSlgO/YvtTCBHhy1US
ZRdxCfuEwI46De+C9ls3mZ2e9HqRWXUXN09ejrS0+RkmPhsHjmc1KFFpcQGlEoGb
gY7s39HYBHVMKBK2Kk6MtLg2C9gx3/mwtrGFAS8kkvJtlX3NaKTOZ7DWSC57kZVd
qykLKs6/ickGN5Gt1YhJhezSWNSDfPDPw0NxGW95qn4+aTZQwuDSXFamysQc2tR3
ekhqL5US9SKtMHy6WIwImgbOUcaAiPhCKipseEDodSFxmnPPc3LZf3hENGsVYCsk
iubU8hd8hPtnSz3ZDlL00r3ofOlqu4xpDlULKnFJ4p1MuLXRb+TPe7pfEhu13M3h
T6lUd+3ngDZduAaKbzShMC4BasRP4GzKx0pFVj5g/pyyWYDNtraZnw3QKBXwrRdD
30D6gr933jXngH7ZnOrocnp6srLqXaj4ejm511A/GNLmDzTivXYCP3cnb0Npfy2q
QfQweBwRgPdnPcw0cKTQvuRejW5C9Or7TX3UxystM/WtbtNkMqIk1i1zF/m4qXbt
3JzZNI/cBXuZgua2nbcMTfQvBWw2B1vxYnXtxcAw30PB1kZ1ZYeRUbz1fg1w90Gw
uRcxEJHwhzXTW2x4BeHvlxaeXtw9jl1bbQu8HU1JTllhGqbtcy3+fdsEk046JxG3
ya7raTyaxLUkq8UAd18P6EFwV6WQud5cLwYc2UrtlBYEKQSSfvS/E73UuzzP1oK7
0Z7TOyMei2JM2ZnuTgJSpBvKVTz8Ms4FSCNv6uGBirX+Rj0GxRCO481OLsGNanBy
TIEAhHQ1ZubZddI/cNW424tRNZiRRT/8ITyb5PJyWl96HESE0V9owcvqBk+7eVd3
rs3oIzvX/piBUGy4//6EXxmKUD9hVUUXJOt7PsxJoGkKSTMYXOvko9k/BUht6VSf
K1ZxMYjEq1X/Ku+5guGkSdoVLqOxzmL9Q4yXJkpgKn30c6ScfePP9xSMzkB9jmyD
9N7u/zMCmruQQBCVgjYzW6EcMEP8ONhUVA+AC5t2iM0kAsRgbpL8oHh+BUbLtwTj
9lPe0l3erIEpcb8zkoPfWHXjEgYKeM3Vioynm5KrHZptLGsw4CNmyx9JHAY7YSm8
d6urSqkLTjU5+rDXk9bnb3Kl+bM7lJedA2c7Bt55sDcuSxkEi20rbkO0/p6NYtxp
Jf0fKaoJNOWR5dXja2YYfzSwTFrsdjAkw4Ihap4xEyTH7q5Zaq0cYMH4JwwLjtlk
Iz9SOm5P5wK4jk1jAC0w6GMrMXrBuLTb5dOUEy2IYaXvN0hRVat2zeQ3fnTXB13u
TqBsf5ene3kG6HuuHADjwwEwt7GHv2rv5sv/xvVRpF/xH+St4GTaVX7aWrXS2Bd9
MiKaBwNbKRmxO4nIRPOu+3T0Lpz1WII4yWqi7wf8s9Bbbrw5l6W96O5JbnqNuB25
0h6hyvisr4mAJtORpLPNHAAu+gHQeCmX4yg+rDTb152AoY+/W7COUWrLqojBdwRO
/wZBSGN/JSZhQMUeok3aMduUAROWIvVEl5dkL8Dgyu7fKtGXhq2QAZs0kehlInum
tBdgscLRBthp4xyN4AOw6VzWNbzTmrAU7Z/4ePjDkDDOtGTnE7+my6mv9hK2sdY4
FMsdiJncXeduH8DQfdrP/yRCh51wVglRozYFMx8kknjoBbRwIsKZmgx2f+VAXdSL
AXNO6RIY1tnMT7dv06Tdx3pc+eny/2QjhiOFwBDucY+nWHm1ImYB8a6YzbWZZQXY
GgKehEbJU84OpEHZSz3Y/OeUgkRHXkeHSWd1xqktM+fL2W4u7KkaQKxjuC4UC27g
szX5l2YuROiXhnr5QfaC8bJp8AmxrNu4KsX5cyJlZCwRTSnhfwoadPAlYbtOFpoZ
WGmYMKXksV9Rfl8t0eEFbWtWtn+WRHV5KsirqHXOxXkycC8HyW/Ql5mjx7UEG38H
uK27Yj8EJjZnttr54F9CKzGse54k8GF/7Y729uwBpugJj2CMphiZ2hOmXmvXa49E
z+3prXDKRnotK6QsOKNbMDachvuBEdjZ5buhdBfyy/VdPqK2DEpB+P8lDXSjY6RT
Knjz+CTDUsmX2OEL94pAkfeDSS69Da+TWwtLnQF4+Kz3b8JjezG9qNUePP61caU8
i9Lz4bubyKFsNwh89IQRLg41mBzrBNNTftbQLAVM8uZYvnt0NixW9wCzRjljQmav
1RQXYn0j6UOvEzG/Qf3LEAdh5QNmTY3jFsOljSrKzCIHda8lPG9CaLRd3+ncbnRe
WGwC7rkWKZHFP/HeTJbQ5l12RB2mfAS8ifZ1Q/ayUr33HB8oBW9+NVufsIVhJC0L
v4Pxx+KhejuMmVXUmkqHUiVyO/UeNjjYIMR3hERXFT4iIL4xueePqic+INFCYZpk
H2aVA66BCqV3kQncCF7NGUSknLW2MtYCIJnj1/xrW1f2wRYei2TiamU5L2sqEN41
Y9t/KsNP6vgazThiZGC8U2X951b/hjk+rS1qNaLf8rulnQXGvk+PSJ4rBOjc2BGn
gdQwVfuDkF/G9lqLArpQWVswtk9iZi4u12aCyfOYgiWRxHMpZn8MyGb18WFx62zl
0opUWRaFLVM+QdPAKsCHN5iJADYCyp7LTeWc4Pyq6k9STA5YQf8EUjj5hB477fIO
7s/9xyEkSr7+gRsRRM6Yi57efH1WdVX6eySerSDgCO1Iqeo966XwlK7KZx+V8BQq
cS3cGpdaPHV5EiqMxNQSmFccIZmtMnQRlp71NBbRVt9qNg3TFdIFy9g/NVKrVNP6
WpEGecA3w2pbCWuaFVWkro/A+iMITR8b3ZQwjdLlROUBlK8WJfAQB3fhdEmn8jeA
nuFLz3x7L8Hpwk6akjL/2E955k25WQzDhpDySIKr1NztTd7tewPXygiVFW6xu4cV
2cKSXgnYpzZb+L+/k5p58X8Z98R5rTWHGDuPdoxT8kW8K/2vt+nGWu5x+rAopGTD
hGSdlGf4XoMzjoJx3gB6ASh6DMpAmpwKjGJCDr/BDLiGxf2do5jLaD51Hvc9621D
TwWFggoJ5s5KKoxPKrGBy32lr71L+IDHQvv1RSFIU0gRdZHcPyKQ4lziITvgaiPx
BeCWPgNZQ/yBiDtDw8Y8yEZbXhtmoWsKMvf2Vy9w3WJB4FzKr0yVaZHV/Xd4FOFT
ZBd9EQzwicqUXkB2i8WxfXpSIBIkA2rcbURl0ckYFrHCDaxe6qb6V118GN22jVE+
FmcVtTiVMgA5QMf+AIlHkTXl8aFlrlrUMglsudwcce98ngkzpiqKKxrrDVs8K+Bb
vMz1RA+nfOXO30FvRQn0oijGFXZt1CXFGvMfgKb09ZuopkvJCH+1pVuiuMvr4/0u
kcNFOxkPaVKGDq7qw514k4YllreoPU8jBxLFOC3PMQZbIqcBpGrjgm4O0adJHsfv
SgC5MK30MAScdZuYXD11rx8EHUNJRZI/AOEqgxr+HoTrkIko4kXUm42KbOQBODdP
rlz8KJEYnYNsnzxZLZKKnYQjuIYDwtZiQynBy1fhvOrX/wayXqOj7OghbleKTpD1
9IMazQA0QdiM3fWk8jNFGe4D5HlZBvdr56KBtekp5GrTyRCEYvHSvh2rbk3rqNkA
l/hRwvGC8yxwxWUQHXs3KEua9fXEaErz04VsAqQkI9dTfxfFiBAGRfxXZt+1/Rl4
jow1LJQORPU1EiR9t4g1dtqUhr9PXpwxHwEs015zaUhO5lE56UUvnmbaBrX8peRd
4GMSO/Sz6+3/5oA3ERjNRUMXpI4snon7H3VEobczZxrRw1wV7dNlhLpLeizFGq9F
mRgqfm8sx1hjy4zbcPHBV239n5MpKQnv5rft9YS+XK4REt7c4KTIGirZsKGLEnNr
MwqknGIwPWWpeK7A+JGF9ygFL1tzaCTbMtpo5wFG7ywf39kQwVKozzYYDs1D20bQ
DBDxc5yHaTMuzFmh7RvrQFDyd+vH3TEnmRzvNYtiTs22DDDbAiXvocZ2hIO73eB0
3R/DrlnovL3vx6qSZQCD0gVH1cF1YNC+sRyeX2qLyIIM7LWxbi+6y9IJBPuK0LsD
s0T+Ev9bQMpqny0N5NUgSh6Mal0Y1/4n2LD70TxeXrQYaJYjHuRULNBfZRmGaiSJ
IoVN3YorknBdiGYQqkvmwtP2gzXBUgp6okR3WkwgGFwTMY+qzWJuPoaBTEkYi/+Y
8flYPQAZkoRbRkqJjVh7XAN/4o2K97Ng6+HXZfdmps045eQ2y1DedFrzQ9waYWmx
OsQMTT/FGI9Z9ArCpk9okZv6YGL8tu4dH6+aNMbQbcwCouwoGUc3oHi+iNu58WJe
5D+7fw5p8+yGgvisj2IC1lIUob7jq4/dMyw0ZAWYRbnb2dQSKBpKSJyPWZq6PIWU
sYpPsiAd0gUtLKuiZnd7zYiOVk1jNRiSexkihDEy5j7iN7TSXJDr8Eto3dejb/Me
B3/Dz8xHWss34h2HHSY5AoCdlULflkr1zh1RvRKkhPXquFCGo6W7yvoWK8bdKX+e
O1RaU5bf+vEqw0LbWaVH5K8GzRr4j544khMldQUh4ciEznBIJb/Ja1k72PysEjJr
JyH8QWezvUmS5ZMvmevUAxX/et5RYs/aMT1f2mNauDSe6wRswvKlUOBSy+dNYfIS
+LgnUhJrhtZDUunc1tu0IwIdICYoFE6nU8ANo43DWkjU7Dmo54hx4wzw/h7nJ/Ze
3e0k4cUW4/oeZ73CQU/kwjd6i+yCr8q5UQGuYxB+cYZY7RASLaISrJCuJP4J7Ard
lD36NUC6hQlLreG5nT1ooW0S/udT5VBOqaRlTZZoV6Og8/wlD/ZimkBdc3Z+zSZy
yhmI+puEqcFPYyATS3eVX4BwIDjY9LuXYTTjPRFPOtN8A7kkO2SGjb707GVbwpjM
4lRXVFS1f1lSRIHutUXQWxEIIGP0BKEM3IOO49KMxI+zFE6jf9h1i7qNhZ8Knwo3
zwjvXqvQagYVACplgx51cVd8JZhlSztQFL9kAoYiAvjbOW+gEF4c+5s95tVqJknY
69cBx0ksS8etMI+O+z0Q1odorrd2pQ855xghGCWcYx9WCQexSjFu3SyVMz5liFLW
gLe7KbV4ok91QKVBCVo/oFRQH+QhKG34SVNWiME2jZw3TV06VTp85shnyevS5NUM
9zzKzO8DP79cW368VVlhIE4u5YUexZ4yoPd7yiuY8R279V4bRWU9csxA7uN2pOIj
cmOXqXOrEkBj0a0X5Mmc15PiYQXeGd7m32fmynxjnz2vHQja4Fz/MUyhNqfKlFJr
/x4K2IoXWgdwtx2XqnIXwiNdUtt12iKOwU8tTU1X7vml74uc14BshZGdbez2p6fm
NhZhjP5U5MvkEozvoWKKOWIuIHS4JKDa/jVaCpyx9EcZtgeQEGmFbPBNGD/Vfy/W
SFd9LbWuRQP0d4jrnpMjH9sL+Kpb0P69zKVotS3q/e4kiy9vJklOQ6vVkOKduOKa
aV2PN0B4VaS4AF++SEo54GNAOujyyG0LijBRbB440sAnzo/FBbbXQAVxKm1a0AK9
qUUP3TCbaFvpdKjXLrq9pbbEfsgv37KqwPiV/A4K0IseX8aKWHxb8YQHDx8NzxQ7
DRFytFNb/h/KHlQ2ed26ifZPvMnkTc3Teg8TU2s4h5pay3rn2cMsQcho+GIlM1hU
D0JjodKW5e+XmIe6b0WJjdmV8zSwP28+xlZLwsrBqh4lzAOKvacLW5mRU5dgWJuL
pHHDlY8/wr3q5ayPxN+ZP9VJgHRdfSc6EMggFzBLd9KNmH9+A6EsyrfP7D7j2+Vv
EqJPe6//QqHC6tYVOCWlsSGpkSibw2f6RLJQvq/cZ4l/0cArlUZZDKIkc4HilYsq
o0aZVA+TkxLN1AKkUW3mnJzWEQvN6qDSmCIho49iS9PhxfsVM2OFFDKIBYuHWm2I
9L70urC2G5K31j6YR+S+hhInlo9Bno3CRtolDLlR3GNd6QyYGOwgTDyA42NTT7KL
eIG7kwn1JqpF+24HdCXZPzXWkZ2p2IyRttN2jfvRYboJD6oldEOepTosRa8jwHSw
AQcqBvdp6u6/idXvlKthiV3nBNL9SGD2N8N8vTKYDFCAGmKL4tklkwk9xP8RKXvv
Krz/FgTiEyOe8n68xe2wd6hGFNmkhrcRnTQgCDgooLsyOV5Yjr8JjrZGlo9LBUTo
IgaxWnF/ZWX3exx6Tn9F6LdgVWzVDH9hojICHlDtru/T+2Rb+4+QVP8G5FYxapP/
jwnLpn3cDC0x6LrLKMqo1+mXTSfanwpGEx70gTJTjKWoir9j/DROGLWpr+7UGXoE
pmDvY9kEIJH+PN8yUqZpPvg0ESEx9LZfti1XMZplwewWyBQ5GuK39yjs3Rj0Vx5I
jhOKzvDM1AMZjMk/7HD5ettaWgJKqXqOfpkMAW5FxG976GmLkplOcfEHZz3PYWAM
O/EH4goQQuXuuR+IrmxzOPniqPybF1fwdGrSaKCdWADoQKgneWLdnCyDnkjtwps8
l4g7hWqCvoE/wOGqovNpO6bfxrqxguwCNV39PlBslBQHCFjellz+W4VFt4sF4gj9
5lBHkit3483DXjrnrFC94XHyCc90gEVjxyszd6lGaz/zc+BJPb5WjbO9VwYTS1fm
DyLAKlbTHBsvJXMTW090QOEoNd6pw1UQzlGAyU3zr0DvqhNW+YPlnaPP5uW2HOYC
GnReIRkJu40cDRdzVItTh/rxD4/yP7wqxM5aR40zX2OVMBbBBSnEQXthM9kVEzbi
b6BQkAdpdYhp1lYaix/Fq9PePB1/iajUy9l5ZIMSu0OETqHI8v/NyuyCL+zMzkgp
r47iNhvDHTh/sfXyLF1dGC9H1Sjsn+6jXPdkZ2hvEN7CVRNyymwuuClYAFWH4Atz
fICY+ucM7pqkJG1Lcj+wFeKQP85I9R87gO5LkQGvCDKk4Omnp6U7rPTvTF/aDDdO
q0yl4NO+yEQgrO4/3uE2Jgv/S+Nmno5MF4JY8bts28Ex2lNz0Ex5wD1x7Ec3phdi
0CJKSd5uqG7rKYUY/94PRSLIyVe0jwgX8+HQaxH4Q/HPlJ3GxnJQsqDBKWMdcAqx
oEsULNTIBrYXteJ17L6PJ29ShxYbiZynrcKIK2vEhg/NE8fQx8WMHkOeirF8W+GF
8VEpMQucdsmR7Kv2SJWLy+WKVQBdquLoKV2rL+k5SIzcOTRhmQdAHatoWDdnMP4N
whUrWN9sfekuvQ4jpossiN/TrwvZiWghQu+DTHqxbuBVvgXABDkd5dFtG5lz1DIJ
WK7WEr/0HIMF8gQcvtpBUhmkTbO2CX4nCfQiiqD+cuWQFoeAZrHayCP7O1l7buI8
uy0sUTmPETqQqQ++8RgWThdOWokLCJysd1trhnlnAVRYTT1XMDGLBcFekmql3U6U
o5oNRUQggsfP8a7wrhynaGAS2NtV7OGPcH8v6UiK2rOFv+IonnDzRI66sXgjlq4V
NcnW/mHBLwp3tTX5deL1SxVxr6zXdljlDx3cgq+AWH42o1ewtoBdDTqbAkkPbFgn
8x7viiUiCKOuAaSyUjgANjkBFDBtYJLb3owU8a91Vfsr1DAZSvXNjMYa8dj8gj/J
OgXFOOkReJB9vKW+PNjE5CNVwpYOasBr0DPJf1+l9pn21NiICqjt71mIICFSa5q4
gr5XJpAen/5lFOV9rK5BPbNfHuDr1XT1joNNQSoIi+n3GuYOpbRsQkVOmn8ke1EN
G6GFXoZxR3P+qIGSJUg2OxY+HNqoZA0O4ihx64sxcsalZvQSga8LuXakv5T6RLcB
mdyEOr9GyMHFeyCwbzNt34HRZH7u+A7XlJ2eu9lftUO0e3vtlakoyyaLrf1fZ+hS
3ct0dL8KQkbd817vWL1wG6gjUOmEksRJP+ETmuRbyqeWk+k5X+tuUx0MUnpcpzxC
KX+nNH0DTB/61TamP+lrzCYEzL/jGqvXW0zdNyuQw5XU0D6T0JSLpJGw/MoqQzZO
BZeLMnNJRMDsghhqeqLehaGngGwbMhq2q9qO2W9XdObUrHXsH1SHN77jpt+K474u
ouZvjyst8jPr8gWhR5gMGagOc24W1m77RxGHm2AyS6CGUU/RjeiQ6CQLahMPULyH
ziAXtYlGZnddwtpoEVDrW+8E3me5TCieRYZzSPYTtL5nnAGZHTP6XmvXgn+doDTN
s9bMu38LJNmO4S8O5zMdJxlXtggCcfA6wNL7mqNp3J6k9HrvqJ9m0hJ5s1Dhf571
wCzExWUOZQEVv/r9cYrihkJlm9elbeZZaQ+YB1AiZ3EF1UwVFJwc/42BPaZ8Oc8y
K0z3FusmA11C0fKdfxUTpDjrkDV4/MzbEX6vAsZ0a5nxmOpbpbqZ6r7mZZCbQ4MU
UBx20KrtzNqMwzdvVJ++VePyFTPu4iS/p0l9CY94NQyzeEu2FfgsGizm9neKflz2
t082CC8MY0iRZYasg5TddPByqdHhLOUi+zwVvQAW65stcbdB5R3KcR4UoT9tuh2H
TCmy9xRaZ1a2yaHiYxEBnQmjAgUdM8j0KTasJotuLNDf2qsjDh4izmUWQgh6Bn0j
lJv2re9iFb1uhvdY9BBkeGfYLPgINcaSQvKwIPHUk9JtI30QxMVSzmd7pRTCtDCs
ACSrsnSHuJsewNBocC400jadf7Rt6PZYPirHuulyN22Q7LHoEfEwQ0NrjxDsG2mJ
BR8WS4bM7RuA2WfGBm4gNiLdKdd6UJ6Fe2+pxvQFaAYUV8Pig933APHNej2fPjOw
ck5BYQkqvA/O66jSzL/8poM40L/W2G7pgxjtl+Zp5owwloxJrcgf44VLHnxpw2kD
Teh21jj3pj+xw0yHVvPgbmqg/odk9n1zBBmGNtD1qHSrycjiKUgRqB22H6a7xRWL
odgvGxW0wXiIWYo0s564dK5CRM2qNpEyZMv4ZK3WwdlulbJr2TGNjl4epsG617Ib
Cy3BSS5+8/gJnEHO9g3ifom17qRBvGookoTPcHqBVX0YAK0G+jopldKTloJpcrRR
ED4o9xyTkcSGRd5KQa/0fydDVredFLUtq615oxkevYtpRlMfQlCTmGvrZSujrYJO
189RRjMc++3LNUh4ateH24GsxdQDlH0phUC0p2+5Tm8zQCKk5AHM68Xae+nX6nv2
99KZiyCuH/FR/zlfMlvDLFRl3H5Yyv0apy8PMTY6wAijdMXJPDmCjcgKsJObXR+Z
Pv+wokcvwUYixiQ8EuqIx/Gxwg+49ZUsT25bGphiRjMMe1GOJFMnOlOPF6Pe0hgT
gs7+Idk36gBFoOeiHB3kmOJa4mRj+WG5OHY2aMzDJkRGlWCSmMDZllDvJHvbGBAv
Gwa6Rl/Qegxmt806gpAc6KUdVhOpTPdA0eL4332yTgyUh5gO5/VCYT716KAe03wG
PDdIf3vO4jzOONwfjfdwzurvvbRt0aGTS3+3kU3BwMaOCejwOF4Ztd/nu0aPW3ab
kW3HJne/jhQKEq9EkrsP22GSKN7US2YYRZGu3uaK8TuqEKHggFufzzk1QrCezDhb
phdfhq97ix0A1lwjQpUZmDgfe9qxVzxNG8LGS+1lz9LWy1gZyb4jY+U/2IDS6CtI
jhX5enQnUV9wKhamtdrktL0s9B330P6T3J+v7r+G05Yt+aT9/SXjxJEYMsJ08zaC
KU422tThYAK6Qe5xN/E61b9QBuoVWNeLjrjN7ER/QdepBWYbTwLfm4L8aFfXsNVU
OF86OAR3McPlvgOw572xuDQnFfIBmve9vepJoEbyqo06Zs/Zqmnb/qRzr+ijwNtc
AME/ZP96zZ3oiPnFCiIVtXNkj32GhV9ZgaMnZOzvlinc5mgHCgwRqYMU180flPGb
X7WfAIIwkEaJjc3sVnqlwqSlDFdKV3bHMT0q2k0x3vlqI9J+u2M9LoXUd9iUODkb
i2bOFlThvpPXCkJvF6ZRzH5++xNrup/34a3WvETjlpygpfxLnKI6w3ed6wXDJQyp
s4Cg8JwrMtmeKGCZnTyHGR8JVbBv2SDN9wGUKmPlD4PUCyvSWHGYAIbAeN0Y2fpy
W63RUWZpjP4rxG7Pbs4ikRrl+c458aUvrFaqJKbLpNRcrWKooywIdlsmDRwGgCXR
Q8MpqA8NfcSvytjTNfD0BYvsqhauUPY+4vrlxoWHPNBo+Gn3EHsfWqoZ/yMUg3BG
2etuqjoJm6MMld+g0vRnGeMxz3DwFD93v2euNEyxxvGfI8HWKFaModJwUJ98knvT
X0GcituKYIdbLpAI+37l9i0eUlmGOT3Ov2oF5RB9rtp1Xa6P8OiLfyKRdZg6nOIA
Ps4T27k5xQurYkCKrxaemEkBmyaG3a4rHJI4puOK4JdRNOCuchwLz3ZMivFCsTpo
GWbdgFV+pVg1LOUMspF3tcoMVmypUPC8xpkM/Tk6EAngLy0GJ3yphgKeCf2G+5PK
A3702I8I6X6HDLPse9Pc2kIUqIb++Zp3oQHMJ3tiSFpyXyd4PutaPDxp41zmTq68
E9WvVpWtT4+YT+qOJjGAm3KPF5NG2CUgZKkVmal2O7wWzZc+hiUmCKBUaNjeoUiw
hHnVO0siwS1j78C1ELUSOt7eCq0goxYJtxfWuYwRq2wELpCT++5+SGSqd+kS0z94
4wy7ldgHyHFKd9xXaBTH7xh6sjEm69lnWXOnTV6CF4azMxrSEQEjEDiGUWp/3BJ3
TPzevN4JBFoICmi13O2QJWw1+aqt/MUKiokVf6cGQooHBb+o5F4xit0dyoZ44H76
G0oiaP4ohvr8Zo9avW7X/raay4HGWDUzTGzgbXWy/hNP0h3dROQwLUyIHrahpEpB
ryiLP2ZmpVjt+tiPsOhTEpvC1gEU4jqkmgpohmkGpe6L9lpJhbtjCO/SKicax7pn
wBml+OCM68EW+sGa2jTWL6I3xKxCn6h5cEqFBiMvMm754yzXEChunJ3UQzWObitl
IBpvI9PmCax95nT1fIBuArYoZuDLa/uGfBHBySCNz2FIowiS0lm4Wf6z+TsFjZi0
4eI9Gdfs9ELvWAyqlQXtP6FNfKAQejIw5QkOXhUh8KPm7G+5qXFQkr7jTWjgijJs
urkTUbpLnsC9nmGYCwgrGtVc6xKX07+OgQ+egHVt8j0pXG86eioLmodjdt6Dr+SH
uY2lryp72LS7SYQ6KF8mG1hXK7iJs21Q6QvN4K4DeD0C08ixggFJwxctWMSm7yie
3eHlo6DgVHWiNVjgVuR06wPy7J7n5rEk4yd/o1VhpmPKFHxHMGEKVGl+KZPprSOG
wPOzuMIYnySpjuTI4qwedAOjNGW1LOJn4z+7bQoXw02ZhOANvk//W9ivRsH8PpXc
EqZc4F9SJrVUwVnkMQF3G8Jr3yGAl34lquPBx9lZkOu5Z+odZohkR0GFqQxtaR00
M5PEnf/IiOtbG76PSEt4uC9n+BT3iteZpD5ASy2g89uVn8hU07CWSIUnvh5f0quu
JlOm3F0s2D6Q4wRF34wAJdTmGxKyn2VfBZ0pW2AooHREBfLk7qU7wKTvlM14Hz4U
Yza/ABfDhqy4Sh6L1OGue3Hducy3SA0FbAi+PuJ7XuoksKirtWqXYrhFoNRh8q7a
JXCZO6lforzEu465tUYi0Kf7NBUyg8FjYDQ/LEDeMeeMJPFbBHYeWIrxExHd/XAo
A93Bd145ctXs/BmS0IkY75suaNAJ8+M7oyegQzmx5qn2SigqzZOcHzOc21s/IYSj
G/wall6Am9KfSX0ZuZIeDRICmdfs6W6BMZDjKNnCpylMozujoDSVjpiDx60LJ62e
fEt50mNE5ejDIFYq1tJvh+r4m+BBituxCIFHzTfLNTFNq4BWCEEHFfBW+aMGk3wy
UghbSTlhdXGqJknl2SRLivmrlFk360WiR7T4dirD5g80UeNJLBBV3XO9ShBsxo/1
g3QfSdnXx3CCeO2prrfj9xGk9/ChK0kUXSsZ34skY93Iqlev6Xgjp6PGwGpPw67Q
97XRO4d7WRV1Gf2hkFlXPb/E1VygkJZbMiwd6wk0CTXNqrWT+4DybrAgpvfB6o6S
sfGIoMhg84i+f5kZ6/wFKbX0bvtpzSx384PV/0lLjsMzaUg/iHUl63hBSWXir8JE
6NmX5Zt2N/lcjzv37Q+6/20VASN4RRrWURiBnuddeU3PGDuvPcD8z7e/+wfedv3D
ofSe6WZtls0ZUQDR5IaDAHTtfMBr2xRa5+YUBKo4lJIRnP8pHI1MYet2J733Kjgq
iHHIEZZioNlknzLfoOKKSKH5tOI8t5wMVcVW3Ydl/r6PVDFuNakGxJS14LhqOt8r
pRNcxr8E/ic9tw0x58iOa20Twyv+9sEUvV+PSp0dlBzXCCRagO3oWhoS+DDgQY8R
JlmMzx4GunJ4nbYGAEHHiQyZzDJXSPgEfc2lJHtHNwqYj3OztouqhSMFdDDHFZ+v
RbiuPcHes7wi5rKfada3hBz936mTlbE11l8PYBLrMYorTmqf02SvH3OpXRqM3vl1
OjH4ohf1a74XtVZLR//lFJp8aSpW3clkoKeoQ/bhihi3ffcv7tGUA3uUKJHo9tye
dsmg5wjEty0DBPEpFJmFOKaaKKiQlR6fTrxins/xWL4nZ9fDYbQosdjKlIJHFS5q
Vx7kYNDZDq/4xOXTo94ywb4JzTQ8u7i10j2wC8C8wemrLK3dG4a3ENGwMl5oeM5H
pTD5arMUYRu11NT3UBoEBBSWwxUxa1DPieL/U2K2R073Gbgbh49D+GCpa1PelG2J
z0vmgMsRj83kbXWuDpGaxlnOZYYxwc/vIUMrWSFmZGdHIKjj7kzxsRGG7LuBhkSB
VuKTDog2mSSZEzB3rmGGnSE4ToL9qJiUUrL9wmx1dOkAXEUt10T8pVzvWVkTDJqt
OSN39Ag6yizHJ5RTZN4NPsegOpR3GGBk0EUajU/hQhOfDb76GZ9lcjLLunFOZsV3
5y4BYfl4aMEnlcwg9zVRpNm31jw+goV+X/kX3NmA6L8q7E9kckY7uKiRdFkd3Xph
IZUTIhjQ32SLyWvRfyJZuG9FptLn3FZ83kyTpo32UKgJu/ncqMqPqMX6Iw9p8ZMy
0oEJocrQyukNht2NtC60liAneH45dgT1+UI5lGFp+V1IzR0kaLELmchS/Tc/j5NY
nB6u33wAKNgUjFaSH8ViB2gu567tr7ZQL88rK1NNVnoVWcFI7FPtoZ0nFAqjgvzW
Ra1kFqO8bGNY1tfLkwGHLk88w4c3fGtzgvObFxSJk4VoS/V2p4ZFJzNu9emVSI4t
iRkaV5a16cDVfVGczh1xG74p5EEOhuC4fY/O624R2sHXrHfESRh2ZI1ePdjF9Pi8
zIaLzHdb4yxm8HdCCMok8jPjRYoICKZgkKS/7K58ZOZREecfyJFJllZ74jL0dggF
pu25Mp9mudzYAz+IAFW4Wsr373zd6CC4FfohjvrJWV3cJueTcxw1XKXlwakXxHPD
tKwMcDm35Czz2FefaI82QvHuLcc0a3qlZgcak7HU3X8KotQLNjh5eKCBKjP4d6Zl
tfUAMQIkHjyvBu5RtmTH1HI0cxzdFymLdo/BWs5CVzNcRl3koapwtdg7UwHq6cXs
GJnoaAwA2mRpfAXQpVTSU5bfvz2JEKLqdMeMIFqV3TO12ImbwT66snzd64UnMuOJ
8+BtKMOI67Bk3OhrxoZeA7XB4tNfPqCn+XDmMYymiJ3KWSB0ONGRhrhF3U4D10iN
pUnNVlFefFeI+/0en24Bt1RwWhxkXW1j397TOJKb5gzxVVNMCPoi10OPgYaVadJw
PVnYVhwfw6gz+NISYay+uZONxrU+oBqtNvx8CrMUj2TupDsVdTcNYyRrJCoeQjGz
/9HuVPUeckLE5Z93WHbsAjPrnCcq9Ng2lE9ZR4JVVf+SaU2RrcPuq6cDTPNvXWJ5
GOXeamh0/Lpm3B2zHYfu5kq63F0ve4dS2rmq2LutJ2RNbjMHtxQdH5NfoYCmd5HR
PfRGAc+2yJKXjp1HQPhakNYyZMCejkj2YReP8rX3/LbjnjS83dLHCyxfQpK3bru8
88CjB7MAqsr4ftx6Mgze/K3IbLaKYZuXha8Vnr1cS0XRFeB/jlRBolyCj3bCFUz2
ngrVkcyT9TAhknBPDOi/adcA+i36Pdgg2mP5S1pxNo3V6WyzAHvhaHqMscuoxRXd
I8J/onKpFFj89eezQBJG83olsZlO0stiLq/8hmWRAW/AQ572rL419uAWvU23kWlS
vxZzFbCiEYfLvtPVefsD0sOKEjj68sgVF8zpZbmKz9hUgB4nEFq+Fifh23Dx9380
50Vc5NuaY7ZvE2krnv2REv2MEVP5sOJg++alVP/j0Gkbd6Ihua84T17NUeoTtWyn
Gm4P7Nqijsazwy0W/UjGP3LDG9t7epewUyklH6DjfA6+LkmQItEujgQdoQz7vCHy
sEuhCgMkuSQ+OD647cgw7FKwWIhkDzxgtNPcZXPc97SATBoViryBP6rMgveBdaqe
O95P0MeEKZfJJ4BtdT+IUK1pl05UlGLE5iZ8lO/Y178ddoSG8SOsgfUAlBvb97/y
kKRtbnKZ9LhMnZ9uyOCi6M2JgyW7eP4xSW8heeXplAQT5d75nChPDfooIy2fN25c
outGCh+eVe+eQaRhdz8adCc2qwg/bulCQhyPfE1lZAui94a8/O5QbzWCVxUyK+VB
XKZJgxCFv2HxOUl1oOyW1GkL9237XvHben6EKr7N+/GR5otd9hvcrxWc5epN+6mw
0Os78y7dnH1prasu7ZHJef/WyeK/DnNny73z+RHbaYW6uTKQANxoZHB1xYt7VAq5
ARUQf4KzZAvemRXoA/bM4Ep9KKdsLV3Nl2yPKprbAGOnvYhRzt3VqszrEHPpoS3t
XM88F+xR8Wwua0YOxSdwTxqBjCSxr1VEqrtOwqOPihAhdFn4wVrbtJxNGT0oEikZ
Mno21D9H71M8VwqvDWSCssZtJy6j3+N67FQBX0yfe6PFAutqr4siRv+WQu0VUbCq
yT1/2pirCupLsU7/2qfpTqt9DtJhFqMr13ZA4tG/L9HZGoB4vsj+yR0JOAlXO5ec
L5y+8YncUgnt55ZHfXmqA2cBl9NyALmjXrIGBY8PchJNp/O7P2wMGYWO+yRe+igP
5IoorziJsFTThblL1h3E/EXiUWwo+wYJWTbtq3W7woDM1hirGTpRw7u8FR5W2550
dJ9Jtjwz7gCffM5XU82GPdQ+sm7GUc+I60oxyGxeQZQNjdyEEGIwlAHo/fIfc/Qn
CA3m6WlxBMWE1GW938tRH/Sz58mryAUx0VhuhZrsxCDNSD/zIt8GV9Dyju5+9TGc
qKufyHWfIfO/ndQfIwaKycm9HUmGXy5I99PEVmXvIgcXPRKU3QOONrvevaYdeAqp
8OhTOQ6UTlBjBeID2yce6hYQf2R9VZ/qY64tNiE6HbyJDo/P7kiCbuw3ct3eS9pI
GLMtjMTGbODsNBqRSBxp+fclga7xR8UwvpG2uPUTV4avdOKAPiN2DHGSbR0grRD1
nuH2ve77WAbK17LdxGwsiM6HRIZTBx9p4vfiirVZxAAov+M7KgPB46564JZf4z9h
M2xlORAVoUgOqHD/OyVpvQl6oaPxkUmP+vFEpHmLk7a1xesfruQKO9dT12X4HF1J
fW7K++vUGcsvFbNNRNiwIeV0Jz2DUmzHWrl8KDGlLkIw/hc87G9EsKgN45sM+waI
uI16+dEuurBxoC7nhcOfrQVGCHpIiVrD0kORLBbzzpws05p5AysPq+BPTOLohZUR
RW895p/F5DpDUThi2vl7U3XEtH7F9GMnRtcIeUfn3mg4LgBsoHW84KR4xg5nIv7f
Bosd3RcNe5//uESe/ye7KuOQyWuMteFTAZuYXIJLkBhTvfqJtbCsYnOEyjMEX39L
ryHM5EzVew4uNj2/aZ2w77LA2eTobLCIDkyiSi0Cv2iR7uo4ykvNWbu0H28csB2+
fUBQVY2cq2sHQWXS9nH09pQcIdnBRzUtAabh1viVlWsmOmUumECnK+Fp5XKjftab
DeDA3/kJrAF4i8MV4qDqZETcGKmzamOJ/RaZaIu+QKu+TuAyNYTGblAHlidrRCR/
LT62mE0rlagtuHFHKwGuhH4vOqge1UJSYwe9rrIkh0ihccHG0oOfLGW4IbjgiNVk
SUuzdBpFYcE7mzNy+lsFyzrm+6/7hcz/8XgUCQIN1OLwkfUUAg9/foZi9eQaahTn
LBIZxbBl3ePJghEN5fBda7jaRL8wlv6ThXtZblWxeg4IiRHMlPpcaUwuAsbVV8yd
7qnkV5h5eRJ6UPG22jn2aNq6sOfub4JjCHFjP7KFFhh8Vp2CUWh+18K8pljB+Z4z
UIPOpzc+wkSErDJePzwDyFBL+SYyzy3n/DU11g3m0P4C9U22gl8JVBeSkqzos+/H
4oOb+NMur7bYPLD7pxTM90hcPhISJ+g0ZgE2Y6YFLBbDD/uP1BTYLn+31IZc96U0
mXIXI5sPN8N3NeJ5fYvob+AkSWRpYQGKG8f1cCiOR1eBf5ql4JEC1WbvWqXMZsPd
VBHEiWTA+gLBopzLNAf93nUnv/3myTduJs9haOJjlxymI0OLD/VmzeD+jEUzaZwi
dYjCsvbxQCPtF97IiD6HDomOn0F0xyPPECB/xEikXTxw8NhA1OxrObANTK9i2LSg
1mwTukGhSxDwsgUJZ3qDnCef0zKYJF+dwGmv2SOJycS7EVBP8ygVFWZmEaQz/9Gk
3ZmmqS50vzgQoFAb9/IaDngAqVaNfjVq7G+vHnOog4n60A7C/nRzcAmwHl8bjgXb
4kswBqsSss/9U3Ef9Sb+W4o14HhUk9gu+XhaxTIXmR8fLgfUliwkCnE6T/CkPiha
afBGBpDKpqBJSinoSxVjMedKa4QXF4OT3vwkejaar1G51mA8KZhaKQVX8pqYCP07
GaGcDWx1TUpF0YktRZqxWcyKvc5p5RKDAoTBCED4+tViCP3EXuOGOdjp6FFIwl1S
ob++o7krPrc1XWKKgLL37EVqdGxDIlMC2dOKsh+CH0VCrIrJq66wAbthWCRvq9nw
RpiK31cKbiInL34eyaYzx71veCq6A3e8nSD9s/UMjS0Xq7Gew+LIVlRe6EdcYvK2
jGVUV8Jk9nydj1ENjVG/OvQZJepKpPgCg5uPtw+19niLAa6Z6jZNLGpfANQhqIJF
hKr1xyAnG5JGw995WjVpJfLiFOL6FVb++DRHTozbO0KtFrriZyEKrx3v0XUXLYdY
DNAMXtCLTMIGsq8LCWjm14CcDISGTJyo/7fz11LqOAHINP5EwWt+3AHVHJRARRJN
fOdNVEt/9t5Ri7f0ymoB6J7G5oGbtaq/aPLUTL0ymKQADklUc5jSC5i2AEAdK73i
2M8VfpWFlhwx6/SKWA3raKDNoeRojzhQP/tLEdk1qqIvKy0J7es7MGC0Vvhf3hDR
kEjAtDEDeOoXBDDKuxLM08CxqVw5fz8nM2NZUe2GDx9vgUS3Xvm4bmrKnnfFbIiz
XSs2frM7C+qMlOxAABN4wZ8NFKBX8apQuRYFpm6KN/vc8VCiVxza2fqxkEnGiExQ
HfJvhe5BSmYHWbbCFsy8k5GbvUmZLh8/x7V2t8TLuoLBCyBH2Cst/XygxZ/pNLW7
xJXv0qOmRBPa/wTq8Gd6uY3YUwcIfA2f8s2i4DkRUps7H3deqwvIsU3ZB/BxfUjW
9peyE6XysTaiajecLIFgeZS4A9GFsI54GemFrG72G7HkHj5uihDKxzXiJ3tjnwCG
0C+BYepQ8SbolyTZfCtvKVaXf5a6Hb93U7RsZZiwZKczJ8sJ4DHJd1KPZFMnkb4I
45ArtJ5ht1erIJU20zIMaa63+25x3moyu1HAabH/hj2E+/31ovrlJ7ic8ZLMJ1kC
HTLHD7B7E4o5lF3AvvW5GdrIzWUW/sQoAbT7PUY+oo6gb8u6s361usETOOM4J9ed
Jc4CGfwSR5PIX4nY190VeF/xp8taeoenEk+gtisx3UAd+YHl8kHoIO9NR20hvY+F
YHhgokDaIxaYcNGCt84obWBAo0TRGuxEIZEtfiOpbh57vb2CK7KublyMBDTnYtcl
6MfANirnfJo63t8hGwfjiMbsqaLJV1YHfwbps85VzuSwWR0GFMKfrziTFpbiT6qy
qF4Q4qShn194/opLGpfbsvl1GSV02lQyQUqVDsptVXayW3nNmex/L6wJjbgEy7iU
D1B9p7ZJxz0uXszXrPFzopcTPFazVc8x3CuQ7dfFl80y5PQVWJ48s5uTd4ckcnrA
km/A9yuOs7/yRQIbfh5vzNQa5v5jtCFtqIVUvwn7TWFp2OxDWh1vamavGXtiTNpW
3w/WwDXXku9n1ChAwCNdpuEhyavewi7cof8+IP0oA2hDRxZqIct5+z/fTTkiRoMd
7LlhGgk5W39Hp+FQYM01+6iAzyCGICXqLbjfKkHz/u9FKPAb7DExi3QaynfoKJNH
IbcmVRrfytXRTr8fi2BFNgSfvoWQe3aGIbpavyUm2DQt+CVpQvTVSlxKJ2itjpaN
ZEHbmjaWC0nbeY20jNc7lZ0lPnmHogwvF4LPelaSYAb/SnWV1Vngkm6Vttww/Pmk
IasgsQb5A/Yf0r6JQWL1TiIKdDpCtaMvHgHN9AVgPBZyk6aDF7lerrvWfn0RSPJm
ToZJzUQf0EBgguROtZWEvaWUS7Cu7w5bJcvVQgHf3a1CDicUL73wpm9Ma/hNX4ta
ZJhLMUh9tZ3jVyYvwjqlI8fe2qjctopZM4WonsX8zKvZ5e3JfmNg66DQ+/nKdpOi
KgFRyKqFDMzUweCMGOMFthzWSyL9zqnmFECWwNOvZswH/RfHujwpbiWxttBmcebR
TkMs8X2hkkyJUHwmhKSUJahUDQxKgIRjkhY+gzmp2oNOdHYC/1T5WdIRm7khWU0a
EbLg9+8sucbdzkWF5FTuN7nao+GYOp+EmG2BJrfW7Oeu8ddvuEiNnESMjFW6ciXl
EQTfh34TdTZapPXZ6FFlZnW1uP6ceb2HoX6b1nKTT+3Kb2qGU4auMEu86kN/j28n
c+2hU8+DCBVg2y0P9P4WzyIB7TZa+zI4r6Qk3P0TlSqNRZ25Vbqa3n+dtxVwqX3J
NBEpwDRLPYF7wJOUR0eX/aVb6YZUcc+vl4hCbpGrwJjf7IiYXDE2VryMX1PmJCoh
B79M+oo4/ioUTk9pP7fP30Kz8048WQ55Egfpi0ftIbc4x/eJTSF6M0rZuxNOLsRb
NVF6Ec5MSK/lxy2oSY0Yd52VRbqW7sLzf4KBWH+TCGS3cCQOpf5ceSJ92H3PFpLj
5KTY6fpe36945khp8dj1zCGr3ZX6KcUHiOBmAjLZKar9u2sog5t270d9lD+dIxm3
+NnW0g1veNP7TTEDx8ZlPH/L/FmC6Yg8P5ea7kFU7ZGU80wu8nbvr64IJhDbMibc
mV8l5MLIOE7sEgCfJNL3bVd6+YI+xCg9L0dIEn2U91pTPMfoIysZFjOfY9rNx9FS
pGLRaiRrjmBCj9ED1dQfLXRCz2mXqAQLpyFJf6fXJed3Mzft0gaVvcrRWeDALfQh
4FAb1uakzUvMxNDBd5QyixjlRffPEke39ikB9iOujSz3h78KB9/1dwSFaWjmCFLH
CAy07fbAC9R0lMJ/SfXn2hb6IQQSjwslJXXs/Uji9CCN7d0gN0M3b7dSB0jqUOK7
VmGeWyuTnfD2DVbdpFSqZAoq6+GhrXA4Pjf8BSZNnS3QZyxaP/Jh4aVLhmYd53sV
P8oiUkSr53i+cq8hw9QC4UDWzcO0z7RgKDgWhrqtq3br7p7SSFFCMhI4AVO8/5GY
jRTBK3VGNXeYVaFrwAfp7Dz1yVMFcL8IuPVxvZYKKT7+8Vb83Ixxks9x0uTxHqfm
0ltk9PtVBMYJDqx8JM4fqMNohkxQF/ti2XJalEx+zJDuf2MyV9M7Y6cdLlLR+sem
fHuHRiUt2EhFOotxQixWrp879vsI6d4SWIa+BhXRP0bChUppZvuy+bvctuZHsvNG
vGQqe6/yfazlpQQmhp/CbbaiLZxT2nK2j/7U76XS2shReQNA6diTuBVavfqCPCMu
uwmgvSI5CTinZJqYsof4Zsd6FEkCpIzqFnPw6p1C5hX/sZbwauRtWvBsvhOU9y/z
OnxgUxAhS344VbVziQpqUlOMascJujtyCCjl/jATwR/HS/6fNy9UMHMO3MTRMy3u
g25w/mMk/xxqWjZrQNL6N9DYYBGZJ96cZ1X6/mCj9HcTVF3z84Ly/MHJV1Q+icIp
Gkx1/dI+SBOsG4SYMZkVFfeynf/VyIo85yAiuJ4bpDSURZjXIBSpr0/vW6gdUCcn
apsKgAmmmkmCrBnvV9+xjgXl8wU+GENydqClYo95Mwxj8Z+SC92y3rdM9tTunPvJ
u30yP+AlyTP7ERU6F0HmF1h4+4lcb9bnsy8F05M6dlPBrQUXpgqRrF02aPZCpVKR
9HL5ZJY5shIUloPehTxFqE/HqImbNt4Pipgaaw2QVSkx9QShrhvCroCpV8UkFMNE
RK/fPPllRJELxE8cWlkllrASca1ppMmhh/RbzrRu/B0WpWnasS0bHO39Nsrv2+xb
smpUIOT9C0HSX5WXd1W4y81XL/KE72WK2vl7d+uSqQJiWMXdw3JwSS38UxY9r8v9
7ko/PDJCwRVIDIasxI5h/Qo09mR62DnG2IADASYaCr3MjiSLkR36ByeyTGrPo8Fr
aKOzLKSQ4YbMcKnoKMhu6KSVC1u+LdCrLc9sH0y68NY6UPCjYD6ZeI0o0nO+XfH5
zH0H+kTyzm0puSPGv55neA0IfqyUEFAQTXHd3nVvmZCvMkfhRBcqKuNAIIg3+IG7
2O/+AM/0D+76XyZ9r6FmSJOj4B6zgo02JZ/w1S64ea5PItkDA/vQaxBp/dS/EVXC
uwhGxtklACd8713Fw+8CA5cQMsN198NfWAMkTHxQXcS7lbBaYdhHgdiIgtVU+Kz+
nynN8m5WetQf1xqAZ8pDkNn3i6yOLsa9ftszg1Jn0oBdE79uIh4rXMGXO3Uz2x5G
CWBSWG9wjqCxGsCLZB2I9bfBhKATwpXZX1O/v13m4gODGO4iGR+/E1chTRi79Viy
XZdBiEmbTjpLKtjGmn3r8Bwthj8YOdg3UMjRT+0+b7/YF64fuYHRuTM/dR+nKlaX
ZhwZEffItwByuQWC84Vf8f+FFGx0FYVoB9MjV3tfitFAsko93mVzOLKvS+ec6vly
0V/uDCbyno36WavROI6kQkAuZYgCkP2c7rOP2E2MOo5eXAIy2Inh3JiAB/rythb7
qPU1wK5fUJDdvw+P8DETjzqDIuQSfzmilV5+2QDjv2LyZAut0SMXO4fixvE3mzje
lm0xNqsC/kFrzNjdnFyGnZw9KTjmCcM7nwu8o7UWCJBz2aTOq8u/6y99Y1OH3k7H
rRwI75vPU2u9++hZFWuS77O8pyhUw19uZ3T1sLJuV/kZPBgpKIYhKmhfl6Mil5Mi
fLiPP5HhmQJLLpb1ryZVHP31jkeMG/FbLeftQud89V8MhLWwa7WynPYj8uUJeRHI
BMbHzCtFzmnCNI1ecEj5fqEziePqEmdjsrKoPZY3Lymxozv6btzxdhHen3iZ2eOK
2AiimVIYnVuSLfJa3rrsPW1ADqf7GBrHuan3G/Eduhqq8pApacsidazot73Sg/FU
5otHevlLRHDTvF4RnuNuRBMgiKQ4UmnAYtQaVkEzIEP9Stk/N/KNXXww6jP63M2J
t1bey7fHhLeZfK/NSkjy7atlCz01ZkGWQ0tfqEJGeiTS5V6giaII5LcuFfmtW6Vj
+6RRJ6ImFaOOptRG+2jfKVqDo56H51j/0uHPMFisDUi74qtBLikAcDemvEhh7jkm
LEfzeza/+iF19JuD+ftNcjJ2UBijiZnH5PtAZ3T7wk1pk/5ukjScvyvPBi7IkY82
bt+mYQtwMmCD1rH5FX4rW7mlfwROID/0oWX91Ik9i9bUnAw2R1vhg0xB2FvTZC0M
xwcVf7DoE+ZaGJt05X5agrV3WAzzgC/kkNIMqiB7SBPbLXsVE9pGDEqUT8/cde/T
xLA837NNXaxZ4LUUvZKTajj06s/Scob/yslDHdMvXz3lq5gc9tUfqFzTd3+12L4x
M3bMtG7PlKDrbks2DEIMjLeCIAzslgmpsiEercYIzf1Mx9SZ9pULKA1RMWHc1dCZ
dIG/n8cMLjo4P240MOYXoCbYJjoJnEoR4zr/w1Z8zbphwKLIq57wJ6fJdvckuBcB
BsJfZwlOyF0E5u+hg5l6F90WWR2MFJoRla1eQhKsTLVvtSy+NQGI+vmhpw37GKPJ
OZSSFVGRsRI7M/GS0drZetLn54OflxwR/VHw3s1qDE+DTR3CZjL/R50lVVS/0a2f
5Wq2yYehzXEygXMfgB/S6PDXj/JgIxcznd/EHvznfTnesaTWJVcbOplHGAuZ3qPo
DG76WgivElGZsV84l6RpzHla7Sk5RWQMkLJumMIzyIoraMCOS0l3hVhJSS/MyoLI
HMY8XBcZhTv8egmhpmmX/ZjGX7ikaT4Qv2PHCqzTTijRjHQVfM764oXZjCctZC7J
FWQ3rMemoDIS9K4NVu4kgmUdrru1iA9WNSh/3+39pQjVM6EWn74k7UCgvK5PMKiO
OU+2GYhseAINcgp2Few3vR8Ag6Yp6erBgghI/A93ugEkCYv5UFTu5dvMnEothxO7
6bJ8HPdn51zucUryhb/htQ7ScdQxJJjw2YKrIwaaQf3VXoSLVPxHHiaRFOfD7EG5
/+SzGDsR96amJlz000Rmmp93m9Ovx40reV3FfSlzzQdEfDIA1wMPlCF19ab7Igv8
nku4yPlJQUEPQq+Nj3AbLsrYDsOqXYDCxKfgpG6OjPdf8BmiVynheaBL49m/XaUe
JdOR3aBavLctV8vZ1j+Xvcz1M1GwHZOB8lX+RwdcZDwcDNjqVVP21upIlrCDE46C
6g6Z01VU6Gn5HSZUgkyVkw+zouGDvjK81BfAZRgQUtor6FiFhFeK+eMEkeaOXsql
/6xak61JlrjpPnDnf20bJQynHrvpMC4Fyhev3JnGNW/YtqKVJbNfuLnrbIAuuI6W
eNZQPgONC9SzFwS5lBaEOe+66q3lI0FxDzUCalobjkBsGrjmEbcPT28MFhapHWdo
s1TcSRZyyoy3cCg5o452Z9MMDWQKEyK8tUJn0kzaEm0/zaZvacVX/prRtvGl79qB
yaaC60TXK/XkpmrwDw+VBddww/7koGcrjjwuaKMBuB41i8vMGt1ttBOp6FduhFEP
dSLyLZB/ORoJ/2xbowvm9yNp0t/C0d7jGPDTA+Ls3VJWAVVaBQ7N7Lgt/5aPUvhJ
+IeRpEYWMQkACdCvOnSVA9/5laSGESPIm5vWFn4VnBBaV0rWcM7Hpkl4+aoMuHxO
DcMyrG6D2ad1tI+IkzQVUm7dylc8VSM04u5KExZAqC3cQHfjtnHYsJ6hPmk0DN8x
IWCQXuc9zLSdEo1OSIPr4U3CAsPSNK0hqjdu6RNxJ3LzkUbtqoXLPXc5J211UkeS
ctIyJ63La1ixW1X88o0bQPL7ExUXK7BkXVmdMETDo2FBiBtDBnJtm0ysTIcqOzZL
KYr98hl8W24UPV4wxycqWee9TpmsjklqsnVBRlY1qNc3eSS+4Zv2LjtvMByTfQDB
GvnLr4dzPVz4X/YROyvogSuM20dLPfBsXXgpO8EABvE+fhWRdDkRsZiVWutOnwXl
WbMkcI41FeMA6DTJVfDhxb+9H1hrcTnShuG84ufHDytKqn9AyK8FVkrfJGsD9gmY
5TeRGbuOor7ZZEdQs2QPggg9ZiQd/U76lVscHrXo6DVdGLFTu9oIlkzwpOLcPQDz
oXwMKNxMdhkfAka8mgcLTykAoHZ3kX7G2IXIpgND3FKAMUJKh6hOt2Y0AypMMxJn
o3H4tm7rUftYNLiW8MVxoK8lIAq4Lqvz3/XOA9IAZwMMEoFJ2KBM18hNOhyqebug
eDTQqwpbwhnV9by+69YXNucSX3qZXegXywJq9I16UL1BXz7DPEahNqcwrJIzh9sP
8tmB5tQIWm4UmWQHSCvfqx2ElssSMGgAOLMFBIkaqS95pEwcT2Gu5xp+Ag44MCvM
ze0TOf7kje6b4RK8JkjMstabAIdLK8fbbU1Np/Go9jhxDRlqrowNGYBCYZjouxi9
0Jm51IowyEkZs8QiIMvPxnzmBeHsaRIFmhTLbEwm3e705oOh17VPMubUF3cYqHTj
YUS99+TwmWetyFEU6arFsQsGRvLdjNDreJGPCyVaAb228v7LbMk+6skDZ9Qb0IJz
1PidaxikY5s6gsfZoBX4lUN7IcclsN0iMpeiSIwQbDnz2I3cUGF1GKITW6bUYca8
N0o5Vc+rKHCXJ+FK3X0CZ4Nsg82E6opPsG0FSk/hKphSlWff58RhZVXMVD33jzAh
3CLu+3iiuRu5E/Mkjq0WY9yTOm8s7CNdrB5KwpLMBSvsmNv04A2IIeHB8CwmMU8X
6obnb9dIPccTqDboXQGHZ8LjeYzGFMHT6ctxcSUJ3hjiCSczizXvtaDGGE933Uip
TgqMRXqR4zH0AzuEIgKGrydqb2QtD0vUqLMZkvazhqSebhf5X9n0NKlWu+KGCGav
3b34k4rmR30t0e+JL12uYbCtBvq+hS3NJ9zE7ivkR5yuuvWrUgofc7XpS5iff1hg
ps6mToIBxZYg77ztLItP0d3RNlXn0X0b3vUiOGy3FYsqlri/oaQSQOuL1dawcT9Y
u5FPmyX0Mq1+KD3OQvuye7fWClexWYTLc6PVc35r+1ndssJJBWEffYCCZEq4iLSd
pSOIX/ZT5612Vz/MrgqbNIgMyluJZkznCpM+UpIRuhnIo3OJv3/B4XdJoltGallV
w/LVt2Okq7adKgUGS3b7vp84wAUSxdwTNsiTXCV+CBo7mZVwn7R2dgWu3mXCEgOZ
HWSAlTjGKMBZCg3z0MEmhk+8p3RAhg9JlBctc0+6ZRj0UULAVAhSi0TpTGE3lEGc
nvNejt2MdAXzRywxCNYPwNrEN63pFLF+0QGhTzCp2A0AxVup7By0Gpb5TQ0gX34Y
pfD7+ZdsZ/LDWW+0xq4DJBzXYrW9ci3r8ZLQR9Wr6OgSZCaUQbTfmW6XKmtagp7r
uqWZ7KK3ExYUpcF1Dxuwi5BClqGN5uQ5dhTJ0R2+uHUoFNYbue12agvhnL0C1WYg
1dVI51XdkSeR1H7dItLYnofqlDrpTd8lWbZB2VdJ9I8m0HhqdTlvdTKyMSPUl21k
ftSj723mIYjrqmtzAZo0g+ilzoivHeAchGqWys7GTN3Lu23trfaTtq/CNUFhjnG9
QIqKb4A385TO7LCopN4mQ1jIi8P35zlIzu2uQVml1owZSh6lsqC5CLMARxTQwqrO
eRtmsl2iipRorAx+xzneMC/AGyxqGWt1c8RFnmLjmimhu6aOVi5CA0ajhHBc9l4Q
oc/NR26jfW5rz3fLbEz6270w3M/sPNJt6UN+zMBpYnX9BsQZBGwNihHtMZ6YwGZA
raBIa4Bv+Dc0zEgoHwrA+M8hZONr81n8L9cnFX0hYLLvvEXGs+2mxYauQkHfpXN5
x3fnBeBOetBdcEz8sAvHg6yPitFikPs71rsly7YU6rC2IUeE7qpXSO0J2XzWirpX
CmZkYCJji3H+KnP6KcnU6CPwU0tWtxFQlqnLMXypDf+79M+/Howgtzhor7L6uqlL
0vHbukXJWAo1WbgeS79bSJhy8fblDEueP4sE4wnGWTeeSiJ36sJd5hfYcCiJFqk0
IvqYxa4tcTHk4h1PsGLXJ9Db45ITLlxWPJ7VbavvMVfFxjDta2gXFIavXp2umWrm
WziCW9knzgJVni7JdUAshB9UTRlp9mZ/HGBmrUkTrhKSmOPzQWMXloKdF4kwyQqg
4KHWs03mVSDWiKNDyegwT2OPjY4EYACYzST6uHV+xPKmVWXcVhV3tevjQ2831ERx
BrgtGolTowPAdtavc+eiFelHrk23zei9ewInV9UG7yOzZi4cuEfs6L2BPVR3WXsE
OS0Xb21vaCXqZXvET0XNi8zXsJd5O2IXEhxLyF7hhKtbNxHmGiI2Rt1fzeZEnVUy
IbwphPdKOZUCsfrV1e8T3wHeGmUo62u1tMm0r2Fthi83USR2wmTcP/AOMCe2fGLE
4ZP89TUXcxgEyh479IPUnGfDof0oqMewTXG3ViDpxKNBroh1ZaT2lbWXl9OrVj0Y
FR8KhJ/YoCRjIQ5Bv99/mKwVXtzIFdx9TT4wV7LZoYSEuBClUPByxNVoeAIeJSGR
X91oAdb/jq97JUw7I4i8CN9aZJmT4OOyRGslsSPwzhgmxg0vRBtBpBVJMjkKtUvu
VFe9WfZ2uCieMOKBZRa9WX0gKg8dwMUObD9RrqHebL3CfWlmDQzeeLKx5s2UM+nS
KaoWXAEBjaCk+ZAds4yrbHC+Ozn9o4V887Sj6ay5ZTyXYDLak43X4byfLUpuzhBC
+NrGln31LqgTPLS2fsHIoZE9DhdFaXqXjfWA16N9aTy2wCqnZdEh46X9XAqUTXk1
40WXMOoyXiYzeg3Jsr3aSfuqemIDfvfzQkhRrCToWBkL9PhfQ6ImLvyeIWVUZX/R
UjPUsm1vu7nX+ji2SOTi6knvv76rLW0KU2kniXCcvNwaj7iO8BAXTSL1y6qEaHdo
zJ7n3zknAHSb7nwaIpccUIWCxSCxJqpX6rBbICMBksMvtuc0mygHETF//aikwjIj
eV1Ypnv1X2bpULqf4tJvsT36NK3mQ5X96txOnzzdXZljoyQ55NpvowazXKF0Cj8X
lJ+wlQhfNxQidbvzdLUbmTWivuRIq2wIuhoARNk+iw111U9OfBabclAsSj5YFISx
2y4xhvzUfgbtUzlQ4m66uOVFebJcy6U+tGJMGm7OJCtfsMvZL7bPfEeaWxqn9LL0
QwRXBBrs2DZrR6trFEec6LhEZnVLLODgKFt/77NVj5D9tAPmZJ8Itexep/nqE0dC
QauGJQf2TO+yw1QYnM7b0dJZw/yYhJxi/PCHt8eGchRvZC1Ysm3wPMCoC1aDikaL
OviIEGJvazCTd+OOHBwmaMjzUFN4Rkf0y2mKZbolyocoaJaSvI7KoM6Zvu1ntqMf
tr3T/vdf8wOdOqUca3lRyRcL9k8+YDYTJx5FWbpKMCgXEs+lLvUpa5gXYemuwO0P
5P9sAlm6t3KKDFeYjI9R8BYn8o0nLgXSvbWimqis7pImtdMp4MMiozGHmE6m0CEy
We6ffSNEKMGBU9erxbbsy+KpDZaeKIzK/laUf8tsn40tkpgIKghdRBzNRcQImQr7
S5BNO15hd9zfgmr3ItlR3VVHEeWKPduWd57RnyadORwEixv7AnFo5pTGB0ht3Q0p
6ZzqiuU8Ew7AhCEmOlafY1sfn2wW8qYKVpQwHq+S7NKNeqmq3atM/25apL2hqamm
dSVzOmSaCPLEO7F74LO/9H9gVCq6R3nJlwhIKwu1F//YJRjwf2cGbh6/LPDJAfvk
rTdJ5aBNNBDKKMcK4fySWXavRQX8ycoShWp8kp6/j/IXNs3DjNAXpS6qTLvC6PLR
/tvlYuF9yyopSNfw5E5vMzGn5QTgTZHAxQ6/SNXCF5NSC5HnuBVpAl3fOsKgwE2L
364kK93wCtqRqqOePLkgOIJXXPkk8Sco0HeBBgg2tUMT9Mkh2MyIReEjOFHMfSPw
yJtQdxmF4JkLi6+0KVq09U7yGq9/peVbwCToor70X/Ogio7HTk1cq4Swrr71pX6o
lV3BY2xCGb8EDQodReg4C1ub33OHUrc6D84W0WMgIjimiGhtjAzUjCkwsZBq9WOU
dhkO7TYEJ/rsv6nUfBww6KaVeIQfkH0d/pz2I/e3L16rVf1/MnbmrFGH8NYYE+k8
pUYx+4vkkQgkZBp2JOdIAwM8ZThKlLiao+4jK3GXu+lYeRCw6eBsHdBT5j1U8Fyq
qSgmXX65ieeuyDSJhZNJPOMtBfzxFgxOLpXATL/mLhHX95v3QYvlmBNCKkiySWbW
/KHlwE5PfsjUr25cI51UOFM4pzvBXBsbze7BBydZ6vbtUPR3+6kzJN7/L1PWyskn
mTdu+nu/+kr+c6ekRnHBEeJ4U79HS8GBHBWQWB2LJ2XUDazLayR8Vi6nvNjSgXV5
kmhRTazi/pDeWYVsceSbFm23G0cBqRDlvkIkyWJyZKRlJ1pTJYdJVNqpsqnyKsvn
vCyoTxgIt47pj2LNuBvLco1QDDHMiQaE6ZDNFDLK4dUnHVgPR+V6zq6SNQz2B4ez
gMogeH2t1srF04uMM+w0oMmis2uWR9PcipPLsPvmc+Qn74Wswn6+sw29Na3KRx8c
CzhxouWtMUX23LwRpHiZKk74J+WO/zKK8jS0O3wQZd4ekPgmcx+nnnGFjkpYxlrz
agHSJYLvn8RDvicJxQ9t111MZUntZdKN1TKDfAVRArjAlirT04kwBrKWsIHoFQUN
qudIIIAVJQ24pZGrhyNwno6kAbQDPWNhN9FcJCAkk4Pf0jKkDuJyiBGCREzumNiG
uLX0hPaiGgL08ZgPUvmKrJV3VX+6KqzaLhh9pBItsjXMCDBCjhH/Ghdl1oQBoP0I
nj+NyufaqYdjD4JqjSOs03TqT77wP+IXBtsini5a7wZ7CW1XvZRHIdAMozmG09Jh
ctxkZ/NzC7kYwDse5BQrM40V0zNvBesmAZDm/niNlVgZXuBkHQswMP3GawMZqTZV
1sR7bupwdJFo+Azc0ujhv4TFIv72RNNh3fZsXrTgQVN4TfqNUsnCKiYmHjXph2gT
3c0mYVYsvrTo87hQ85YAcMvoedPiKxD5w+BBEvXlwO2+X6VJkygYCli0DfgkEUcI
1KBmfHMG7Puv9j567Oh7e2tu/hpHhnY4uSPOUXOyQQu7/i5vDrvs5Z/+dpp2IwIL
KK4dUuOuszQkHbPTXPI31Mf8XutyjeoqACQnAGR04yAe+YYT8TL5ycmfT3ecr6d6
WXoMg3fVakezgwxfm7bQd1uRIKVMWfH8SuhYa8lcy7FNLTIBCewbN4AKktyJKCLv
ShsLLJz9pAbEuWPWpSct/hrKl8vDJNqzDpWVoEkLheJZgVpDGAdI6zZAZ8QLFYB6
6PHQDtMn6L75ryalk9cSicy/hHxMkm5HOY4CICno1CoSfy5OxZHnVhWgw5pvDUCd
Na90IVw0PQQHxeqaHJ8F6+1LCgg78m/jWMSe83q0LgAjaU6b6gP76H1rwxmXD5cW
LWkyFuro3i6wRfsD31f6uw/kbDUdOLtNBt0FU0ho498GNJV119GCWkjic2MTjAaE
DcYeb+TSGFJ32NCY+E+Si4xwJd0BvCJcsCHTDgHXPSO/fo2WSGrX0t3LpUxfRpHm
udG/Jh/bPK2jDleiA30YThq8kybj4AGd00EQYVLjqHbPv0I5FQ2DL63iA3OPJAMd
ObtqnPFc79BW0buh4aE5W9ZVaVi7o2hZM5PYcCNcjHrGoCRa1EAhlX1eaX8+DcV8
XXPoUxEbrsNoMe0qMm+mNG78ykBwWj8hsCLdpNBDXwaLGfT/H7fjMKxLuPG2suiL
XIQDmR9Lk0VmIk6x36jc8WV2kv5JoKzn75Md/7/I6CBd+iNzVN4BUGQJA9au91Sx
UNPB/0WWOJ0eBUfuT8Y/3lSa51cu7z9bytzGoVD6adKn/u45iZmaAAmtCnJ2otPp
bMYMjAIAqow74HUqyrsAtNxBJj6YXuYeTIAivHakfGmQPyeRcjjxbap59N08IQ+E
u60lg4+gpFnNy1ryLKaJnNm49f0D9lKA2q2jlRl1dIy6FlsmdIc8x8TGcsbzUnl7
e/D5zDqsfYfOn8/89qLg5cOZlrumGdvHNXuDPZ0IjQGoO7/2tug6zGSKaZ3YIvlc
WmFpuo89XQnPFP/nlBDRNiPpLcpLtikM+w+KzmoNNXzwVHI0SFFy4UONXLLILue/
3XGPN2SY9eowy4Co4hhm9SH5OfCPCCV5xH+Alj2G3fje2x8W4T7kEo+L9ca+0N4f
iBnakpUnv6LFXGmdGI6B7GJK3MbiNpCsfLg31amFH2bet2ZxCwxdqLXShpDIronp
WDLjyFcDnYMrVUNKz4vQ2SMDXJjYY+1I/LyedKXJjmZ5MgGtLEk9VpTzgQLgI8ou
jomW66FvPgg306jrM5egPV8OEKc7I7FsOqRWFBStLdsJXQE/yx5D3VJ9Necrl0Mo
GmxJ5YipKXRYnMq2n+weJW6/pNRk/IU+B35KIzT4ozuv3jlOKIGZnOSzAFxdd/yU
r7y+k1YIZ4wpjMmmsI2UbjngRSr9s7gYb60xCgJBywC6Mnb2BceUq5d5sYUJ47Tn
kGkm9UlGRXpN4+fojuErwOnsmwuhtQsjfkJ+hRVNgbFPmCOFgmR5HLCoD8IC+ZIQ
vlky4DFtH8xskdQuGbEljhrfMF577ezC+dH7T58KC+yG7Lv3WusechWoMJ+1EPWz
pZDFwgnoK8bbUAdvJ8LhJgckOK7JV0sxw4IxE+d2J0Ns88tdHLZhpcp5JoKHIOYF
kPlDyxXhMsrN5y0xd9R1jfe3SjvcFHcWY04jYBQDJtGBqE3SCWfOxD0rqDAeAp/9
DwUP8vv0J5L/VSMRIAZaDltUwRunH7BgVYZaJRpyKNX5GzsRqEEJoosuchMeSx0W
weVeDDrWUYeqXXCiNlAljK1ZNmOjRTDsMb9kjQJSo0KFTeXCbyYFHsZH9EqiGc3F
ouc3ztBqq5FlK+xoBpU8SRH/Hdarl5/VoIkTIxDZrsG8tgMMhl9B/lehDEPYBbw1
RvaOytd9iFdNdBPxg+lTlROSTqOsimYLv4/GAAZsjRnWQaIt4K38j0Ye+0Vh0h+R
ZwWKng9Uy931O21l34g4eXfAWer3/yy/FqP635o2VzdM+TqAVW06yyolFFy3y7hX
Jmq1uW00ai9ezJUq+7T31rnXe/RnEfopLMMGqlZMWOwh/wMjce+++g4drSNmgRuY
NICTex8Ial6WPNCd8R3RcsGYF7H5c6sf+XJJOfiCM/eLGGGJz2D2LYtr5Gs0KEOP
TeyLJ9lWNzzEyII0vVQCOMliGasVrTqE2fuS4Ep+cTaa50Y4OYSe81Kn3Kk0frT/
bIRvGDtT0wIXp69Ul+ZwL58sgmdFrZH8+DvoXDG9MahbPj8oanMLyAzwEQMS5LZv
UuhK+kE07DJHJN6OaOdL0El1AUYpp9efaZktoYzKfh/QvodeyEs5mTApoXFD22Kj
L1jqanYd9VwVsa6j43qQoGjOg9BC5LWDAWckulDgWqf5AalB8yR7z3pHIrEfo4Up
7zwVMbIf90mjp/alYJz8JpPup7qg332D9EZ4IsroUc17glPD14KhLzzI52r65AuC
5hS52ReLeO/VQ+Qi2o+bjqO/NoPbnbpCTMI6VGMYfREFXgUtuGqgGbBEsNH38nAM
hje5rRNKPqW8Kdl4KC/yFholA49zs2QKhUplekFxPDWEok8fbCjLICVIap8K1Wwt
da62ebIcEWgdOQD4KcVfywBicSdzJZyb4ZpqMEHDN9LgnUz0IB26Q5eJ21htRLe3
yatXsFBjy8PE89x2l3LNtyP3cNekJvkfEfn7Y18s5lVPgFgf9iegA6wtC8xYUidd
ml7vg1vP3UQGtCQBZq1+1t5SPxKLSSp2zuwv0vMvlv+WpiSCZN13pu22ZyiWMeDg
m+b6ET3PAyUrcZqx4TIYEYeOVEZ0pYUMGezIif+8RNUkkViu6lcj5FTsRPXjQlQe
wT76uNu1M0nubja5hGqZAg6u73TS0kwZtN4CQXWH8GifZDvM+vIncUJbhFjwMUCN
z9Lzwfi+hJV8WeYc5nv4cuGwfM4zEI1OUJu/1GTrK8N4XdykSHN4NwnwVILp47Yx
pJvmntnkzYy1eMEwttGNedJ+BCS+MLYRgbclIGkW7eZEK7RGgq3PlpQ7ezP1/xds
52xazVY/MCJr1DSuUrBWHPMWrizHIaPntWMR5XvJXt1MHd3BK792I45biZ3Q+UiF
qSBQWYPjxOi35xnkSyfihj3+fas+6pRccZg7VF1IJX1dUohUk0+1cNQrBcRuH63u
5GLRDmZpb15E8+51vljWM/V7y5HtgeQR1rzzSYOBYeb2eRYQ8ddALFnjQRg30G8q
6JarCfwqOHZsVxdSMWd3JiTuKUFkOz4DFXPNbvi76kEz8rbgNF+ugB8l4QfefyLa
mYAqgiiHc79WR5pL53GYttbSX9u6ZfBoQXV1fZmFlhYTcbitOa4j84jlBiCmErzY
vW+2uYaKfWg7EMtpCnv9s+RzCvJeWSKKcS/0tQpyYYOEN8LnOgCDpIpd7afbeRch
RAg/KyAsg7zg1qP9KrycCmj6lIVRJic/1dDkw1uCMlWdw7rt4RJqYb4F7Ks+0gqF
WxVeB2hweIfDFEXSFmwV0H4AxaVLy4/HSEA/G9WLpQZu6RlRpv2452y1dwiUiLaH
wfE9fUIqNAi2CI/TPHaVv8iIY4o7t6Y7dXa224Fsebv3mYk1SBnQEDIZx/HlTHfR
NMTaXZfwPAJ/WAgBk+uEFLATesKQHyzCaEPyjIrB3Wq6WOadYx+O71y7habYzM1d
sDDXmukxr4i3xLcP5D/SE8j4IoMtNOWXNbD5IAGVCnKkIt985kxNApjkEYNWsCrC
DVN1ieqvx8zGIat8zQCMT/AYLP2B9JTusg+o2VzkcYVM9OLuHBpd+RUn/zvxySpm
F837zlAcBdtmGOk9746zV+lxJW+wZ7VSsPFWynK2vfiDX9my5fgCYKxqZ9qa2P09
MAXKTQecXqWPepXcTUPhojo7u00rmMw4DJaGQVgf/GRsmknsY4AuhJJw//km29uZ
p2HrO7dftq4b6s32dPOHCDncY02hjpUznR2vk20EX7rmx+ulREvgq8Tf13mIgQnW
pUYu6JQtNZ8QcuOneTGL0i0VlTDACNMOCulhxBJAe5CuaIWEt4kKqb1gT54a0Y6Q
Hej8i/as4R4fGKiyg2btkT5d3Vae7Jv57SXz6n+2fNMjlQRpuHSUXryZb6Kd3HIa
sO8b9h38pX+T4YtWdDpao9coz+5Zx74PrEAxt3SLF/UkoaRwhXngyY3Dx1L977sn
+mpkVkN4BYfuolGbLcwp7paCbrVnqBTL/UNxu7s5RQJ52pwRFwxSOSE3DgNJNmSG
h6ldWpz3M+rPI3IwwaPl/lyd7fVfFYiGq699qt0hA2hS9I5R5DC4Te4TVdBkKrDO
IY9MC+CFmyMUKvFw17uWszZtqbLFmqE/t0UM810pWnVHIXZgi44yKK6AZw62VOF3
9heAJs7peTuG+rLdSdEidINtdxT40kdsPIq7FiL/B7SlGXmpA1H4hdyOooJzDWGz
3UOfBKcDP5LzbLmaxfJ1pfR4lTT3FVSTgDkWClcMgt9HovSr1bQq1zX4pw6D/bHt
ZOm9y1NLp6WidVRkQy/Gx1E2QCH2MUlI7SazJ+4A2DOXO+TiG6d3XHf/dL+mFAd9
cGw9g0IRegU4X/fBRTwzA5UKR7vPlz4yuoiUadiApi0F/JAc/Qt+V+ofcIF6GF4e
viIT4YeCRlP0I3nMdxQZVHjBXfUtL6RXZnKpDDHSYNMZ2pysKHbhk80yqG4iSC9s
r+AqVxMSYGr2z8QfzkyH642pmT/OUxYtWAEoN+Mg6g9xFvw0Ws0ri/y/Ngd0lmZH
S9U5CyMvZB/+nP36kc5DyrJ+KY6ddHBGK+mHj2ckrbNwN+vDEBSoXHwIMTS1BH09
wbEOeJBm3xBwVwrH4rZ6872F2ZurxXpkw0gxBLFz495e3kwS7Ojb6QoRucP5voPo
nnTgJlNulmTFb6e4UwjHPpdZSYi2Q0M03NfdxAgu6Eb6oCUQ02rUqu6ftysdyLb3
mRTHkLmsxsutGh7jBzGmh66N7aQ6BTCs3iZT250WomaBOxxmH922jYsdLTyYjU6K
IFA/XkovOggXSxaIKmnWYUTEeVqbhJUn1kUVm+8J3Ff5ZX9rt2TEWx3xBruD2l5M
de9miyk33bMuPYA4yxVsrW67o2PRvy1KhXzYC+cHrwtfUW0sv+1QQHMIDOA+tuFx
BMvQxwCsdnVRSHo3ZeY5/P5130RraqqmGaVF68bbw6ek5vKgiVcAkJlHj1xTYXU9
Sq+mjgk3F+7TMkVrDHFjuCvXjJfxnrZHpn+qqrCTiNFxN0TuzjcEr5RZR+jAWTYn
JqmjBHr29eqv2mTiF7dkSwCUqEp8Su33thqyS7ixU1YY77mMsIxjLtUuJjrDFb7F
f0HmkJlcVfX3z4Q9UUj68rlpXLEiivYI5CdlN32oMy5FLkg/PmQFHAwTnrJ2wo+R
1HsHi7JHfTl8eKW1zYjqXCnm9Y5pXt7694rLm9vNhDdlcaOPvk0lBtbbEwKmTcwm
04wg1oWO8cZPgHJQMhOpZuZqntwLKdMb39TRjVLiW/0/cwocy+p2DGFwS4S59ErD
evkb3kJOaD8Tkxl/t19MwkrLnpv2vms+ovLwW0ZpNG7j+rNlHdiiVkAMqjmhJmX2
2zeCCJdDhbVZHGa42xN7R8wfvzPwW26gsCSbpxSKFU9x/14q1wWCRj3QhnOO+2aS
dXImXuMnPjiXdaTeDZGudO2PRxrBgS3RPZNXYjmQOdACgRNDqqmMW6pKGMGweYEu
XMqaQ/B7Dsbkvbd3Lb66ozNQt6+/UkGEMZ8ITBCLICmazt6wm8oqEViPJWBwtPm9
Irr4cuxRDRanW+LuZXAx2NI7Nw00mt7YPTp0O/JrcXvvc0U5i3Cv3M+xV97j9kdz
ggyo0xWYACbbHhDjxOFEZ5eEd4SZlZhNF8ThI4Wrm5PvFu02bXSb6Z2/crA6CH3L
8WZEBkGES157uEItXN58s+n5ts6pBGlToGfxe27+KED/R4aYzPk0ox2954fiHw61
HYKt98lEjJwXTBmpwgsZVXv3/jufcgLjuDvXvO1E0Qp7FV9QGoGFUI+PdG16ch5/
ORJ+hi+rL7ZF1grTJ5ipzM1yRssqxJh1lhVwP6GHRb4jA2T2yYpa0UlAOBVAQ7Up
jfUCigZPzIy6M7t7EEx+n2gfnKT2XpXRJR2VmiLZrAneqJ7gBD7XiE059BH6N48t
yI7vfhAjy4QPwMjBXa8alLkLGMThCWu+A7JcAUPIKyova0s6t6Zwm7nS+rN132GU
ZjfSQ8zM+bJnOrj634i/oS/hz3oU6M0iO5279XHyejG/F59Z0lREHli62lsM+Smq
nMDRqBzaNlOkD1Lv8AZ+O8l5jY9YBN+whcLcLwPI5EDItOYkQIcL9ZVL9Jmdckrt
vIr+QXTXK6pibmbP1+K/CnaUMJpnm9MyJHbEGrevBMOWWQwX+0nwHPBTJWNgu5q1
CPqBVNkMuFhGEEKyOZ0lQIuc9NTaXjojDaNceiQK7OqOx5I6LCSXn6L/cAo96PxO
EYzT3BrOVrNEgN3f8Zbt4ze55N5/ogwNkNppMN8A2vnnrnAW4RFCwxe9kczGpZZz
8zMnTEhT8wUJE76Y4lqtPI8GUlb6LA9fNBdOb+Le5PzEcuGrhQmDVzkqZEd+CSE3
FwMfCOSTXORRHg0sjUBRHTN5irFZRTVvsn5zNN4slm9544klqSmdihmuZocHyeGH
7D2hqd404nz4iun5o2eWpq8jSc+6cIh2UN5zjJ/d3Eu6iVdTUBhWphCEULnj0fK6
6rGLk36auyBq9gR4VkKJ/VgE3J/qFIJSo3rC0RIGK/ywWVNZaPH/cS0zqpL/BhtG
ubQv9nTM01nH2yef9ThynSANx67BluaSAv7AdTgldMNnBnyYt6ruGl8dVT39uNdT
Dq+bZ2ZqMoHQ/4XhXvXYv1ulRIzx8pbjYx9OsD2nWB0fP34E59POylLqqNvGM/la
GH0Wz7xDQplwAf2k5rq4Kg2YDODi201mkGO/NVaXxzv2qIOdAXAwmal9TDzqAh//
8yNt+v4JXtBYsQzUili5zxyqPvYAWyk7oQgItmSaRQSr86d1ujgXAgznhg5Kwp7I
IyuTF3avCPm+10jgd2sd2Mg0djakuXz1ckxCiCK0heYU5xKxTZveLMb4GT+aye+G
TVkjMMAg5q3WWNx0DcJkez6SI9Dy2vWVo4ZMU7f7p53DPMX4vbAnrsvQ5Svdq3nP
9KZmK/R4jrIdfvrrFd6Q09mc28xrgKK51Lq/aKBMt2X5/HibhTdSBYm7yL3uUvJj
wL/IJOG67gB1ajkh78QmbqDLRgigSFAGauq9pM5/2kF6OcqIWGOttekkHKnRRsJj
9eAX59f7QphSjzsie+1mGFVxGQFpoAF313ltXUHwX/bhA2NJI/3D5gKGAHxnqmJu
PRTeMIaTGrzrp9ePDAXQ8YNbHpUEh1piz0hFqI5sdviXY6iKwDAbPAeNxQPR9oSZ
GLdT7lp6tp/PeyWdoTDH9XC8ORoEbdZ8gorkXSaCMVmIdsyPrPyl0OaA+cpvgmq5
Liymg5lckPk2xVMfbS2+l8BoSGWQ4pBNbBPwla7+vBiGSoGC2cTDZRr1NRvkWjqN
OuLF8Zo97lcXPoDtaA8Q3f9gh5CuSH8RmZfHamgp18bMtfxEr6vPgTNk5icisn0s
0YYIRzfvDKBpe1reZRf/YZ80or6URDM18J9U8fGPUzVnx3YVJFll5L+eafZFjHUU
M8Ni09rr9Oy6fumnKyqnNzMrTN4guWYQ7pTy7pvtHpuIPbH+4PZLVj6y0/nRk6Bv
h/Zu4bdU7rvCz0nrfrEEzUQTyyD3tS0INC8H/+AkJqEnrzNs43rB6SGeykxB1/CF
UL7X70pgF8YjQePjQhwI9fqynL2XxO8vF0mRaLQ0xhQBQZUe8G2N/IbLDcoWT1c6
f1bOxsl4cMXRnHk8ffFJMFhpYJcPbhvrDwQBEfvvxMge9bJz0qj64109RbKXniHJ
3csfGC/4xBjW/Ch5AIPC8QEQnpcFN7GjWE13oR4xtjYb2IAG96EXWn8xPu0ko54E
KmxDbwaStkMZQMPtMvsnpXCs/yWWYZgdsHF4q2Q+u1aycFkdRd/PQMQvFNKTGJSG
RqpilufMTS0yuDuT3PasBJjEvSy6kysIYDNLZqaZRRyymCakPWzoqIpb9g0zsPP+
ZGR6rwcFYiu9lBLRNEqzyjHjK6fGbFYKfkQrfoE0anUIi1uKEJ4evtZ6kXtuefUr
U2j4pGhnuN1py1+eipqN8naT5G4Ij54wtd+r4co3AcBIfhSVj6Dln7PLQtYctBBw
6GNQ1WsWct8XU2zqdymNFstZSwtpTKGD8I5kk9DE9epn8AIdTpUWemqydImOH5Ao
QGxFZLKupcRNd9Q2evias3TEzN9rvsXeFI27eAhQRoGVt/nAU6z1L2/t0e4o+/IP
HkebplsEYwJ/RANQERcrw9JWqXsQ562rnIOX2SvH/Rw9yrWE9u74x/o2+doy5j6w
GfyzkgfOYds8vPD0FtIzAE9pDxvpBho6aYUCilIxrmaCflQViV/pVnvoxqoAewWq
xdDYLgEzF6qjh6S7tIAXunPwdAdCtV92iFIRSbdm/4ae2jXvN8pqm6HfMqz0R3J9
Usn69YOhIT0Dzak/P4H2caOD/O8fasSkZ+FGbDlPvbvzYVR5SMrAe3Ybtn3PTJRj
PYIKHtYiEsnbXP5ZWnRgpjyCqDmbATZ2VlPr0ARVhzQ1xKPaZd3fFEERVrolgfDb
Ezyl25Yp3GpHQwsDuNAch0X/f2svbx0ORwomhXw1mRYo9zjopBaV+5WcqMDAioVW
KmDU/KtreEDMWoth0bg7RlWreSvjs084U7Fk3cD/3w4jJMG2Hz1vOABburuccyfB
+/++M5Fd+U5MSMh4reaIPR4i1hiwvxLx2iAaYmDrWtuCVQWTgUqXMvYfv2Yi32f7
kde1SWVd67hUsran1J7u0FTqiW7uj13RF3E57Y9PQrSbpQEtZYwJT5YlD+q/H7Uz
Yp1MFRWf6A4QH7Y59rIPGfLdewChgxt6uGdP35LEp8kUfIFar0tukLWScjHxoj/E
XMPAeyguoehxsooKU7+yt2pUnVaA2FAKek/Jt6F1fK1JibyaeXdyk9I/j1500v3O
bnzGPn+dpCF6i+zisrEpj1Eqow9S1qD2VYG1EF+cL3zXV/yY7PEOP95gPoQUqfsX
Ic9e2cvMWjKLgA3GaGZdP+TRUzRbkVbY7Rvp/mLgkBVFdcdn3jfMZTT9veJKBmhA
WHP4HgJHSwEy9j1kX6qic7Q64A0FQEZi5IaD3k02Gh16Y8sCxg/zGy7oil5vEqDM
DtwPnY9X/v/1HV5NCts8Cal0Y/DJ8Fi/BpbOOAnKVZ37GM96vVJ8XXoHRMv8k0pI
z7Vx11tC1sZ5tOm9qgzNWKqQSarz4rfQ9MhCMlmrbZ6eoUv+axRp2lZso0n8SAEX
4UmCMxuujbovej/tnM7CRTvB+fpsQaOlZoYdWId5yvbEJQq458rkoGDqllL68bH9
NV/Bm1FjpHV6GSm8mrznG0cM+ye6FZsaKt8nHIRqUzmCnHgPxZXdWx8NobQtQVA/
O9P6sprB6v7ZwGgbJlAmM7AtXTovsK3Jw9Z07P16X4kqxsedlRkugPQug6ZKY/Mn
2OGL+vKYrdSn6ZVqvy9egYzoCf0vk9l64T+yW3MviJZUA/AniD5XJfBwOTtz6QKs
5KV1aSWFrNGgaz+Va6TnkUl8SX+dB+vBeOSw/vEOhn1NVYAxuu1KvkkLkAH3+j4Z
9LVPUX2UwJHHdPSqvHTZb0vltbtvn0R1z3WO+c9U+P4tTSEO3sx0qbPp8gOIL7cK
9IaMNb+kARY57eF4D3xAveUWTNDO5cwKH1goH7FOK6I4qhDYUQgTlacTSCq+PvB/
4IrQFOJ3/QvtdfxOJrm8mbs1ZJ45G7LOAEFapQ7cHlqyyu+84uMnOsSUwZR3O08Z
CkPmVxKWm0ZJrdkwv9hWTDIAo58PNm7z1i+1eUPSN8p5iWm1hqli0oTxnPlNcfY7
SqgVpwgRlmpTvKayoc9+HyvQOuS51A3a/QFM27rhVbYDCBPQPsAn8GpcX1YPppbq
/RRndeWPQ4I/zjp/YiGzkPQ+Lxoi8frtxEd+F3y1OANrbbEkG54CuTbxyc8LKQiR
0AXZPUEg2a30Cn8o7/2QssG5xzypuHCICnB7kqVNZCx2RRAQzqB2P8uuzsVZRpQ9
KHNZDKdtyrsFRH3ZnoSKannSFWaKGP/0H/0/CnBxs4KGxoM2Vc+h5M/aRWF/M+FF
SH5qkYocsi2ST91w5hWXarr6ZTulJaI2JquU87OVvNtZtUdz95OAyOtYkG/PvkU9
YAHHKP7uLeCzA8rmJ9drbRm0biPTfV0z5mUAEFka5JqO5VvcemMlmAEmKDq3ZYuV
X4x+5o7XSY+rY2vnp0EZVqZIhvP602ySmYt647tnZRXVSmktU7AvFJujZNUFA6j0
6YjyqWn3ljXCm4frZ7HSGvO3CjyLxxPj/BFtcgJJGFm8/uZPoj/UXLa6M60IWmPO
wY0UjMuXKxfq8mi4C1aZd/jF2jdgk6qLX2TObSSdpSg7tMbotWFz+XF9i02/LUVF
+qqMwgx5VYV52rNsWZN7MBh/Gk56XkdPNAxPKFm0O7OH5nBu6Dy+HTi+MkGJ93Gs
SzBEpaRXwcMzyfWQAxUyg0cNtKVmKhS0iGFMyRVETpQ/hTOqdQ50eg4VAgOtM5Jj
sYKFQMtlGyVFme1fhX3tw1EfXs8SA3vvQjRem7e/TpyCiwl24sVbnl72DfHiV1Co
YJv/ku+Uq2t/Dj+vvX5STpw+NAMevL+OWTyYVA54TK50hhbGqIgmDtu2lcACsvNs
CptG8yLIxNzg2GuegD2+mcd+gWLgammjocc5Ey5lm4kHTS7RAyhGlehDsACdAlui
DG7YSxqJUPOYh7zygrZvjzP0y+5CkwcyzNP1VlGiAzjhTeo/NR50IypCnRcw7uEX
1uvaf+ECFkTFaoPpnQ0Br6/EdYx5pl9x1OvSyvNWws5wipqsWCEkBAoPQiQFELdH
/Vb31TNClimOZSw4mfG6K9GoVo4uaE9Ibrc9q5rrQGe94dfXooIBdR9rVOcgpg3I
bpcSsf/5/a/WjJiyNA2LeMMLQexfj6keIKn3wroLcdZVrsKAo+C0tSrKpNNm0Blo
kbBNghJC0INmGttdv9taAZeSW8IZ0BgKB3T4a8HrG9WlKNtdx9+iWISxmQ+E2UyH
xtuHrwGPwOeMbJpiA5JG6GuDuztXFo/MjYtkaoMJDR2sKU/5TNib4V59hm7dIhBt
OW4LDuSnhD1UaHdnLtpuz9hyWhFcS2tHPJFi5rtsy5uzB+rz9tbNw/YdDRhVDI+i
/+6BKhhAsGG8mMXWAxU/JEraTwdy+inTQW5IgQNTcI/vtYK3RYHVUPwPQ3q7gT3Q
NeUZgLSuRRxvIYDWfne5oYgWAsHkcArEq6wexGOru4WGIElyMEpJL5SiUHqOLFUO
wtxdcHQ8Myg250JGYSpqIesOAe+gVKQr2YR5aS8qnNsmVg54RJSJZsEuaFUjtXAd
0GDmUOQxKklT1wUoBN3w6FeQlLQ1L+FpGjpus/G/lbymQmKU30UHn0h9LmuFujtu
E3Nup1ISdXY8/EnR6ItQoUtNFwEQr/IkM2+D50WkqyDjLb+uKMzPtydhYRq2qx9I
dyI0CgyLuQ/M3VOjCGNStzaNlXn6BvBMyltmTaEGANn4XgIh9al5GUSRxD3Pr1/a
79E76mAZeqJ30JqHGt/WyQtKL8Rm8vG3fuxiHKi3NcYV39B1bK1B3MjNk6roUtXu
WpyqbMuLBEhoj5nysxEb0/Kl0u38+jPQe9YJaR7nzt4PVWxrigJvbM0KGAFt4AZn
parid5WKP3Xiw3n+v+m+zqqb4tSWufA0487JWlVUF6JGLxToDQul8tK7PJHwkQ1h
N2DldTI1IggmEpx/MR5TZpagilHLfUOYxspHCHG9hwHTg3hfRFgSJYCVtmlIGMJX
kdN+Hf8M47VgudF9+QLVC71VWQrj4RywQ0RKAdPn4Lg8PIJ9vWzTuj/12UXu9Qqj
wRgdiocN2dLFdWXHQUF/eJBhBaT8u0hS5bVrmZovwvLUStwwLtohAtfXdZKABleG
7Wxxf8sd7laIUyEyTUJtdNrIfihMcFHbc/FbZYswyrDOhejDYUy13bsCNwPqA5Gq
q9k/P+0GRp562YdgpCfKeCW5Y6AEW1I8sJmcGNFmA8WneHLE01hHA/T4tI8cRomI
lV13gQ9az88tQhwuyecYNej9kItEkFo24RcH5xhMNUUZziPGJ8CibgNgc+2AUK5P
gewVpX0QuGIydBUbcOxTd7CaZABsvE4JzV6r9cq8BDuW2h6yuz2H4/EuyFHnONSl
YN5u8/cskDu0/S+f8cLEMMOXMEklzUib3NXnIzdWw6uMboU+b6lFoQVTCR/g98ny
pgzHfWQs44fSH4A9IhpXPI9HHTa82cZZChoYqwxNRtWTMUzVPKJcOM6WEJDtNwSq
XHL6Nvyv6jlFnO+W6AOHnpSYPEHrczxyCjWA5QqN4jEqcZ/hLkUTc99j196xq+4E
+OuDNXLUzZLgzMPg+z8jI8Y20ENH+KSHjkCofR1U4MbvHEPPXM6PpuC92OVMHHBG
SsKmKsHzgxhJNE6j382XHvish7e1RaWjvCubtgg2cKtInqF2no2tKJWo/Y3NnkiQ
wSKxsitlp77IIyOElk8Z4EIRXoenVlndlvb+8cRwSaigCgmBRDRR1+xB505FiqOD
iw7SDNf1lpq8S1rWVuIafjGlOxXnmBSeoGQqA3ggTEYy6ZniMXGcqv6EQIzQBMpB
j6HivDNbkGX/YeZHcN0zae5DeVEzXb/tOmujQgUL2PO3L95RPpCRDz6ZIm94f5kS
YBpA4izEmXxS32x0gBIaWwLjWyTVU6vnBn3nCRugj+PsyuX+ceBft864uiUl8CMq
p8oYtMROYfy4Ozu3j1pVWw8VrxleHuHnoLDbg2mFzWVo4//1AaBUdremkI4GIyLx
NfP2Lq2UJVoTdR/8ChjDpihamMqbN/6LTkql1N7z+Fl2FMHNNIAnlDWk1XH4ISI7
nkrNTNUWpRMgP/VmoUG9h13A1C9YRGgCO8FjNB69c3ua2uByyxyQu3fpQ3jA3eFu
8GmDf7Ndm6mBKSzSIjwZEIpb1ZOOAC7fIZ9i0J06tWT7nk6ApEX87mr6qROx0vgk
pntUyd2a92pzQhS2mjBYgrODU/pv/gUziQx1W8n0sZCWvJmObDI7SQYvgHz3bH9G
VFCv9AJwIZnzB8pbN7Emg/mROoJPwQpNnKXvCXfM8OqqBy639NQDmvFVonUUx1Zn
PyXKy0NtRKTgNLxeJdhWFU7LvZJM1PyKVzTv8MTU2dd2YPOxTPZ8R9U8ZD4+/0f+
OW4mhIan/lHo7oW06alGUyFGkE4nbNIjHihQor9ZFhooQA4loxuwLrozen+T8IbC
0SVHqGr864AJWgl1FxbnS5129B5usOgl8IKmP3PZO3hkMuyJbKu/D/9YJSUSOfeU
21WCUt5982IjaUYnRTdIoUUXshFo3RbRs6+dNZWa9WPG1rFdiq0sRgxr0ka869yq
ILWXf8TecYRvyV1t2lEzKYWREOyiu7sQylT78DR/nr1luso7J4mIO4gBxV8aer61
dfb7yfSJ1xiQqDAhUGjTjjaYTb06bt4hIquo0/fbkEUVl8/B6w+hETg9xvWr3CnG
MnW6k37ZDuFZJcLLuYzvlxOevWYonH4RGwJhJsjFi6A8kdzY9uyn0TsXDrsyfhET
Dbxm35rQq77rX/2XqmWwRB7I/TdIHNaPSl4FgqOOYVsqBjewy/dvSEe/5Jq/1ESQ
Zq0agkseB2BJLj81f1fDXZXj3PCFOG0Aunyx0qiVit+DZBxGOpAzV6Gs/vn3UEBP
Dcy6ZXnUXTYGL2q6hsS9WL+FWR1g26o+zAhedDGPTFtJvVmDG/jOsTNt0F5Hgb4B
N0S2NIxAO07QYj0c7bXFlMlia6mCibw3F5mAe354Et0b04FWPYs57VwQdyUjNBQX
Tq/FUkxCXcvaT2TxDaMnprrKEhZ6kXTw+wSPQscF2GzRr9ktJERakAGTspdvBhwH
gzVtkfDRnr2aXQaELv1wp8I3GGkiXlrYwYKyCK1tloDl6s7U9eRtFa8qZ0IkNgZf
g8WD3Iq1i4XKb75ZEqieqm6nt4evtp+xpHbdHlhFN6W/JC+fNJp8VwEQFUYKbVgH
kvxX/GG9Sc5ZKONoPPpg5o5jKSCIa0miqSX+ouFztwHboFw93LgxypjYh+b5iX72
2hzMYJ/yCotlu2Z7Nw8iVOtpoc5JTR732A3MM8oI2wM8ks23aL477BZwAK1wnIzj
amMQwMrufaEd7dYsVYb4m7zXpa6NyUhamN+D/0sUPiHypJ9An7POP0pOyLWgZIUm
zPtFi1SqeEjT83arzAALdcTfKNMG7k7etwzCFi3IpZJUZldXNXJUCjWAWWyJJ2gd
V8hvTo2v4wUYir/W3hD6fUN9X9aTQOBU2UKx32ztsp9Zblt4W4sn0r2LNIS3mGlI
FwqqZlnGZU6fDpkeFOLDiB6ByTPSDs8lY4dYxZUMFJO3g3Om13NuvSHl1Gt1sR83
Bv4tbfTdrX048PJ7dYkynm3tebtXdzy3MyXJrBRZMHst3zNIRxC/oYt84wFFqod8
LWFuon0jsV4fSaN+rDd2b9qtE2Xxc0FBVIKk4osDflccnvZ5fiYOHwyOsZN/KQBk
jYNIJU8VYeNHxEPh60e+HywB5iA3WrxH4GI5xRQZjj6Pytg+rHRd33ZngeTdPaW7
eG3mQl3/WVWOlQ1PvowSnn0M+5aT7IcGhKmxlqjBGcU6DlnPd4vPVsOohjrAw+mw
Scxw7n/wyqUT9djpw1j7Bp7EWUFWi/CF3e1yE0p3j3bgQfIh9RNBN5qkd/oGB7lB
8kA90JgHk39jTT5351ZXEgzd+exxrxiCnCGF/OpbfWfRQMEEN9pu/qR3y3iP0zvv
h9NkwrNjpADA+1rAHbO0YUqrbhlX06y9Yf7bERKhqPdsbQ0Owid92mASEeuY7Fun
FdZ/won5q9giOjJaGwkBIFLund5UNOC0pu6ssXNT/5jOCLpupTvpEG4OsZaJ4Q6U
mOmGVVfrWOYVETj9ANMn7G+hzQC2L4GO7Nvu2J48Xsr6rd+jLwXLsklXm5eTLh33
dt7OJWipPZV32a8onYufFlkzaaCupTLQepXPu5nu9yk/xTgg0umeoyUjQmiIMQDi
/q3h+ujyvtaevOnJiki4qwM5SncVrWCb0E+HMV6FXclEOB7ni0snUASqn2QUbdEU
DdVyBQvKL6o0VKBZAOvLxKzTq9TCsw0HYlkpTA3KtsYIM7iikjwsckzb/E2cZf9D
IpiQj9lwm3Efn+fEDSYmduOqxyC47j0UzhO5pqnPK3Sn4pFpV/GWYWUhOOfsTnH+
rBK+gOW3VWgr9zgdOmuoyOxk1OdAFzmnF1eA5FLkMG01nu3YYz+hfVLfx60JWJhE
nUxpmXSiUIiPM5ns04p01kEzpvHIxF1HlcH7XVU/HvblmU2UMSDZTLoIvANc9Or0
6MQVfDoS4AKykBeW477heoLVVuxnXLYGSJSGrkei54jfqkHlahV/8IBzFHZhEyWa
SbPSCKNfqYJlUjIFiDSHqjzggB4nIKbmTOmN6h64b9bIMEMggFlNc5YI25nSfuog
yWKGxBU/XgL0SudKxD++7PzXL0BZWZxmdWW8O59vK2Wnv9xqV8cumF4AZvCtOXCt
s8YGdIHy+YRcoBKbVuATsI61ZDyhSjB2yyWiCLHCWtYtaapnnO/E0gUoz6QYE2ig
ptZo5BD3aCV3DjDHXOZLkE1DLS1VPu1DyGx9I4WSpPllDW7iRkFltGgk1a7JoYQ7
bDIj8Nf50baJwQZz2aZssuv05c/eDknZRlhW4J4l85CxPdJH6ysKhYK+1UqScXhO
YFLhZp5CMWO0Rv2kI2icERtw0EVAFXYdCfoOrJ4UdnRGTeapVPjTtNsFO7OFCNjg
J6srdfk0jayY3fOBn3auXZnYE3rppfjgZOPvkS98BDomLF7cLzRuVtM4BszEraze
ScK8h0z25Hu1RsbhGBI2xIThm5qiBRxaQTFuYIZPKbeGJoY7mx5mev9ZsVK9ICgS
Q8Ru8u51IPGtEoQMI9XrdvobzSS68R2Bc1nso4xUQetk7l4SZ1clFlTNNiqFbUEs
yvLsoRRA49oiv7DuLiiWk0khkS0Q541E6PYVP8G2QQZ94OdATDcL6y6XgOGcICeG
UdJrVknKcQCBo/hqd0dhdWRglGHLvVEAwlofgeneTaosn09EXaVon7nzue00wSWM
VMo/L0EH3bG7Fz/Oa7AjO3fDGd2hI+h9pGDD3LeF5IMNuExiT98mofUqgdml04Rl
Qx2ZWrVWj0mz5Ox8F9ccQuzPfuNIxtZsYzLNYpntmuh+HBRJvNAJl9BztaC3+9GV
MEqXvpkquL2qrOB92b/lWKNf8GVzUW2zOeekgth1POR4FxKfknNipK9pN9aKvcCy
37+yiEzKMHY8KjVogOxvyJZygyEsji9Rs1sFJF02UQ9bl8PkdYARuNLB5VWPcd34
Xxsy8NENF1AexHsHCndR4JPxtnKKfL2jB2F/QQRWEAnn715M9lRs3QwXFAcKZXnc
4ZU1hkPQYhL1abZtkH1aCoo1XMC+ZQA8oLn451TqiGKgiLiIDtO38uZgM/O5kd7E
6Ah0YYvgYytL3aGWgs72/4D4VE9eOo1jHTiwe4q7pMZKgXPII3tosZiKG6FcRWLk
rozIZgqyFddAgmuo0FJ7BzM+4gmLtIC8sJ5i0YrbRvv6k8V2CUrjJgh9vsoVrfMV
rbdtSy/TW4SaXcE8UHphhujRNuMEILw2xRiEaNieD9yzq+THsF3Xwurn/1CFTsuB
yZjY2CtQpzur/S7raO8HPo5kMCFyA78s2no50HyH8szSTN3nKpzXV4nqnQIDEqBK
saPjd5Ji6KPO1pnGD3XybdP8T2JzQUy5y0VBLBmPcws/4WmRqj8Bo1Jc7wJs2Ud3
WNov4Ofox13sJbSMUAKeEyXyvc6fipIOtVBbTFlCZuRdMD8vCmMjei54H/yPC3fn
PdTnJ4klzmowhXNjD0057Gw6S5FxdXtCfmVRNHIZLgYqI86pLlGoxTvTPMya6Q1I
y8s2sHC1fw0sR+IJtm8Dh07PoolJPZ69elCO2xareSw2qTXpdLU+xFd772AsWdJD
Phi3SlzfvKpfUDcYo/81SLicOx+KePYLVgt8l2P1ljmBXC1Ot0RHUz5SFCUG+Rg6
xnlctzgxmtHLeQpK6LtLfGxsQM5b36HSPYD5tRu90KPw/uBYg8cgbblZFCIBCO7Z
yQafJcKO+PARH7wTHd3l5FSJakSu77qQ2+zQeGDO59DxlFX7tCR0MWyS/QTja18n
GkMSzWt4vo2DLLiYPhlLCcAUDLO06ob5PmQyTB+xDwWA2hfaVW0Pzav+k8wdfcoc
5Kh8LUzdbVmNvgzQXRUhDykkii1esH/EqWS0Zd+VjK2blrPt/Qc3bMo0ltwr8GEc
v8CsfBxULS9Tf27BX73Ybd0FIBlu8E1V3q9F+H1DQljs4VOrAJiJtZoLdhtV85+6
XBd3cXIlfrulxVL1ch2FXTY5eR/n0sVOUlpDwtiz0MqQtpVOW+Ec6qGqebDz3ffp
vgOJbjYzFo9Tfyf04CDywQDsUFtasdFUkkjmJgqRdq0D3ri5hJT5J1U5GcXLLKyM
Y/xHzDhcLqYZVPuFxEaLJEHCbLi5BADs4X8Xw+FFg2CpBxScUD1gbwvWfFn5bVjo
y52s0oEE3/v58UgZIYSUku5yA0zlJe7Pz8voPd8x9TMrWHUfWXH1LpotNMSX7P+Z
258wpAEkZPnXsGBwhySZ7VEHNIA85lL53GgksVwBTV3+AvD5YxF4J/Y2K451qufZ
iT/+sMAuK0u9u2/E1OjPdPUHodhmiQw1o6wXcCFS463YpNGP1gjfl7ONyy/fAc5N
/NH2FysGeja5T0nD7QyxOBAl66fre77FONyQ+lQf4ZOBboYyr7mrfpyUDcbE4KF+
jtnRcB2xPTJcZgQkVkRp20H92ZOs38TlF+a3dPmDeEWHvwa+IoGFhWpxm9u+fSDg
jvE8ZCGsRNl8/PUcIqZqEIb/O/zq2juDcAFCzBGoZqOypnlSwtfUAMJMZeWzvkxU
ulksXqQRUyhMTNqnvc0c7cbfTVJdfBODWIqPCKUa8aBVdvQ7MJRR9in9uXtLJRa9
tL1rQi+KUdj4F7x1tZCslnrPg/qEu675ppFUaD15DE+uHDJVg0VxZ21x0Z1RgrRI
VepH697MQRFCD42hPWa8lgnHRS4Ifbgs+SmChalEYx356NP+veQeY6VbmpPxsq77
PvoGHWvkmsFBgwQF5uvpOPdmxBCiuftOEIk6TIyD32Bh3zuSgA0C1j21U36xSGf9
DR2Wko/Pi5Nf9h/o1q+LcuRCK3M2UGThNftBOhAUxdE+DlbWSqezpvMt2XctYF/v
hjmluoKbYcBvnGFN3xx46i32lMA3VumxAkjgr0LjNXzSqDKJKJ3btoYBRz9W8/nD
syI4GPdz6ZlgfEALSya72qhX2nbdj76d+VS5AkAzWny8sWXMU5YDi/vHVDh5B2Sy
YdFTpYiGlitpylMMRR/CeQRqpfXq6WMWEEers59R6VMWqz8eR+lw2H+vxk1fR3cr
PSX8lm6nJrhSvbTeFsD8OohBUyDY0iFCSYoYJ6gAZu90gUGfVh2JnFpkWkPKlbt9
W/ln22XIl47qkcp76p3ZgYsYsYjPaJzQhAQtHj6I1J56tcGL7isVp9dyMk2MR9fP
r7zXwuAVt1cS5Za9Y9duYkMW50OX9syc7V+Zu2eN1VjTbGin+pTqHRKUGBVBh/zT
lLqp1Rxbr97esx45C832NkXyJc9QpwZl9dZSy+ZtyOGzCIPfAJD5/CNEu4mSNWch
yYevTMnpkFoh445cDskqaS4I4HV5Yy6TXYbsNQBKElRGF+Hrps57wQ9jtYu3Vssp
/CByyZyOm7rTWO/1W/kp2WmdIEt5j1e4LTRmJGHgJ+mWtbH8Xl9x+Ih6AvLwpzvn
aKsKXb3uhd1rnugi9u4lob0cl8Eb+4ubJ5+InP2L8Fmf5whh9IpZf34CAkNfM4H2
mSLNfk3JwQfip15v2E8T/JXmZXuKWrdtsLGcSkQLs1qeUeY2dM19uJuOq4aCa3ve
w/231wDKzT1E6jraKhdowiuyjqnONpoE2xympucG8dcYkjnr0vNbdfvJ/eo1OERI
4KUSX6IFB1FnbAXIdSkKrHksoguHZ4sHNnkooVMtt0qwfbLc+/tt04B/g0T1aI8A
qTDF2L9WjZapaazhM6p1IF0ZCAI7ysqtKHDqBbAVuNA1Cu7xtUnjl6M9v+hH/BzE
VxRGnqnzGLvy5mbsEdbFuM3vpo0wf3b5Q125xKDTUyFSS4VbSjpl2paDamCmLedi
NZBPgMBjmxtX7+/KUFGsiUxCmj+ciEvv6pvMeIWgwS+sLbc3OtcxHfNR4ewvzYwH
c59hyB1Hbt/VQBmcgz+CKZDMckcY1HNeWiZIbitArlnnWcWudev2FOT5CBn+3w1V
JlZ/m9c83PGCHc/aFaBYYnafyDu+JRGpOMH1PzUAZF01DJrhOdUd2pusMJ0Du4iT
Z+wiNNjNa6joLvZTflC0zp4RDxHseqQrBHm0kA18KttdiO7itYEasGqEhY3ShJN1
UgydRZSlM04CDK8oLr1zLJ5Kpv9V/5aLRQV/Ynj0B4wZf24d2+Kqn4MthuvFeaSN
NQen1d/osyGI0l7mpKGkGgO3c55MPE7zDEYmBLRDSf7Hmr9Cpbr69jZxF6cvwt9F
PlUqy1VajN8kQaBI1kXKBKzROscNLO4ODnid2dAzakYWOB57DW9uMRsAVzHVXS3v
Gc9oyuS9ped5YdJcEidylwJ3uIg6+KcQ4cnd8OsLF+rnI2NPxFgYpn46x9LpgVdp
pkvgANaRjZTFEjdVXOoT6AIOybzwMri88r02FE9A2dwNyWXxcHa4Xuj2EBpGKilp
nEKXK9cT1Iqg5l9WjvhWGIXad6yrJxqtCPYUEAz6ZwiJeqlNhB1gvcTYqlpc9NFu
QG6oj34l79EBaqWeTWT3iYYlAOcJjNzFDBA70jpCG3Pgef2SAJ/HuBkBfCrt6lJL
txSwXznDTQLkISMZIEQsVSRX5uwfPTH7HbM866rRD14tKxdSIkc7gHU1NHfFuVCR
EUukedfNw7jlzO0YYA4BhD7JRYi/Dqj3NKFEiT1qfe6pqqmAr3KPL32Im+gjnzsW
qTukkfyXrtfdr8dZ+szT9VFgn6pt8DGn8F3fQEupM7vDorcDMviVKR6TRVykpgdT
CAj1Y1Kf3ATg3JuvY2otTLAdXgOR5sEFGxNoGmomZ4mVMv0ME4tyylu6KcaCivpD
EqIM1KevmYpTrtWMms487wzVpLkxNyvd9hUc0esMeqyeyf3hCamgaQHfzBAMMws7
YtgboK5VJwVTQ36akcRiF7SOrrxckVR1AZNPCknJ7WN8oPH/9ZudKL304WpTUZP3
sM1vLLc1UIjh10vFP3HVKZHa7t1KEt9sK1vBjceDuSgBwoIkRgUwDhYgN7eLPw91
Zkt+EuOC2Gb6B2OXJEoNveHHNasDzmwtu9fzl/vl+mDsiHjFKxx7PZG1YxEAG6bv
VXfdk9djsjGcH7TJCrW6L6+isbOqb1mR/WEicAdDZtxKIet+UuSSpQZBhMktkUEF
Od9+JtSqxSPUSsZ5B94v3KCiRVa1cyxatpEV5Pp26r/VWcbzcg9NHlYX4qwRj7FW
PkVJWmdSdxPYQYDqFz1dD2NnOfxa6tCN+XskkuCt7gtn6PN7Jua7L/MsWFXvvEM4
dmSa6DgnA3wYrAhFjk7Ben8wy5biYgCBTez+uQlb2yWfEyLKLG4HuRJHtb++XjCQ
9AWX1Xpac1WwEbcCvno78Jdskh2WU25FN6T8ptEBqgI4cZHZ5xVg7WSVgZ66CrGs
q5+UDQdfyzG5N40f120x6AoNWCt1au5rZGx2UFWP2HJiYmXU9sFX4ADpGLgjeZcZ
SFO1zibaOMTIWSEKcRJj63X8uHf97hs9d/10yieOb3WXc9unnE5h8ZGX6wn4x2wj
oLMMlP9v15rJSfRs6z3IsHnhtM9kS1UxOgZAp9TqoT9Sza2kaFXIncOWSMPT/LNJ
NV1pDp6jQwIJ/lq4k2K1UlAhgVGEdkdqyAIsTCMY0ycsk/AcrY4pxGn91I4oj99/
cEtAU12/yFo9/eDfQAbg2udVhY5mdidLheqZlRMauTsCprtHrEeIjszIgjP57FPb
Blb1wb8F89CJMjphT1vbI//xlKtHKTHLLglE+tRA4A32BTEG+muRBoHNdZHog82Z
+1djt4WcMm18mHGYypwKWQMfKP/kVCPgbK6hxfAHFpZxTANh9wqH5VEDDjAmf1eH
goAKBwxXnulC0Wgd1pyjXKPYh3UKVXI1SVODsQGKkG+oEExrV9s2KhEWXd2QnjoU
QiMBSTLXTO4imbAA8YUUUp3EE9f+cZuYMkYTlm7m1xetj9iDjZt62KKAps5wFl4z
fvFTzRWrYCo/SZtRoAxungL0VOOi0L/Dj2FLezVCLeXYiLOOGzur7PFtHFdncrVb
QasqNcduiFdJ5eXYb6XpNPAEWx9RveBI9O5lauUi4wAgz0NhIeYJqqH8hyegmbwr
1q6r9AkHudXbCHhB6YNzJE/uuc5SXBERDCgNr7z5qf0g7MKOgO+Tc/wCOClMe5Lf
UooeJ70LojEnWBSwvSR6AtgVuC+gN+OoecxlC/gOjHiaezkKQ80htwETI4fVfXg/
Y4lfx9wBEQ6USSrIzp14awOLwQ3nC6HeorxEP/8cM02tO0AVM3Fg7xnBouCXlmLF
mYuO+IYvvdalNWsS5JAxvo2leyLebtAC8D+HhsDoXCNd/b1uK0P91bKs2O/JA2EU
yPLyEDKMdjxrp3Y3Y/+9MJfkrQgCSoiINYxdA3bbL5EHH+B6IujIBIBFf0TmxSFO
OBAES0FGCNSJjhOF9a0fR5Ael9d4d5a7ZGHmOfltBIwYu4uWNwFmPuZA9iibuzlE
GJe2EL27W0REN26MF8WqjG22bEKTvHwSpuZCoOWEdce8JKjmkSdyrCjR5vm8D6NK
ZUoMdvCogTZWwMaGzmXffeUaJ75P2Nl7tZlJJoca5JAWHLigPjkMMK+mNfNtieAg
i3Q4CxEPdw12W+IOrPfYMYpAWsYE03JAmcIZQUK2J6elIAjBYWJzng+/dhE8dITR
ynhHEUfx7dZUDcx2MnQRPSgKJBwGJ35N/jmiK053UjTokLNPRlPlq+6eR4mmwEv4
TF7djyllbjp6VQiiQBG97FXX1ZlJEMn8tVLTaRq/vxi/o1+4FEo306NmJ2XKpS3o
jMi6Ha7B/B6Na/7Rw0YlewNaaKr/2zUk1AYDtQ/5nOGPf8eufV1Y6K8+tHFYdEod
KqlAnFowo8lqxG2Bk+y2azapsrM8zIuBvw3le3SRC56m79LjmXuefS0X1+7UI1IW
KMJTZx0azsh44ntAjKQ6KPnlEYXC0F3ksWPnZUByOxp0pLZ3KN+p92df2NOzz+oZ
DL4eLYdcoGNf0ngbzTVuSw2mC8J0y5LaNeOdrjZxRhX8lPxPmB6G7WyNKJJ+NMwh
Xw5vrnfwLLL2LXsfr5pXV9IHp7ewhhhi1XOghDMyivV858dBQ7Zz7iRy7SA2LaCQ
O+T55PtyeKaobizHHz0AuzeGUZjdh2ys/mmsVL0FtuWHWHqibAChUNpqtvFQqYxC
uknJSdezhoYm7N+jKABgbx7J4Mox4om8pmmR09VY5w/FKHe38N5Ioknjq9OS69s9
MbegZ7AE5OuMIjk5AGfvXHWbdHIKVIhym5LdnEDlM7Ir6bA7jYdMyMGA72UbfCUY
UYwMl3xUQTBT0EOG3ffM6U78zt3FSMsjRkkq4z+OqtRrhVKwfmipAQrE835CGt6X
B3Co5OMu8hAVHQlxViL7pleCOdWCYwRBaBQWBurQACtoEPHgca8JnnfWW95TQtR3
LqLkcBWmTq3T/Z0PREBYvQQXP8/cgCh+yCgtfaHgUqgwKSr9VNiWH/5uVN1Jr+r2
qPhzStZn4Ft/ZjhMEJVmKPZElGTyIs3fsLytRBPj3n69EwPBBLMJ7P4kwoH1r4n5
H48oCoDdIuDa2k6tLG5sB00U52o0G/stCY6TOO/2SYMKp+RjtrPW2AZACY5a48fd
Q0XncMj80EP0jS1TFXLAG/vHFXqCKyH8Js4yACm+hCE6RJ7ZZUiogcSMoUNgo5sQ
vUyPVXUo03dVZxJt0fvx3wJcKNQtvjOgfkw2CLZFowCUKaKxYe/THYub7mv0g6Nz
kvxe/woocSXLPyZPCo+WwmntQn7BZXpWK8Q/tx2GPPdYJzi8INH3rzEFWXvTiFuG
spgjv8ubZ6bn7Q6308sliypuG245p8JQs6zCdryE3bnHacAT/VJJC9z06A0CqDb/
JptM5am+uvrGH10zEkTnHFyk4/laGyN7cnl5PTie2I3Fr+pDrkEySaw0akcwqbRu
ztXPPcR8vKWOFngJGw//VMVXpzrOoTc6nIabue4VK7/PNmGRhg9dFhulaIeakyi/
3bnE/i7acXoDlL8L9eyhPykJ4NFs0iMHWWdYQPlkvXcyigaAxdqNXLv7qMnVuJaA
8//CdiyVyPG4v+nDfBRwbv57TPAf9a8ylhCatJnb3bC007B/w2WbZdSEt0GVVIBY
feUW2w56nk8IvlxaFNQyRvYtM+OKOagZHZGzfiCvaWf/DswnmcVNkJXi09q4gWvI
rk2BAQUwksLWx84A7t30FJVOLc20TtXCOgsJhdOpYdo3FSahKrydWm2o6nlWOtWJ
qbmaMnaRKzgycQKy0pCBXtDXdALnqQbf/qI87oO+AyGNdrQqcDPPogKH9ic9UDof
o5MskDz5q+EnNPndpwBXodxozJkXTFPeNjUUiOZtn9bPIpqe7zr+DG0zZGEU2A29
v5zlrK3xJLcqFpeB3ghyIrfD3V7F8kbAM0kmg0bF7p/jZ+Tbs1Bu2uHsk62YRI5x
yB8hgJq4+ZbJvt420jfLacduPrtKIsMqHhrr6nEzBDplLcL5FvHISg6hNWM0OHSJ
wYWnr6pfpdY8SgFEgAPeo/LKfUBiem7mwm2KDRMGP3wsbD76akZHxvV79pdNNU+y
zITaWLTMA58UmwMWQ82ks0ixLXQ79aVZN57Tjxc2/MXcyLPh9UWo6XyXU5QqRDBy
sn565ef9/OlXEEfAwP46ZunUrkzQdUFOHcQdpG4RaBXERZlbrd2CaV3gSAuQn7eW
pgfz+P/sAS8r4LwUpndl426si1IAjdtMi9R3ChkjiVch+HFJH0MCSDUCCu5i0eLy
FkJAglHT8Q/BTF89m30mMd/4TXYvZoh+ps4oWfLyoPPDUtbLG2JcTeyWWAuM/2gm
z0X/achXTtQdXVPlIEeRZOTk/Khy/Cpc5Squr0bOMyXjxZJtm8rCVkWhSBKki1nW
1YTVSlHTLASYa6y1H5BMYom9vhoagdei/SWYlwL7gi51UwmksjX1Y01N37EDWP8B
Vp487EfLA4biDgSiJDFz4vIWlQcPOP7aegXS3jbviytcJ56mizwu/M1wsr9z+qN/
z2L87QaOyezLgiw7t1EeK+zzHmXFk+d6U+rcmL9vw3PA2pkQzXIIq5AN6v7l9YQm
dGB5ePl7Eqz++bUhBJU+CVEzeNeEFPJLeYg7zNTm9KmL2I89ekI3W+mYfP1B4X7A
Wn8F0k/J0V8rcTA5b6fQZ3FsWZJYttoz9G/qGOiNLZzjayAvsb5vAgOF4jqYxnOq
t0DGlhSjHAogHx9NwML78O8pV8BjDAjub5isoJGIli2CLXTu+z81qqeTdFk4WY/3
jVR1zdXP8sXywLsRmrIqCIuUOl96eh1ePmP96tWJideQLB/dO0Tnl2LWUMv93hb0
0AmzN9z3Y2Ep3d0reJDgOyHMl67lluBoQ31qZ31eIT6x5V/hzHL0rxthc599yFJm
C7t1PK2zU/6J1+8wmy06GSWaUgpFl3LLwsJvf3GtB3+JvW3US/gfCn0E3nIIc2nH
B+PepbIofZhZZEuB7sAk11fzYZS0hYTKa5/UDPvvzvNTqFY1lhhWcg9tqp8VEdBK
LpW6lxvLRvmfAoHiFMrLwaxP/ltfwkhbzMoOCLTKpZQeEurnqjy63mlwxvGwddGM
5Y2HuF8rzX5Gc7jQY52u2ND9PduqxVrgBu7QUHGgJa6BHboaKtDGmtHa5dIT+hXp
PJSDAaviPiuMb4hgVQZI+lFn6IC/af12czdxcNzPLCVGsf1/tmLF+nrH3yWaXhpk
knm26cfp/LD30boAHjvFNilsd7VLtEn7m1ru2myzptAEfpH/HQzo/Y8DcLDBm1Oj
i/SXXSlcqV+f/tVJnXPAlZDw0w4ycfO8GJlYbDAjyL8Nhg7ZWXoSoyhqzIfX7rhV
TOMSsATCJayyUfLr6PucPFlpmn/kK0AUYK6XRCUo1NFB42lmc8pKhb8EgMmYBFsd
fHwEs+KpzWstSJtxYPBFZF63Dg6EjLr1H0Bzstg6r7uFPYR7FQUfgNtQ/1oOIDrZ
SgI6S+qgk4l8ZrLb0GanDZiGXpf4te9BsI56k/HW0neaQ+8XlZm8PAyiHaN3U25i
tMtOYHBOerRzhEJxveHMp//bbMMIU3a7jXLqs7thW42aaFvGiVM4vwqDjYgsGLrc
LrjTRATfud0AojhAdmJcRnDJhgLfLN1jg5fgwLTVbYALJxTFX5VGIEkHZyRB27cS
0IBvhMxDfwfGXouXnN6wrT6NGdmEQqAnJc/QOtfT8gRRTPq9uLjl06YSuJagVKIT
MA1f0EZise6sKYJG1S1x0pjiarsSeQ9AAr7rRTv0ax9+efSd36coR5ZolovvIePk
4Xkp+D2+OXqQNL6lwRp6x1tyQ1S5zJOQ3I6gqEauR+uBmKGdih/EjrfPjGd0mU1q
iv38ji9yH3QOqAR09J31VQsTTT8v9aHY35fd8l86eXl4Ds/j9lsAl1vEBsNIgMAS
0tC6W/2MNPNtIs681lSLqQLEtth0Hb+P5VLZUWb5NZnlnlq5Xl0FyGN1rpCAO8LX
lMlmYnERpODCKH3HPrFZH+Or9Ne5Kc4AXsUNb4FNn6+ZKVvruxDJkok3t5bOsIEO
Wf5tOvx1acvTSIQX9N6CSPoM6Sfn28l3Nj3pCovR9Zikb6eW773yaPrIc6cmQdIX
f8CWk/bFt+kiRQNi3rwRWYIae7G8rZi0FsadAMwO6Nojr25/h6dCQ+5izMOtOpMQ
/k9QuPgPCYsNsRl1zyA/YgIhBQUPRM0GoOcTFZpQI20rVWKgvRsZ21FGqEcgvoxD
VJR4YqaKUTfvpTjrXWheFgzBO0b2OBtF1oXkXmM67vxNiGsqRdeSjcDSzGH8jlZ4
1wNsGrL+e0WSOjOEApIyPQOyGIKamTlZXmEZnZwfQ/Br8tkYy51Y1TXVJFnbW4TD
4ndKfPu37aEDxU2OvE5RxP35S7o+eLNHm+YPIQvf7uq3itQD0wR6oYIowvjnVR3p
Fd4vDffhjxAaAeA7AY5zJELRhr8AZmZFHQFr8hBpbPvvrKFyyaWQJArk6sOPckbs
LVkEX7k5BqJSnmOz4dyXWQn1deGeEKl5cwkuifk3yUbxxMHC2IVcDGb5Xn5jYCMu
C+mnds4xoVz0SM6hqYlBiw2v0ZHl9tcBn+lyePSTPR5I9W8s8fxEzoPa7JKjsstb
VdQ2G2haAmpI3krhgqM3q3dvUjc80Ogc4qjdQjYQ6BX2EVMFPTsc9x0knXbfXQ7m
lGEXSuZobqytjaF4c7O0ctOS/eYK4D0ZNxdKTXmb9vUaFOdl0kkOuB/RVSADnaqD
/CCpzTzsc3oppRvL2RR/YrYvqzw0XhtPVTdfAwUQBCgLyB80XsJsS22pkMt5FziH
BOcvv9kKL7k/S8mUQXchotSU9VO3Ex2SWAEPXQdMmCU0SJbgB3VH88qm+TyUNEX8
Tm6BEbUDn3PL551LQPqfiMmS39h1msAcZ8WFismrglr0SevM530Hy+RzT2lEzpBp
qFRNBJXnv0jCMHvFMd5eFKRDWRfgl/ikSQRJ5euQIzmorhQKobr1uFDrodbrbJvG
ftuLM0WwUU7RTa/+vOX0XwaPvhLX8B8ka8KHkZu6FVyLxqfGS6co9OI3o7SjpMsg
6lv+fhFcCIZ+bct9oqTfP9B8Z8A2a7pJuflKw8L4bMBHpMnn7Yoy5pRqQtHGhLrb
397WeLiblsl+sX08tsEa/SHyUaJ0oSVguCq788fZZUdyotyqvWjWHCiz9anggGyL
ZWOsqKF4C4veTBVqDR1QfSols+FQr7Q5oEiSG4rNlai48IC9XceSpNabVTnXQu3D
G5Jpa98dSkB8qLZHTBDW1gc9m6JaXWKjpVSPOz1hcseQYQGTRt6/WlIXprBpX79s
3D4OhJKrdu3RRw3jUCbX8fdcSvS64sKIvFzUbkswKKPdNcbqDgpTQ788ywiINXr5
mZYOn/Br0n7iw8cJRxAOQQ/l/8T3pNoU6rLsuki7HA1WY4miu9iPMzG1lbXwcpAJ
tdjqQfKlM+5mZHQ9GA0hbbf+TxZrrwL90PNYy+flUNGsF2wmKCt38ayJA6dCUUmX
A6TyOnEe1eUB9GTgtv+ANet2xn1rQ+ItZynCmZNyaI1BKrVb149YZTxhvPzBT/NB
e8oEVEyDIjR+Wwq3VLM8hV1UJlRuJpg0rZxxOtvGM7Z/U6VRJXn14SltK172uOh1
7ubI4ojoIcLK0w2PR1KNkyoYZpCtetu8SN3GXMUam1lAIE1gOsJyR92+dwaYwzDU
XKet2PUYserlLZEiXwDe52NSHGcQiSXZtsnt6rEn3X8A2pzA2u47AsEtBT6iHI8y
X+yEw96JFcgXKNlbBugs0PN5b4gfyvdeVjgpR470L/z/LEok1JyOl0gDf+1nxu6z
9ggaqyu4koNKfvxchEU5rN2u/vsZmMB7W0T3K0DjyE8Fq0+RED2S9s207tC2r9dt
AZB0Aq35JOk7M1lF+3ICMLrjHeSYWaoRr2VYWrUcZNY+RcmkeBLBbyQSQLbB4GTm
N8JaYZMSNZHEbuOddwwUew0OKurr6RljwIz+s5+NJfzMiOVMZSjY/THa3LaEnJu+
NdnxY42NPwTtng3bXBaQI/O7wcwDltP6q9F1FvYdeUdPpnsXh7BFGf67tdD/ZwQG
StLrT1ApD36vKLyFqcdmMpZtvw+oqYEmnpxGFEGsZ9lNgXXmlJcrilvx7b8wCV+B
c5sWnRi3tubaUZXzCOl+mXu0lY6Ew0cUPN4EATVG60IsKoLf9xRphTZudxB/hdH2
iH0zKfxsbKVMlpl4b8kkvIhZWfaUHwySfFsSoOyZrkbtQuTPA/J279DbjIrR+Pia
HKMD036MvV/+942xtjMwSz7DbYHzUZokGguKwBAvQj1ahkYBe1sQOj1zKatqHU5b
5nsgzYOUTgZrJwLlj7rlvARW57iVeXXS7LNEH1+ejKF/2XDWLIol9W0Bew91jQku
mNEisMleASpFrWxCV6R53uQebL59kSZDcFVLTQfruaUNknZRzhgz1bk3ppVWj5zZ
scm2gSBCbNSfB36BDxdtt/zxHkj+zcyWPHj9APyuHKPUSS0ajxDxIntCvVQufmlj
jp6Prz/cTiMXr0W/k/59R+ulJnNPboHQYbDyz5eTsTlWhy0ySUcRvLdiLat2dxS1
I88GFAWkP3fWDrOFbWz65cqd3r19x/Pzchs/sBAtOGN/Tx2WnPtvwMThV8Mb7eB/
2Nz0NOrYj1j7sdfUWdjh6QNkT24nS8yyvzFsdFmnq2ZXMWXgXplZhbcu7GC9d/lM
7liIkrKrLSBcyNrgbTulyxqjLj4GkDHB8u91s9HYABasQbcfmpB6jvjgksH9vIt1
0fQDyXM6dWeHEdO4oSRrw/1rc+LDiDvUUbiN4lrwScMJaKlSJbxPL9bvLn7MCc9D
HzLvDLu+LEFmuLVVZe/E6MgWO+XLY/PTm5khnaYjDfc/TzWB8gIsJlXqJasePxVk
8UDdVvpYvrtKZz5rMv5WwmFjfaYXJFmgrfes0TEPhMQOFufCVuV3athw6F84UArn
djP6EHpn8TEnsrQGEbByOWzKHz3uhdv0pr/Utyou/7DHSmHJ/NqKyIRLcCb6qQA+
IIJRUlMj2zihPiWJjK81euF3Ts3UFVGMowP6zMQMZJZ3hHHFbNvhnW6+T80R++XX
gZIzofE2FfXbFeIVrb7h3niGOL4FAVM9DpmGnp8WT5WgpkRkihspSIo6DYeKCsbC
BGwkPj7CXi+NrJVu86laRJ+ben/xOHNHShK0k1t5ISdxo/T0zFg7bMIBcp8o8lf1
n6jLGQ7c78/UheOvH69s1n7c28Kqy0Ulqyw/+snntF6SEiblCbDpUrdnRx6MoyjP
zE2PkwTd2/bAxeLIFi1rR3p8jw8QusHoBpzDjkGdSZDHgMWvzOvu29d8I/ONK6cj
vkTi6GtCbL4ZBhmvrSHXgNrJXPqwEws/Djm1MX1Ewrtk3YyTcDDipRG9TaGHf8KN
WMjkuFeW5puKwK7fu5HE7K/rBe7s+98/AZuZ/EPXbeCz0CEGHH9Kz8fqFCjmd2GL
wZ3eOuIWocZrkwehU0xPkncHME8mRFqVcXjrtL+IjZUpLUQLKVRvmQZrJ3sgmohh
xiIgi+cyq2VnodKFfMPtO9Lm5eLtUk8O+Fvy0XRSPIlnwRzf/4jKeD3iZgR+NJ9K
/j6zNfE6/pgddeSRpv4Dl0rEV0WbPWbapdk6nO/U+4iOouZWQ1Fr0TKjs/mQ8tiO
dKEM6foNtnnm7mbDNvVAX7RzTu4nnVTEGCN9Gs8JMkHUWXemi1Yw0jWSIMV9YvS9
4R51t7z7Bob3WjsgDOYxKQoapT3tU7qF3Bj6SWpnNJxGXhXOP6CcQI9dBO2hZ5BA
klizdh+hIk+X62ye5yrHg+s30C50QL/b5T1/OxqbZAYyCfHcsvAV09zxpprHvwRf
xoPrn3hRNf7oMUPkbRvxRzr4e0kEva8yr7CcxZZDqwTVJymq3eZtKzwOF+GGnqH2
ElrAEIYUrSx0T5Dnt3DtybJ/L75cL3mvcCeFjDUnw2hfZ7NPuOBKW2Gu//McP7nX
fBnV2nkf3ULrg7mO8b6k/qDFgMpSapMfSPoZDG+HCool90uqBIVUV3qxTdqpJk4e
LW1IZUuDJqFYcXUdKNcPoXnOKLqP19aScKk3B+XNNZ5IKFMq5atur9cKkug7GWJj
4qb3W96SJLd2NQWoV1eBdyRfZLvr9bVeMG/n88OhkKHpOv7GDCwGMHw00SYyYnYF
MpOlyM4UgM9LLq7AYERk01c8Aj2LomW6RZOIXcEEv51qjtA5Fr5LueXYuAqMfcNl
9HQ6kibez82FauFllnA57765e9oie73cwHJ54cjmoykNaywfxFhbQD5KlFbY2LMf
sqZH5vgH0vOTFTBethvpi734zGNcfiJaH20Aa0Tqn3y6WGyk/UkmG5gTOe3RJW9L
uOGBVM+TyavL5gWNEdUArYg/DV6v/bQrkqzc5DXRW3EX2ubRl6m884XUtonTJIMM
LgX+IMFuGCc0xnvQgARGZFnf2SIxrlyQ922Rx0XWEaPygf1nE549rxwkveeYPUi2
SWy8ACJy/t1jtgLaIZI1uh2o5U5741SgSGm46RE9ztPyAesle3sNv8UQuMNHKJu8
+HxtK18wSaOpCJJ4QVBgyOeSd6tpXLq/nQczAFdoPmjjqydXNrKalX/xTArgQ9Fq
vtBxKVlz8SPspxj5xFh3Bdcx2B0eLoq48GqlBHu08Y6moutCvXN+GmrWAc/QK9lf
hgzk1VlBx0dsa88B61HoBQEwI9MEbMrAJEXzjSAuZzdbI9r7R454pDcBNKAWuL8N
7ZIfcYzNYM9rBVUq6Or/gDUG3C04nwXpuQAdt28jzic5xheoAtkeLpxFsnF7L78g
MssBbobCEBbKb+am3JaJtKtKk2yFyCGX+n4NRNsCUFjY3z19rdq+wNHY5+8K5Zkg
pW1Soai1u0ksLjOXemUmX8cldCNCa4XjboKUmRsqBgk6+Jx/dUq2t6oFM9TYQB+P
sw1lSj7HcdqIIJ6zJjIR5F0TnHhXfMMW8D0F05t+99QX3nuVlDqblP9DtKq3LhRI
cZICJTg23nku4yV2t5STyANpg9y5p1Hst0IjWjJKlZGCycAOgiIAg0+4RVGObmn1
O2sqesUqFeavHHpqeL6a0Dyv0GogVSnR4oD1PVf0V0eg+U7oHC5LpaSr/8hpFtLq
2s56E0Bm6MOPZN6rrx6R7i06gWMisLQSgKBkYleJYhvkEgEQwTWK/mTsh1Fkt+yh
AdYtWKFOV5iDFVYCuzKzycZtccnGrhkL9WXIrY7+v4YRTDhivnWh/Y8Lxfup/x2V
xFxK9B9tC4dfWOuW6qppHohlkSsdrjflKrJwfB2+2QYLtH8X5Tl9SvX7x0CMD9P9
9HT8zKKGs2srcxT1O+pNZWPt0IkQ+gUcErQ+B3B25lZyFdfQO1YYfi1GpeknKKb6
zsX0BqHuKFqciKoZGOVwIyXytu1i/VZsmCpldzS5ZromDg+X1vWU9aE2W3gPvkVf
UBxHU1hH6gTzyQWi67xo6hHkl/mhd04Tz+lakzEvG+D4PYV1TY6cgRvsk1mWL5HS
IFUIwL4ZyCa//vFVhWG5+MM3ydQL2RXuUjETBV7G1eG/lgmbAa1pOpCjyjU6i8OW
0pfpu6+zDjuIh1I8Ws8C7wk9FIfE7LeJ+44GmTutTXkKbgH8qH8kdNWLTZkmZMIJ
P2VwmvlL8+ygV8Cbi3Y5+TQwwYnFoiC/eY0w2ndwEBh0ffMIWTTwLT1htp5VnqVx
Do5Og0sto7nAC/dTi0od+589h2KeD418/v/pwocURMP+1KTrU0NwzHmUqYLFMhiC
jx1Xa/dwIgZV6Kx2Ib22USiCimdBtJtgoAP7+3LC0rZPDmyKn2NECwAbWLVqm4Qa
91CFuWDE2CBjG3BBq1iL9NC3mvxcold/lNXrAYdmQEkKWKgqRuALDRznLFoG8egF
Okm9u2aDOguHzeSK0UCiBAW9yBmrNeDLnagDol30/Z6w9V4sHwG2wyy6fKdauvgZ
bMls7S3pFINlcwdlzZQzgoimQaW7SavV6BHIh4FWXEAI4NF7Wr3QqvRoJg+rMrp4
gHE4eLJPt4Dts+DUjoEWE5CXKtYoVc22BpoKc6u3o6NWPZTLTPics8A+zayjGv3Y
W5bZjQ9nYORWRZnG+3KcBMumW2zuBDd/flSTU49l3RSY++JBB/mro+nqsTeBRu/x
N/iLwxU2hep54MrswQKrto7krygQfajy2gUpKeo0ASVDCtfyGmEuw0foilmwlLYy
eNegYts/UlUHh/kCK3w04BK7xSVDcyWAlNi72YwrBcLuOshovqaHyE1fu0Gb0Ouc
jRufa0kB9fwBE+C2S+48MQX1+VoNVR3qSR3aKaH+7zMC3hVJGrfLCNpNp8bMqSrc
PanBD77UaTFnP2GmfU3spZ4P8aOSSO1gM/pHvEsq/EAG3nShpOsdTdYH6tx+cXBi
XB7hKXNZx7viJMqOmfKwKqu9zwcOebIsG7RnuK0flSJN89kzIlTaVki4K6xWl7aa
79fBSjcxJSzOi9XOAvmgGbRJhd1RVLcekUgRjpzjDkptsR2OeLQ4bS07aHJqJ4xy
CRv0QgSkh1iF8dFcXtQoxeGuvXg6Z7G9JYybJmbszBLSNqyrS6/2EHXxEyfZpiPb
qyWKQTUSKY/b0ESIfTByaT6cF36uCrUW5R2KIukaZz/XXww9z8M/gRU8YuH2KO8q
F4kHzi/x5WV45kCmDMsYv1V81RiXBc98dHaXYvbRMtTm0ZmdQH+Q8J0PC1mIGB87
vgjrP5ZKtp5Y7i4frs/AIW3U9ea+i1bovi8lhh1k6+DYStGnHR5+0CLZGTiBqX4M
gaN4kkiSxk747aKya5gx9epwLbhS1CV8uPSxeBJy5rmEwxfn8pgMcdN8mhy8tNZQ
7PL3RcMplIoYJNp39Edm/prK/UJrthXU1R4NBRk7asOhqgEGXgGt0i36EoMv2JZA
OS4KzlCp2f0Y+p1jQw3S+/oS9LueM89tmwGSLY0tXXt4+0Y6wwd/3f39dhdzAXN+
wM5BxjfoTqPhRUVEtCEKAMEhBdGksy+Rb9sZVplYemXYPxskP69ISbXXeO3vjgnN
`protect END_PROTECTED
