`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3WM00ov1wMQkriqjSaAt5vUzTtpy/mzCJywu8oHW2H/i8C50/d0akJwMmxno7i8b
bQ/WNqaLLIHPkMTe6Sv5pr6n6fFxqFneAZyGU4r6d74YqIK+tnEfvy4Zkn+Ihi5V
ZDa3rKG59RzA3nPqpD9PRQoyZcow2LC4BgezbcdOsXZHTrKEuXY95+MkC+U7KWUO
3dJwJhlJaVbvtQoH1pWhYAv2U58nfTRbQiUU5qWJt3NVjtKfCbtkmrDVKmoqKyRu
FkY0La9ZUaf0nsRALkBm3bD8p/tit5F2d0zy2REctheLygIv3IYYLnSySr9H+D65
+emC6JzLAuF36PqWVf8W83zmg6Dg6zh+zqQMbJ9k6bIinpgEvlMi8Py9gqelIY2T
JTjoviRwf2aDqXKh9Vka5Kyyk/YKRjqF6E8LZA8G61j7tgVBUcUKoVF0JsibSmOX
/tFHDS2J7mLEzBqacHVE5c892Lg0NVSO27891X+QJRFw/3j/Acg6GMwrwSFRhwQs
pR7rsd7mQSL3JjR8k6XQDlYp2xzFw22zvof1XiqKG+Evsxw4VbLyZWGEiPwY0Si6
GS1TJ0ZCHReyK6dm72ia21/zw/rEJzS3wd9kYL62vDqdl/2hmGzThZt126dVqBrT
TRdW/FKpuxHnKiqgOK8QEezy/kSGZd3PYvo+aF0LtQNf7ER/kwildwv+1TQpBpnA
9oUQqZetg+8Xpcr7HqTeotbWr8AS2keRRkBJQox0t8g9oFqeel9BodYDWW3fHhul
hA+1izMkhj+t6iRjzSgTVHP+3YzavvTgXUcaHQi0zNmyLzF7D03N6gsQY31tvs+r
96JirIQlbVKP81oVAplx8ByP24/KqABtTZ+HPfFnzsqUoCmk0Dz4EgMpMzxGrs4V
64fsCB7yR9svKYWZiiYHjjAqI+alXlLJVBGD8dtRikXxMdBXZ6vL+oT6r92uhbJH
PQqoqEYPxF0pgr0cjqI0fOV1HalcNHMTAcNiEH4tHVfvspYdxFovySZGQVM4mYEk
UX6Z6dbSx1FEX6NyyQbus/CA6ln36nNq0xFTQYknhQhjL32DA0ycgHDZ6FimhUDW
icpaT+YModF9s48G8E324GChNTopUXK0VsHDXkeLtb3dExjq5N5dBkHWHWAHFn6+
p9CKdrGa0UDVbKb01hfkZ8aNFjWXkk5zRg4LczO7pFwPb33o63jqqDAD75MAfkQ1
F8s4S5dG7Fw6UkbABQ+a9ssdk5VuPnD8Whj80KmzomEh5xn4v5AbC3clR8M2neOm
hSCyNMeCB2uWb8yAXg/AONx7cEVl3T1/5LRRIrMuxjw2nfOvnM9UKFDoLQlDTIP/
RyTO50YrUDAzp3g5tltGeI6YDS2Y0Nt8vgN1/9Cn1TnQNQgxit3K9QzGN8FzWdOR
5ibyJ5uF7q7UDZjifSaT913HsiSXSxvoxrWkqZIUkw+2sHa0pmu9SIZxbtSlcwdx
gTFj6XTeWDcMJ1ycg0MIl7fOw+TJCgg0/DbBo6Ml9eOD/ktxvd64wRoLLC2NcKoe
kQzAFZ6xDAkfLMi3t6vgGklz4NZaN85FRpVZOGHIZ0bZ0pZ+I6KDPTLDNPSOcSN3
wjavHNQQa6f9qZ8yMXS+O3M/6c32BgnHfe54tHVMtyfKDVsZclup5Im/gTdILeGL
m93TQ8ZFsoVCfATJda2QpigZln59pd6e9Na6XArwspdhw3mxDuwyT/Y9xcTzOjv8
gIZ9vOmnr3wwr+F73Im7ygVXO5vM02u8RGDvVyk0FTSgLqIqZ37APhZmlsTF2qu8
gV6BwZNyMB6N3ukQpPLAWhH/LwAPeB94B2S0x3TYADmB7xJHuOuHrzhpWsSu1Wx6
B9GCJztGbVKZZXG8iXYIW2R0Y4CqDBbD9pUhKdGtN3SIjv0s8c4e3ZIooisY0SPu
ZeCA99NMI/yAJin1g1pRRg/AqG2q7oATEMaQYM9P286HPpuCwTN/FfinFJWW2OAH
M9MM/ANuz2rUW4fHZJnudWh8ZpMD3ZAS644JMXVUvLh0FnStphzGieSnVra1NWgb
XgxGcWgwFEMfPO8y9xQrpnVGCLl9tgArk4ENh8V8m40Nc5TySDhZyovxz8VnZ8fS
eWH4CBezUbU2NeZ/VHsaRltbN18y1Nbk9HeSvPIq+qIENE5OkogQqEURDzl+EsJv
X+PplbVoPWYBP4ZqeFtUoIPX10qFNM8xQgkl1niDTXWq/OOoLbCbqwQIHfPnL5vV
zJ3FMivVV4vH2+3rLsUDtGEZjIAkWuLouFZYZfoIoErZJOMIDPBHPcRYURDHt6ZF
c3HBx3YJxOvinY6iQTw4yfBByYVSFBpBCChs7egGrtrsD3uXEe4d8KExIQkzHAEA
hxa4M/IlfytzZ6qr+iT3fF9r1bJidQAVqstgGhQa+ouA3dl7gV+R+W682IuTIadY
EREOM/EIOmF6Vq7AmMIQLblAZM0Xd7vVRGo54lYpN6uFXluJz1g91gRKsjtug6w/
p5W3Kt7woVzZBj8Z9lXcvM1QpvWxnxoTYuB5zWE2X4CW6ofGtEZPES9Otin7yRHj
//LPOurTRwyaxkYiPapnOj6piG+d/b3U8Oj8T+dGL9CQp0eRWWCVWP9wcQm6Hgr/
Zvi4EWhJjEeRmswrdsGgVTYfQQfbUYfFE6+Y3ZFJGqtS7YdeArWrSmVdeuWBEljS
LupxEhYoKMB0T3bINeprhUfWzaXERFnZC1YGweDeufkHrxt3PtuvTlNLXawh5OdA
X3IGohQl52hROAzQFGo+2ZAjQfAEPB0fynTCF3BoU4/vgzYCGIuyZo+rzgkm0Z7S
NBlzG19WIZpdFBZup9hGJosxuwRWZIXV4VoFArwVt/pbwk67oMM4c8ar1cFTQM+n
vDnxFZjD/tntQJqcKCnWAvRwfYFugzY7Ta1n2qsT6xV48m1WTIdUkwm8WZGWxtjs
aqhijHSAcLl44nDmTSkwNpjjkaONJTndfXd54D8m5TYmLF1jA5tpwi4VFleOSi9z
FamN0XCYcgob0gGhIxrLzmHb1vj+okWjfYywNhqnXfPvy/h1gYhbPCJVhEYWxMRA
H6GQrwrKhlk8sPyxI1K5DTEpTQFbSN3vJTT+Hv+nJ+2Gk5640HXJcUEnIqv2007z
nyATUjx4cgUuTMrMe1ngKXaMSV+asMsYEUYjaTKNdECEOZOGXp+X86H4dCpGkfq3
DkM+y5hpRoG0HDld47D0AVSiwOtehCN2FCGIl+Bbb9S+oHs1YGqI2cqLyqfTIKgJ
Cqpmol11WNPfFXv4q4bmnbLwWhp+RABb9cRZmB8Sj+vr3r8qTK7Kn5ZB2CsDEZBx
jtuSz/qk06Pdv5YkSJ9InTpC5dxTIcRdxBowrwqfcoQOnV55n6UJnEvKOLQILF1t
jtgisOo5XIZpDpivH8ixn7fX5eySGugrkuUznwnKJ+Z1sYXAbS6YGqwHDr1riZhP
xWfFVFttgkWn7rO3AIXb0/pTYbP4CSjIJzy29GhSrMh2KMhQpWAw6NjcZTtvZb2V
YY2mMyGK+lTKZ8B7erLsFFZBs+MLqgr+q0c33X05MmhdbiG1eMQBjY9u+7PrgNN0
t3Dn7eiXvbqBorqxrI9WrLw4jJ8Vb2bY951lNjwjUSYO9B+GQ0jnGONc9IjT5CkB
TMb/mSEG2yysi5wzhBeZMKrF3ou5eaBQ6Sm1iW0WfZx1uGOBiglX79nedVkJyziZ
l84jXEVgAWhcAEIuAhxvAx2pGaXHUnuonIcN+iwVN+EML4nPqzhFPR9/qZ8Ndw6g
xI4VJgREnU721S28uI3hf7IWQf/r2vrk7Hp9iIV10ZFbpfydRxHAosb381ePN1x9
atDcSmAF8bRO7fmmi21M44vrEL01PXuxcSKwdVQJ1bp8TmhdqZzuQ5250Vvxbfh2
Y2TWie2GNHut9njBFp/DW/qX+S+X9HH16l1Egegy/T1iAzWig47sjMlmrbQFoe7D
BZX+U5SkUcFYdoNGbQccuPawfJiNoVxzb6xXE8nzu3YxKP3V4BcfvNl8RcACVPcH
LY4VYfBgsNajdZVDKMQyPQkkvz41VUU2HIv5adjCKP+uH2afJS6Vbnvpo2CTasqu
GYczJ+Jl4HBVWl6lUSeUlG7iJPObxwiBkj12Bs2b0cg+JG2fJ8iPjGSXxwWD2AS+
hZNZMtbYeKXTYl5XW2tTgjQRE+cKd9Te6cNDOB/mDyZVJtH3oqfhcAWMHP9FKyN0
yA1GrVJvN8HIecf19oYNnCB/KoRfBW56Puzon1e1fBn1p5SBp5WktiL4K2ExCzhX
cUCc1WNHvhnEDB6xGaekzhDBvqqqtyWNuqiQraZ5yFDI5hnFAyZWUiZB54JUqu/n
a6iYugkxHhuFO76DLbREGkYzxWqYK7wP+eIGXaOa2uLpmflGCQ8MbKUIR85WnhXW
60ZOwqSbSOrxQ/pDDeaXElHMX+T4EPJ3JhmAaFbMbc0zJRaCqT2uWwTyFqCrjy8v
/JRErLU4C1cXoXB9h/01tEPhqFMvL+LDbG9qWPtU5nvawQFDR2BD6zqmhL1zuFf3
OkcXwxNTsj4sp397wqJE9JoxzCz2WGOhK8l5dFLsHfUMTykMoLPQRDasyb1YxzI5
wcEcTaHjGwT5+ezm6WV4f5F1VhUlxlBV9wCD++aRIlghkLNqyyC778kiqkwm20UI
uWmyi/9tFtRTrh9cVPVVEkOgNTMYhL6FwERcnb7v+BcPaB7khDdQOiyitbzx0YJY
BkQYDzkGiRU+V6OaKhhltzAF0NTmbbMVHuXvE8mHeFCq1i1K+6HMmdRFBkdA4ENd
vli761w26ApxooytAcQ8Oon5DVgbBiVTnR8G5gDkJitM6JVYMd2c21aARS8ZsvqI
7trQG1LrAn7zsunfypkXgVCMF39wy1mKbRWT7xilOFZfKCK0Af9lqBcJLg3K8q4S
hw+qHxGXSmQukKMkbI2iXQiTNBYiS2ifYz0CsGbvukRM13yO9rfIybJNPJleKdRU
idnvP9gyxgAQC8+JKM+YSn9P9slFA6h5TlFNRbe/zBX7dr1UbMhb4kWSZOSmj6Yg
tzAkc8BlyMLdZn6vaWocm33dhYt4BrLuV2IgyPl+3ZkytJ1TmcVHwCw8TPxPTJwM
OAJX/KxAVApU0KFPWH3R05WJz/Y747V3W8QvpX3emeDEA8EkqS3az+uBL7k91aon
93SiL3BwhofY8KwZetwN6VyEB9PJYHyr3qW5GTFKRXqlapguYrRFbZLe/VRphe1M
eZno1dTHg2bitsGxLPNB9Sn+rtdqiPxoNLdcr4J2HBDMY4611KZU5z+hYJ+soQrb
q9vN9qExcUkk1cfAjYhj8lZuZ3xG4ikjIgbvrUC8a+oXyxIv71BVoCwcFQ7r5ZVr
7czENEb3fcJIFzcljKOZNkWYYzWLoKz7GKMOiPhcAM5+T+ITVTGtS/lg9Dr0IrRc
fy0t4honk7ucYDFTuijcPTfC2V2bs+Ukzq7qGNlF6AdYKXA8barw0Q0+bFukTg9b
Mn/+NzW5oPqrG0Hir1MKCrz0+9qTgiy0X6kjW8/WNwEpn8EeOp9p7cQqdfR9x91k
k0vmP9cR6GJyy+k2sTopo14ra/w1IBK+3OqTFq9eZh+jzCSNxDT8DbpHC92v1E7M
jkIzdCxVpWceSLTUFAEXd4eVeytLuHA3vnnNoItamH9rJxNnJB4wVIwbxaDosH2K
Fjndml9+yPEOjo9H/MCSuz0gSZDVKmFNXkEv8nOWoM64DTvrd4qqX2JuxqBTWCyz
uKXczFsmigcVzd3RjIsUzLxJmIqEVs7ZCNdCva7P/Z9u0sf25VwneQGnGOWGDZn+
tQk3XcWEzx9Lzj46fOvoFVpcOVbgZ65hqLKPpZO6zlbhnHRfkytkv1nPEqF6eu3m
OrUtbN2HrmP2q6oeOhf23zPRyGD2qQK0c+UN6cTQYRqF8SQJ7beDf5AMJqkuTStq
PxP3mGr9VWziF/I7wb1HV8oZ2WzuX7FlWY6mRKSxB28lp2Ky33/cHzjDqbsNHhhd
t/VwlzgmWjf4WB1iTyWzoAe3eC2Rnbp0AIQwLedTsXoNRGmSaPtxH5sML0qJ87UV
NUCubfldv5cDyXLe6zs9iieVwvm8j6HhWSvbsbcomCZ/6lMIjnYuOuMpUV0GzSd0
qlZeCkEG+O35WXH+XJI+B+ciVVXJ759aakHyEqBxTCKX50dki39eZbVoSK9wVs+Q
jArGdLQlLM1oJ9R+KRhmNZZED4BWJAsmqydE8MOeBLOXEcFYbEWmQIawQNeEQyJG
RFzMNTDH5RunEJefK0rdNmCVa/eyhZgd9f0bK8BSDP6L214jMteLRpmpojik0w/r
pD7TkDJfIUwZbcpC+cqNKxNXFJ7hDnhyozcTXFkRXFS7xOuNrXlcfzkru7wEtg0q
z+qtKx0EJp5HF9Tq7ITXLg+N0s9ofopaNmwR73plH6OHCmDWMSowF7Mv0mbfHtTo
OrhjYZD8pV7LrJBsbUa+WDsNUaxNI9mcjezRZmkO6GQTFbbnilOWm47e48gFB/Df
pwd1X9Zas46HG1QpMioQ8fXp9YIEJQaYRtDG114KmswQdOtOjynVR3e9AEZyTcH8
GT/6aBr5ibo7qZDV0oYpy0UMInyHj9LosE+otV70v21VPrWrBnEkLNXA4atzJfIj
D1xQ2pUA+W2ulJyjcsN0bKGzA/vZLXzi0cJNYVIOGAZq7PZei9LXsaj3W0SteRY8
kJYTTfoEpDcEDtJP8YO1iiR+9fOed2xaKbOj2FSncH9HOt7YzZj+bvxPvanZ97IG
ws1YC+zuVIl5zf3ZM+a3si+QRaowNsMzH5uDcGzY3hL8rtUMxbswCwqwJCq1YECm
3papK8LbTecTECZyzvGtXSSCKPXzb5AkJ45mlsNxfK7ijXSWx8cEBqWF0Ox5xKmF
7xgWY5UgPFz3JtHhgD9gdT1PDzH6Z8gILaxzg+fA1mQ1aFDKJM5gwZU/XL+hOdIm
dacuSZn2DMT9RRUxwkYhEiFVSOy3MTuLSgPP2vcfN20gPQdxw/4ZuZSjzpFcLaNI
/wGvqjXleKhYdNx3n5pQfYrKKSVDlM2q4vakdy8PHEEzkS9020l/Ql6f9b9Qk5ot
BUvMlArUj3bpYpcMYZlp4qD8snlfNKZYFc1d8uT1W7R/ynevKlBMyFR50bbSjvQF
i0NsByR1o6p5A95deVinCx73pIkg64xqfuI+9ugxRGaKsx4T+BIyWa1yHQMv1JCG
h3nFT03l7QB7k5kDAOcx8uJxWsQNVJuzFrBbi3A/Ae7tBO5oPE+MPkAj3Xo5EdYc
067dljG92a92/PGABtu5iKlqspqUEU6Nl8Vj1tO04herehZUfnaI+8SJWuQz/LJU
yJVX5gtuhc5iFoY8gmVH3685eFcmgKXQ8zhae+1ei8k1o6U8fsCq7e6bljTVpYA4
Ao6FshRYz2TTZc5m6vWJAlDKKbo0qVBw9BqSD7yWK+Js8kMvThI/bRXG53FMc1oV
uYmtaRDKlXDruCvQrSkyrFFfQ6RPXA6Mr9/0TFYZkmSSFWO1/mLsqZAb1ZQJ+GOq
swT0nepnF/Li0oDLVYs/i84TwYiaI/YDTcfgWAt49CuFLd9FZPZwur1NQTdeuaRu
XOSOgKtSDlD2+D7THZcXsugNSnUxeYy3tTAzrezVLrd+ZeCvSMUvYu7R7NKo/9UQ
D6AjKbVYsBYxEeNMOzaz/fpVISbjjldZ18NXkjSfMyKXrzbMezNmHnBZGXQt26Im
dOSU7u3gj1tLDr5QiNybtG9bF38euZyo17lmv/OvZLvXEC68QmFufk/VTXXJRjIg
bMi9KZrVuFn7ggCsmAwLJ9myulmJ9/pi8+k3QBh5HYEmJsIIh4bOFNE9kYIRKpXR
6tWEJknNOrGqticF4nDjLgEmJQZjdwWqKTOoUzTkQdI+ihkaMxXhoUORctGLjuds
2BqZkBVYAkzz3UnF5/upaxP7jNfBMgJP7FJ8Df3K0YPlGi1XDdPwpJXgSa3zQ0d4
l1jGhIuURRwwSGcKd100gpHJE+7l7S4RkpSZgzxFPNDFnBVfxNgWMTPeNgR4kq1a
bWmagVvYmyDGgR+x49EJglgEJYPfO0arUIKqjVoKiex2EZbNqcYggV3gGn3BQSe+
+Bb8hYTRyYmyutL3KDum39t6T6RRJvJjMUSc+x/oHWKUwjQkzHc/tGIwkNvh5QHQ
aQEzvjAx8JmWmSPNPdnuRip0KZZFCs+RMVLCS/nCudyGKyhiWYb8xoVR92uVj3ji
cC42pCiqV8QzEgqwY6sfVloVAyhKx4AxKy+lCIZ9czNnImT5hrQ9dTM0+fY+J68m
B6oYkx7An8a6Maoea3oLMhUJeepKGs4MJVnPV2c5NIn+LpRzSdU5ndeXakDnXEb2
/bqqoNjb8VumwTIHELlBn5vIVOM7h91epHm/KyJcuqZZt6/U4hTi+allypvs5h7V
rwqhbSO1BJjR8wwwzVqc1Z6jv5o27XMOvs9UYP0krP8FS1JT3OzAcj+Lo+px1W5g
MlBNZEmnA3cbwlWnLDogFr7JWCIvo+76tBcNFAgfr4nLzEqB/L5QKROVO0QjGmYP
kID+fIoY1Z2pyuIcgARXf81XSNXkNIS94ik+Hgeb/Gj+JDSLzSRq9vfR2Ddit08j
5GYkoI27F8xM+hWq1kA+piN+E/JYSkbAJZsPdWBFPKSscxmkN+iSJjtUZKbvH8JU
TvqCzMWr9qSWVNzTz01qeAqWaRoxeftW+z7+KYBhpPmi0Eew6+G3AJBOma3DMc2D
J77jCEWPOIlaAueprtklEMu4prke8G4IMkUKTBh9UUoU616F4rW6J5Ha5AIEMxnZ
4DjyzeoPSFNCGDktSrSMQp1+X3YFe+mBxws9MgxEl2O1Vf2oTl7mCoUzvzRemzGI
z690IwiJPwBpiV32KO7FTPqmQ8rEfTZah56nyJBn1337FNpEXPk6WJkHnTmy2N76
u0OblRqL2DtFEBWTN3NZHKpW1Fn9pWQdoqY7JfnLunafqjnVLexQywEw/roQHeT6
uNwBZ5t8d0zlL+TJ6/pVkUszqesK3DvvV/38MedYDo9CX4S3LYqvz+JJNiefWSfY
hZdhku7zxjVWBSTed4hbG0Llr9LdLPFpi1HR6EbORP6ij8dm4ncuR2hR/gpP1VF8
ARXxYmuf8DprdVqXvtvgWBvUcl2nN+hxfstSv3/Ybl227sZIW5GFBv70PsRTMpYT
fb69foIMUXEB7wAch6mkfz/mLgiTfd3BbLHPdNonJKtmhaPlmpOLMtG8yPhEuLHF
SE1k8NYYlSoNsmgstEruwLsxIepCPgvtrjfSXM/l15n9B8i4Jmf2QPwcddj5mmof
0+fZ6xMmyMnxVvi+T5EsQoSTzU7+e0l2pwYYW4kHcJuuWz7OpcXAwvDiWHJMH75Q
we+rCK/CzDSf+mw55S1SU8VPQQBLA8s0yUE5/v2rZsobGPh860vhlMVq9GQNBo+a
womhXsj9Kfq+YVQD/XyBZDFBczt5rbwhPmBDnFuXwWOHB/ZgvVXyFeuCUUxm/+ov
oVqlYS0VbX7VuAb2jihUGGOvnjpt4SQdUU7lODb8J/SbFUxA2BfWU7vJ2sIrUWMo
pOZEgl1i2/uLI9ZpnrN5dozk4/TaN5QM3bWmRnjaA4UUynrFVmI7Pm/3qh57x8Xx
/NO1rYuW+nl6wppir6JRZ06rSBSkjRqsrwmDy7rooP+OsTMBqtXeU1dcDiX1qlgS
w3tgAhd8ptX6DYZ4J4LnRZKL8kLZCNRe7c28gdBhgOxQFItAX0BhV6C9LR/FcGI3
GTbXbSUIS5tHjEngJm56pYscNFaHV0Q2QqNeqvUkPwZJfCtFu/NEPhNfnLa0qAuK
jeHJ41DNiiizRVw/6IDLR8vM03EGzOmRnu1D/lP7x6O2w16sqTYEfr7BeT95LYh+
U5atYIfCi8SsqA3zSWBDz69arAGrh0Ktx4PxLAjzGt2Rmkn2b/iOTFSm4oXIIYN3
+avxHe9IqJoyYfUExtabb/nbF51SJVCOmSrqqaI5VHOYl3HPxptodoVtKmyyaIY1
oMPqiBgqlmCmSKFUn9M6CQm21IxHiM0ur/vBXI/v978yifSzFKEHI4XeHvKhw9Uv
TQj67VrON+IXih/3KjU+V5gkHqTmMmrgEVWnyZDNfkVf9VMNBbUCHpFZsdCuMh7T
8GoJiAteWjwWjea73F5rte9gU6HBUkunuSrsLJhOKe5ucrc6iu+3wLsTqPdWlBVm
PtgEHcQmxonGLrwcjsIdyVxT/uOIWzocQ1qUtWoLe1KTNECKTcobk7q49zruw36j
76Tuf/zrwZXr8ZhwJJlZLSrgFt9UOvm/qxENK8K8uUhotykc+MqV+UVIHn+DCs3U
9uuwMU7liKvbaD3BLjXfbr4sX5pugpFiv/YSbtG8QL8L0BkmRF2U2J2ouCXNa2YZ
5solPmP8rDwGYqyvN4+oNaFqxefOo6ivf1QeSd87AQtqxGqCL5RgOlQjLyt68o2C
x2FLFZcnVzw04dE+Wl+0ltirQrk7MsJZVpgelpWc7T5Z93bIXtSmVJAjSax2nQQW
ueKjfh2njnhk6520l3lq5QSnJK8Bao1v1otgAwlwypsLfx1uXD8jjJniNtTrNrT9
FAZrcXDEhQXP5OLBkY9dk0+oARhsK77Y8MBnmVmt0MwX6Sz6mc24TSj/7ru0TYSf
d3JX+tVN7rx2plmwODvqSbUEQ+cR1NpNVCQ7eCmaN4x8Qj1Q8ILcuB+lqhMkf9EA
Z1U8etSs9kSK6xMSnyFxWin7k8csJQC0bKBRySgqZJLeqaGtueJHM/yhsiBpDvrR
TaHHqI9K6TqwNRzeXtwp3eYfDZMpaSTWpniRWZ7pE4s8H9jWSzI9CYBzpGdV0O3m
x9/KHJ583PrwXqWsgDIFkMiYtLog2wZXsCcjuMDNmTrxsifJYGIXCi1tBIHPCgiR
hBo/fIdxSGqcxFU+GQl7QHr1h6/E1CUF2hBiV97uwzI340oE4Y9Pf6V32wUUoLfN
YcEi378202OT7e+bjcCNTk+cOvg2M2yoNmpYHhtmsJBLNYSA85KEkQbWOCGy3MCv
q3fHlbYgMz2z7Ic4VShaxFDeTG3b3Db6NbLfQrfnijjXjUTYIYpbmEjj+PwXYahp
vrcQBeHXWj7H/YbsA6mWB1jyCR9qOgfhGmr8Pex1KlFWmeEO/opBrcwa7if97vRP
5Y/e9eGPCkHu0COYtXSLNvUszr/iUe5VUJlITgU/6ddvD+X/m7ppFIpZn7H3Rx0X
DEnzmyR0f+cphbhYmWJjoeE8FyLlQCmwcHKxGXFmvVG5y+mImzi9/A0Pz/CGbifC
wjX2cA6RErJD0Pr9BlZ1vwTDCL0kmQqSW8JhxccGkSf3PjiUx5dx1jjXDBi+VBX4
b55+NzhjCSEkB/vrPJuOglg1uTGfTBaktLseEVRU/6hGMW02dccCSXQ5DrATGC0N
SJiSIDnvmTPvzska7Rorwi8Z0anngOVepRxR3ZRT9Nia+7eYqRgGlvrbdVu/gHiA
Ofe3ZF77JuGSD+ICa/FaIi8SYKWUXo3OzMt7yXv1EjJa0XdE8bbLv2u98sIHR0rC
w1W0eVV33dzKZW0z0fT39/I1PdivqyDzxBnEN+SPdFLX7kgdGBWHJ1BIqKYi2Bwy
nX6FbuTdNJUCgTNEMbeu+41j50dZgTtIWdtHvczqT12uMT/VzybbNF0uP7JEYG84
IJYVKs7cWF+5sLQDwC75YRnpmWaBvoDbyjLRTNi2s0GxlmL7M2VbCkEM4FDfm/me
WooubNlJ8V+C1VH/gEklUZlklT3nwgJf9YuKABiSzcd1HbIOEapc8nihNaMvvf98
qrCuXvqjtdY8Z6/qSW4HAMDHPcWOJOp/3GMgJf5R3WcNu7t7dMBsDYYu2eKQbkUM
l2yGVL/P7DwaH+znW25vuMklKHY+R4A3JHUU8cOM98THedIXgJmKW5ThWzxxXRHW
C4C/rIAetS/1aEvz6fldtHINf4Xe8Xs/fsu7HyTaSTmxPcIbSxjwUPOk3ijFI4dS
f15iNuy30b0Ust4IiVwKSmQqkvLU4uA33Yd+daV7fFUfxsbi3IyzAE4BzJ+fVLek
R5NvNgTeDmHqDjA46l+7qXbj8ICSL6uDrUsWWuzLxnC6PUVEP4OD0HmWXhhpUZCU
VOURgeOxqv+z9PF0S4M3FRohoiZcjFC80Lv7wVyEYYYGB91AHNp9AMqwYThA4GOn
IFPWrDKGvl2UrdwfpVVa09Oo62fedeOPeMFREHAX5Lco1zXvlEp8NIjQtTGNs2RN
N9QFniUEnbre+T1ZAq7ZQ/pSDSpZZoaQJ/CPjT5SiW5DUEfBjSg/y/V/ETCirWGm
9piMQvlgXqstFVXaf6JwZytssY3XREY8D4AraeRPtFI4gF6VHXJ3YxzR7s8LZDzj
rtq0Dwe2EQ4JBOarcvAWMz01CrRvKzsmtvE4h00vROP2OY4+ZCSFvua5eAnXOse3
Lp7W13ePIRx2/dFgQ/3vr5WlzmYTyPA1tQPZiHdo41I=
`protect END_PROTECTED
