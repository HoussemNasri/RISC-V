`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dDWp8j382yJSTO0Dv/2FipUsb9+yCVnL2Cvh/FZ4hT0FDEFma8tu8K9eN1LXRJpU
kMF8QJYwJZzP+9rGAUsi9yFv8rhJ5ngvml+2JgpNGUgjoVAxUhDVNMj0A+Sj0NdW
+cTvCpq+5rFApq7XK5TSjljwTaWCwg245lEs0VG3xgLLa/l20DsX2R//KL+W7YGq
jzH1UobvGQmTaiZuW3njRHFd5AXV4ezVpdWnKeEeTEfVZiXIGO7074fMIW4LnAmG
OFf39Z7hHtiWju10j33Gc8OZj+zbB/Kpzk8RFQyV+mtXTlFvJxYEMcRIgkm3PDA8
0B88Q+gk/yj5v2G3NPfoD9vVcC3dM5XkytcyY/O9NfvB9b5975mzeuUryMpWdT/h
3DK4NSTiPiubSoBhdWl9xaFU1Jo/jc2yQMexehDsVU/PmErSz4Ng1OWIzqDgXbpu
aj9nai4XnvNJOXLddQW6bwok8dZPBsKQNDIOaXyc7x6R5sMKiZ87GzDxQ0fvg8MN
brUNRhftdomhCzP0YJbqrM+0zIwh00lpgpVgN0lDxA/3hymt3gl6IXgaO9WNvdc/
BjYAkBbAoZh4cgcspGXR41Du/zMA8tNmVDT0qP1O/rAu0hG0YwSFZZOWXz977/dr
XHCfELJGTESsgpYiAxpTFSlg/NuLEid3wvrXHpABH+mih7rmtK90SDRcUSaKEMUS
ManPt1OSIoIg0+DHfHfnxUACqZrFZreSgZA8VyTYuOjAEJr8MCVjJ9B+scvYowv0
7CrgyyGs6KPslIWtbA3Ta6SR15ZfmlcN5/QE+wfURqZcm7niAtXMgFr4KvXY9/cE
DcBzPFLHZcoIzZIMy/q2CMUuge2ygl0rMn6luT1YgEGZVS+7V7tO4BO2qNDM4iX9
RA7G55SLvkmsvPcVCQdCDfgBZX5kb6rkb0VbLtzijsfAuCdYDjnbpeVkMM3Gf7qy
5K34ArRSjmm7FdeRooK6zPvxaWtCiZN1YI233+zddhyfe7yndnIwp3uoZGcBcgwS
kRmMEVr5htidr1plvlPI6mbx2Maw+MJ4JE9nq+uJy5wPFgX0zObL4hLSuCCYg4jI
`protect END_PROTECTED
