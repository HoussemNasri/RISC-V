`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sgld31P7JA1tJ4pJar97/X/n6hpqhTkGGyQ53fQa3Dj5/E2XHmY2qwjdbpgvzRnQ
dpQ7gAcaeaF1V9WNh2XX3xEYtPSdm006HznbvU7Z1zNcfF20ugTsUqL+LfqvW1QO
/sVB7L/UYPyqPTSig6I7tf0PkD0utnKY9H9edyYoDCu5/w/MAxlrgqKSbxf2pHgx
AwDSjBqK1nSajoRpcWCkqMtA1aWYO2J6WEwHP/piDxGTxObHRwwJzTnUdXkeL+TE
RSaHeNhIq66Qp1Lpmmo9Hg5SxSZwwQwgslgtF05QGXM5QsOhQg24qhb3kEBzJdNH
OEtrCfuDhCZW8TNxAUxCNud0rGaEplbCjj8XxRhbWr2YLqe0ssmOSRk/Cz/VgkJp
713nS6MH3CHz/nt5pVCjDg==
`protect END_PROTECTED
