`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVyf/Zn4FGoHCPHyNZ0jqDFe8bLVTlNnBg8x0evcgu3XBz1xrO82D9GomX5q4WPv
HoI2SKN6cG0VZB3L0yAKgPNNvzXXFXT3y2gslm/MIlmaJotd5nLWZGq8Z1GtUwTj
2CtfTIfIsgrbp97MQnlxo0MnMGJI2OAyXtIRf341vZU2URmAt2Hw+CL61xdWPUhB
9iOYP5TXgImm0IiWGssaGVYmvLPYURto3et83kJf4w1LRNZEueH8ElxwhX/cjm3U
rnS9snObaqzwoKHJDLvv8JPW5eCI76aPFaF1dYuPM2VQOSPoGM6FfaP2gFSLR6ZD
/YPdw1+9n8YVR1faZA8xnLBYq2qZzvxEC1zChpY+H/YTqE79rUIR0h/WXaPaYfYk
Wpnfn2KNBdl9g0uObBsox2kJISMI3acqpxvKd8z6Q4KK7achE6WiIjIUnMr2vpc0
v9NP9pu6cB+ZEMHP+V7ZnjQafwi6eKcWMrrMbijt3p4H8YqNxKDrCYEPQZO88kZy
nVNPRH0bbDcPxNafafu33pTqaiw84MsGnLB8c47Tn8D3a5JMXQDGMmJ9unjfCNmc
730tgvNvtiwEWEMAGzf5ValQ4tu73psj+VY5MSiE4osXtqbJ3kAQy1Z5bqiGrVF2
vu/X9mvGsOEKXun8TOzZIeitOBOIlfOPduglnOKfXIvjHi7AU6MdT4+O7jijdMD8
U+XBb0HSo7sIo/ZGZLqYz40mv8jK8OrjZ+LDOrJstcTWFDmFy5irsotn26kMl4NQ
FlkTbWFbbJNEXRRlfzE9l7iAVytpideJWPdpRcqFw4OPvhOR6hB8XRdtvhle3qxW
a2IqPCwqNS0fOTFF6euRgYPpzUSQjKDW6qtid+517lgkTpdnHm6cGaeeh7ZwKKud
bhszJUzmk72UANn7BOzk+q8AkkIyDWdxLqjyY1ppA9Z5nhcXD+PrcQyKZfV2omfN
BdztlO2PjdtdQz1i5LcOzrCSp8rTSvHSUISzFMAhQgPk2K1FnJ8gNZkcp3vJmW2Q
X2KwtpV4YD52hAUT7MGxF95NaeDsKhKYGNmNw7b7VJhHF7wfsJSip4qReg+bGJgm
p0V6mX0d7BCCE5rbpttjqDxFZeD1RX0d8eY/+7uedsHtZXAnRvXi7HJBY6E3aXuC
9ZmILCSFWkO8lRGUeo2cKy9PTbofnRVuMMnUun2/G/xJrAmiHVfXYX3usZF7sKzK
bvGur3qswEQwl3geqM5JLUwNZP9zDIOXy2NXH51u9vfEhPfr6BbyYr42qy7TCTGd
3LpLxeO/1k790wYD2TTCFqJMKZ8q8q3bo9COc1+x6+lVZC4YLTeY2Gj+wlVPgGaP
HD/L6Ge942ID0wGUuK9fKLK58GZsu3zLeSD1IB753vLvRI45YVvjreOltpsRCCNJ
YKApXUp/a2O+A7Keg0NU2w3sAHAJYhPO0MjVYW7UOJmvPpt6vTQxmkOoMIgOkKeU
/jMxZDZX3ikV5c9XXHcUYQzY1q+eCiG8dBJt3TjuJRMckyRFgPCDGOGSqGHgfWqv
NisA3q016cocoKLpV1ERaOGiH70BsMNE9O8D146oyxITUiWC7ta5UCRKDptVFfeO
Tgq0lPOOOm6I4ol35/LSVtc+2Yx+ddAWZ8ztteWm2TaMZO/UKZVbLLY1GIR+qL8L
RKsmMiwReRdBRrlOog1iwbu/BPTOXbXktbkTXDPouBOSz2O5LNBKTQWmjQHjmq4g
fdg+381S01C6rytHTDur//Wxs//1I8n16L96PerxDS/fLtX5aLXtw9H5sD4yT+lQ
zaNrG06y3Xcgh+d6F0MAvbZIKFYurD7Rdge3LjurNp7wvkUe1EPLVvJPWOtgNF95
s6NOlgbI1h1OuwjiRGemB4NgnTVjYup6arOyhjicRb8FQ948IOWOoF02kMQ//HHH
RXC9CPJ3BsfuPzc/rXy9awLndjVQvTAqk2kUTJ3Tc2m9MmkVBVbzGdke2jPp1cmC
f+1v9oU2TyznOoMjQfYByz3I++GzGcdKjn6+is5ob00iKETfgaUpus+VaiUgFB22
n7gFz44mlHcvsm6OaGPz9Aek+AfhIxV8Ur7RFRe+/yYhaWSDzB8Ipr8cEvEX0sFE
NmHY+LTWk7aix1ZEPjhjX0vaC3gi2y5RDSD/v9CjaoTBo12QzK4Ti84DvgUziytW
BkTpQEh9jytcSZD89CqPHUl0IpKFta9IN64799pdo2v8E1jEoo2nTHqBX+dcVzC0
xV4hFr1MJ9bhnfbXB57noKW5yt/o51SW7M5GEssJNYFU5YVsyOy1pxkW3AcKcH6x
hXE3hbSOy2z7g3fxQUjkSiVrn4QmpKvWNj549NQBoW5qDdl5SuTj7lPDeasFaeEq
IbIl7L8BpHjiyQqX+WtY7U48iEP/rau8WxK3o/2PYmEJb5EAEPkYAAN22iGy5QyI
p6WuIAhrOQgIEGh5LOgV6HB05pWTzYQhdETR/gvlAv7dTQ//TBDtRQ6v8lD9pjcO
gtrY4FepGcdLbwHJ+5qgGPKdw/LpiLVoUtubUOk64F8W26c/babN7dMfeX9FSxmx
mZ5fGKHRoCqc3+qnCXTBWYJH98Tqk5Nug8vOq1KJbMJX2uKuJNN7xFLN+0DjZ4fg
y3Ai0OlQHALoOQMzghokXWjGxiOtkKKqqoLll9lG9DUj74LxOwrRu7Gs/G03fazv
slUKmS1VxEewoOQvYJ9o9L0lpnkvpPE0e7gEwq6Xe63gW9mh6rLlKTEAIgB6m3gq
ZVXX5C5jPVqWyTIJcMzGGxIAqDOqXC43VZ3p4tnOzjkELz4/ih4pT3taiN9DF7LE
GX6I6HmrT5nhj/k/DxVTkP1Pt/eIR8kJX0bQH52EqfF+2+41MNqLz6aUMC9yNfFV
TYLLxnOrbxYMXe3IdH7949sbs2hBXbdidpgc0Vq5nvzlikVBapppN3eiITGbrgSj
eG5//8pSesI0DqQ5BabvbfvqOmhIVgPCFeN9BHDhV/4zbHeVX7Ycfok07m7i/o2Z
k+5gPs3ShMrB0N3JSKdiBnHrt5o0tTh78CvysyXZSS+s13OKDD0jVsHGU32mf6lO
aEs4lX9qw0GI76kJcJAoqJ/v60F4fRx1s8bsiyBzrmYbzHph/iI+jDvOw7yNoTIY
0KN57j9V4E7rTYLODmKZQ9u39A9TKOznPbTRlcv8EV6q350kZHKvQZbZHX55/pQn
5+v363BgbtYS/xOOqPEtdCcy/h2B0KUsolDo+7olIDboOAHhbWg6CkaD8GXelFLh
SzM6pVgDDGye9SlYlOrEMXK1oPuq1drkFlkLRsHultLn0IZjEpgyzFIdUZaIFYP/
IxDB/r+G8m5NvYreBgupJRXWSllrlwCyhNG8BxAMhUbu7CBFvXdoxHqaJMEoWclI
VPoQqohp8bLkwB5kQzlsWExz3k5KSKAAGTKqtwdpx/pnBbgb239DaLCpbToQaojh
vyETYaPsitM+AYg+EJD+KdTif48T+LqYfl8DdXR/RsKLowQDb2suOcPXuShP/H8k
bOi63tQOZQjKrCLSib3a5jSLIG7NVsq2t8ik0S9gvqtNm9Snrehy8ECve81XzNA8
crI0IGTK4vqF6rrg/gJvyj+H3RdSQicpd+CxmTm/A/JnzllhK7del+pSLE1XxQaA
j5DLx7DMWOQBkb9HaU9CTcgLkbN3JPDWGWA+tWPDnlr/CK25FRflLvFtVfS0Siti
M0sLMzSlyp0X4d+Xt8vfVBEd59AdLf8eVQxWWQBk938TaNrGCJhtE8NUfuLcgSsh
0mOkyN76KwkJ19/wk4DxpodrmGDlefA6+SyNAyk1wFAw19KSiOVmFnZJdumxeFVg
UuaWdo+B/wLugeDBNqf3L52nGQDogydr43iCV62VdIaMVIuiWLmNzVVaE/xRSQ3x
+ivD6EscglHUVMPLywF7azF0pXjO6zK/WbUrz0TGGDbELn5hc8JyKCmdU8X4pMiF
OKVnMV6UfKU3vH46/We8USxbl62ygLWoKwScRGTogJTHGODwFTx0kvgV+/lwTgpS
qH2qZ/W1FFmy2JoJE45+BJ8+gCOJKKZCEqfkc/7pq55stoJIMEA5/o9malnKs0ih
AyxKKldFXiea2bZZQCAmyVJXrx9wyJFZLsDiBTdtEh+2/YLMjI9HhxPCFRJf+wqz
yw23sqe4gpo9wRfaaknQS12va/UZSBKtalPzFqxpDUzHgf1ZRqwsZEoGYVNLxbvY
hhIYnHvAKOfIdxlHkr2HrIvoCBymMXX96ECfAKuWOO9Er7KNAk8k7h9a65wldZEC
WZXbANtdPzvFvpovb2H0T3zvKw7KTruIym6pZPNzAS5sGI2Z7cD2zsJVcR9d6iy8
w7Ija7MnUAUJniox3gumpKHqisPcAJWbfnm6S0zUuEqeJ3jO07ZLG7NoQT8y6mog
w+Px/r7vqVkk2jGf8JsWqC3TumaIYFuluVfp6AbXVxps0SvdMCpJZfHEou87T15x
biuuUcOI2Br5sdolkIvTu8QpSdnFcWmPFTMS7KzaYOYf8ulvT170MrhYX1mxS6gT
P8g0uRm3ZtRHru0ZbUAI2UxZJpSvAy0KkY0bP9hDgxlFmXnP6JtmV4j/zyZnSBXX
ioSdvmWa+fdZkY/FKTey+8YS4d/S+y9nuK0ox9C+Ee7o9NfMitJI+kkeV1AA8ym+
cUbuuo9RUqWiDFRIstTMWdVYAK847aZCKfqcZikA6V0+mPQ129i3Ewub/dP6rC5B
L2aTLrqPOxHWAHxA/XwddBa4ib4idkhrSfYlNQ96xLdjD7UdOIRTeSabuemyYaxw
KnehDqXqE87rDCC4wpyZCfeVJZ+WQRfLkOi23zv4WDgjtOCJZaPu2hMpAzLvPNEv
8aVnom5OeNAwQa04p/lTmvWVkaXAeFkyLoY3Vkf2HhO7NuHOqGsx768DD0H78UnF
UvLDrrMA/xGZMrxMifc6C8pB7LcbXSDkvKW1avDIUHyoj1ggcityBY+GYSos3ULm
YsveqdkBGXhRZM1TyobD2107H24HxDifos++CPZYWCaeFSXGKv5lWNllMWYiORgk
XvtEtwkI41RhfM3rrTclQzmnOeab3mevr3/Ic9dn3hjfHsvESjEXSfPTV7G5XQdH
bIaXzwMgK5hT8LF92JA23ID6NGoWG2iSN61y16eswhh59uXuUWgb6Bs4ghZSmAeh
mr0v/cjL5t9/AGCfTBEHc4hyFZSRPYIbtePjlymtMcQ3NcaV69e9C+iYgYYlSeoD
wgvrx4ry/DRHQRczqr6u/GuOjNBIEDxRNF6Yc+5yoXBUrkOmVSnGurrh0cv3xNPG
fKuQGuDBcI86y4IybxvnktR5cnkzwhjtwMKSA+pIo/nIElAr1NDewkaAij5YkIe0
TX2D28lPWZWHsyHP/1N3stLmt/8Wu3ZdfXWh4noE3VhuiQ43QRuCQnjVM/maS+uc
/l0o7hdkM5KCbQk8aWWZPo/kKcOFgDezz/Lp9g+71EH6oev0/7rTlTf2pqzs1HFa
UVO/dVjxH07HP+WFV1mVpbrpFdtXQ6yoUK1K9+0EsXJUPwIaShQpnt7ryh99w+OK
QrcOaHaZiO2gq1Xd7S4y8Tky19uRExD+kpla0skwQiNXZxiYwXjozL7baNMvlUCA
pNbHACgZ2/Dvfu+xJ7wHcxN+0V7wmlo8rB18EDnJvc7TWpkH1uIz/Q8Nob8XUP2n
lfDkDZREvomB4naR1ZLygErEbWeuyz/bzLpfVrHk6zrtfIr0f4EeQUiKsY69OjLe
eEQLvoWT3uRQe/rZjtyhjregl5dvAQuaKELIoUuvSrZ6ahZC+pDsAOP6vhgW2fMK
Ui2mnULGUyN0givIapseMU9UbVz9UFHfrzW5IUggpSWAU8QqQ8JOPERmnBaNDdGC
ghBmYzew0u39Myb3L9AgK999NBCm5VIc/ATmhH8dDga9abCbUIkAkSQ+RdWfXyLf
mBNTh8sSKXTo2gs0wVxeKK9YdJ5W9eKlcqgvgZDBUnkr9UiY2oQ6daJrlVALLw6p
bd8WT6xbsEROBv/+RkCZXNDd/mtIKlzaO4u4mz9a4EP57/bAeUxmsDZSmGs7Wpz4
s52aCxG7yTLjRcsyk3xfoB3hZdL/7/o3zciZ66yqVvl1bfZ+pW47gUv7S88jRbFp
CBOVc/vKTU3O7XwPBu1TUPKQ/2lLnXTeCZ0Qp/RpgR5RV6yapbReJBHyhyO0n6vS
uZ7C7isrT+0yMMmv4JOCiGS3KBRhv696esAZ8yRA6HWWH+V+76l/JVZCqv9qZXOP
cpqJIxHLVYwHp9BrGGQBNvOEKYBeBlXIuzLnhwdGXXVH96RXVmZ+NSL8/qOjli11
RRK0zROyyrkBeAJA0/+tYQXx3oEcfeNur/3NbiDs8fa0bl6BbmEUPzZgPBJzQu+B
AHNnyfRDrkU2c0LNKjSMrrtFrFsVnRuNlZDAjh8GTDeaOIZSOO/KEKq0vpo6Ggjp
EO4z5wsKKfytlxKzLcmP93xs+ec5hrwc1lKCmsFiNXTf/3IYW0IbJoz//e5gxrCb
gfQpEwtZK8X/qe+00s+YdHRx3Aa6yHsYlWhb5FR49jSo9OXVKMdIQEy7MPxVmAyu
PBvRMIvgiCC4vJnWxFef90g2keUOEm5Z94o6HA2055gnDxGxZOry7aXvf7rTKKSb
1rfWvapn8b48OA+TT3/aoN27vtedg3hb7TogD2YTcq9+jYYwyGXhh9cYA+0bLplu
l7lI6d1lCt/Bb0eGmfCEk9IY36vyrpGHLNfV8WMwmP2B1eqfpQ1oH420gtfrpiOO
84IZziIH1ZTXVf5utQwJGkhAVt1RXEnfWKOELyrN8cCGvE6buc+9BFSshl62u11v
Jgq1+sW7neoR1OV9sDhqZHXY/C3+4MNPrc4w3Qlsgiljrw9HRFdfFekp3zwOowd6
0fvQLS4blIBp365x1oj7yOs01j07s8DyRrMJurl4r/RcOLZ+dLZMDFT6SgZrJ8sg
ZrzYOaF98rCFEE35KpWJzLPy8WsGjokNLYZRq1987PmIb0iVmjNvhUGNvSaRkX5h
EHwMevF9qLDOflCo7X2WyoGFAADyn9D26YTU8y7VHkqNyBnah3lN+XhegWs+2+0l
tX28ufTXA7RdLeM3YhGCDk3rnYe6GBH48s8AIm+/y3Zvpde1Pvy6bOl0wrjATSNt
fjW3YjIK5qp/pNfCqEyZSp9r2IoKhq27Y95X1ykBNOt37PCDUaRVFfCPewlobz3V
ADucG4jRFwdv6YENRsf+x7p5oVfP/IQjCqEkmqoEl0Wnps/8wJivLVXvpr6pwzqw
ng9Rd31j/vMsDEMRUS28nf0zbn/HJD5BJEuV9gPPalVewc5Mr0aDPoocH0/HjBdO
doZeBemkwWJS+1+c1RbZrp7Urx7iAwxm2FEZqKyIIVX2s8Xjy+tTGGZ8yGRk9lj2
VXt2k+oOVW/m9MSKqeKULi5kJhq6KFeNHCd387llBxsrOdR2IPpV9y85DfzlLS82
7T6b3AZkMbTAFJUryRck/u/HiFT10zT3oZtZz/yqAIZ8CJoALrekD22x2FTCudh6
jDZcyvSUM8PXMe2aKVrOVQt0IrW6eVHnIzygfRH7xGAWALV1oMxHXgw8gjaOeMMC
9VYMqV9s9N9+gjEYJOG3hntCfF6e+507R8P9WaUns9BErA/MTOVseQM7vy/5sMHi
EUAHZNMGsxrmzOoFeDgMKiyuls0RcCKiNjzYQY3w8hEtneM7Pq3+LoJ0d6fIgb+c
XXgyZOeqOPi6DA/0qfs2Z53f8eqE1DY0UHd2/nZjpM20wTYWnxQ6jqkM3pVCltXx
KEIgNjVHT7f3EDIw9j6e5cTgPjVPIyY45VY6UTJSQBxTxsfK1Y31eYXqxLoWdBiR
wBGrxt7+/1VcF5bY52mJ8LOo9PTBMVIzF54Ry5XUtEXAvV4ELdtaEEZkj9WMs211
Dz5l466fiCq7qf6PkQmk/TYdf673shGfac4CABaKOn/86/S7pA+lh40jXqPrTdFD
LE4sqTJ+H2+rE+VDt1lcF1880TMwsebuvWXF/c78mR9Agaqymo5nWL5o+fZDs8V9
LHujJdEyN9Yqz/S8dbdPczYUqNHaf6koBiN7D6dE5p+wU6IDYUxtqiYgcYgOJ315
iZwRTdEemhkTQDBm/8EY9LlRLX0udvg+Zp9kpeGCkAThg1K2YnESvM07soT8MBab
+/RoDMdI7Dc9OE2eFjm/+01YNgartccxdc0npFQq3Ncfph/B17xEnt7A0/YBXnNq
hhawh2sb5Qw9pbfIsSU8GKYgMMhvUGWWBGXRJm4kKKv4ruGhttF8erVe/bRJNcDs
qqLKm+vXSXiZfIOX+89W6F+2yFsnzHe4gkEcxhbQnqusaXdkDmItjBpVJjXzHSPF
FQSM3ydwLF/Fk37LaOkZy73ZW2divfkiluAUg6sLulaUFUL/GpTiHNy6g3yLdddO
C4ipVeJyisEULLa7LCOfuqdku6djvXJA75SlFSVsdBfieVW80p+wdLb5diPc2iCE
XdTgE0LIChTRvbs1WchFh4vB8olF2oS1t9Vxfdd5VQPbPzD8I89rkZ2I4nRcsy4q
wm2ZshLN7I2V7j6zLAljyTl5AyhGvGmqcuKKx5nm0TvGDNPbUb0iuqnsv6RV3yVG
91gs2ab/yj+tqxPnYvM1Z93+vKJ+GQ2+qnSQEXXxo0yySenHvaU+BymdayLKx2NN
FW+hcHJ92yHUWV+6uKgNlY0ZRq30RGoQTu8CKfHoPoZuI6/OQWbgowcoqEIIKvH1
r/Dex9zg549y/kRhXKIsH3C3h7Kz87HmctsnsiPqyNRP4mskpFn3Rt+sU3lqRgVb
bacn7Ro/gkrGXzg2bfBGRKDM+QyApKmmpqoI9FbDjaIk3Z4ek6e3bgxsPvE7PANO
AI4y5+uheDw/WNzz+OD/J0oZQvednc8U4beLrkoMjpl0GxSvPtrB1+noFCQ5lzQ4
eXUkAXI9eOcZzcXQ7Nn38um3VA1VA6UG4hA6V925pitkEcqx5AIuGINH8kxKs9my
jlRQS0MUOjgFD5saql3ZAhxrgk3+403IHcfkcygbMB65h3+KA9svj3jaCjXyRxsw
dadOn1Uf0bs0sG89r3yWeqwVSlXMJB9U/3iDGQxTeJmWu4CfLE82BRBOdr3pJyXJ
6JJDItBMQ2Apdw46iFK2pKqWJo26bDzRamQrBJ62xjLDbBRcFD7M4GH0xuU596D0
4GUcjV7uhL3au40srbr8f2ZkUvvRSh16MbOl1y74+ihnfZeo7+4htZMtl/rt61aa
JhBXG1Mqpjx/6joPNZD5fctk2p3ygTYxQ/wLX0+vojA+04so65/VTcM2lIFu+y3R
ugvR4EApshU8jYyYrKGYOIB/gXwc7MZ7VsY7xrRYyu0V2/LdOjlMuYQ2xCJobz4/
W/CoLysW6PFwYl0rkXrvx6McpIyXroy+n2jqgIhYA8RJo13S/oFiONReQDIz4Qu0
BoJphHov0eaLhwPnBMlz3maoruwW3MSJCkCQ13c5FLXKpg2NUsKecJC8DObuxk1+
s6eYkpqzuY19LPz5/PUO+8e3Z3HJpx0bif+aMt4h/+EooETbNPYoj38n6h7EwLtQ
shMNXsGhsG4vvW6+m31DF7N/0QaKkVFatw/4DZJ9Ztw1ipYOF7ZdnfqUp9LLwp5v
VbdwezN//7OG4Y6mcTs9fOs/XjRaX06qoQhElyKJNwIBzzQuj7ehxinUSaXXseak
mHeDLkfnvaCnUTdPDJFYPmhNlp6wfFg1DZx+Vs0TyV9jTqh5qML2d2d6fJ8Dq32i
6EWnwsczdcIpbA6twfyVYgfWXmqeto4luX72OYVyYwZjcyrRLPR7pZCg9EIBw7pf
QZS0MZOdE9wkg1RaUR1T1rcg9DN4hY5Wt5kPTlTOYK9RhC4xk5kJPXnDubs+8qhC
PjsBx4NNne7Al189zJk7ksYX89nRo1k7lhz2iZ4wQT2GdR7HdjxnsH4vLxm+lHn5
YaeTSbCUc2PMXpSEJhb9CkVTUXR0iXcXKmi5rl9lRUw6ldu/gFXiO5YxyHb2A57/
HsI8Ncf3iSk6XGjcDv6BFszfW1txJzopTWhjQwiry6YbkEMQgCzdG32l/FaA32UY
HKb23pZv99MEuFTJh27D75FFXZN9HfBNQDc0gpYKcmSamoDVzAjiftpB0aY84uO3
55+b6s2rOu5Zc5fkJuqbKNDJO0J/AftcLbfCct0qWOtVlCL7PF19b/8CCqjOZl5r
cKfKEmbwbVP2lgI/DH88LY2PMO/bItfoVSTbRsIfm5WqWUKrRj+4mOr12wb9nyyY
hB9ZZFEgxaPKqCJdVOwOb8kH7nvtEDL9DIFbtd88f0ysAWiFxu7NbOXD6ljon1lt
FHrV9DAfgLi74y4xrac+b9eZcdNYlRlIozYVUODlaK1mTHp54KDLCvaXBDDYKL0V
V2Yir7RBORAn4OL76/nvbZxM267qkmK3si+3rFXvla5Aqk57ZwhjeXQTASBfV7LA
BrdnMUdxeqQjr78uioXoYOxfchLSsP36jI/LmBjCa/7hmgDXSaPmUyWVUxH5tPwv
odOZtJvJ+Yfm8CLePLkiMUhLATBlytjKQJ9CBzdzY8mk7pkg5NbGmRKonZEAvJlZ
m3EuWeX3xZLCIpemyHEZq7iEpxPZJvzJPrd89lbiyyDZ6V9I2Q+bsCrTI7Q+4jIa
/f3h9h9+Nuw5XnF1fXLSKJA/fa5qQJIBiuJV1Hl04V/Jes9SeIcH/0Ij78p0Mqmo
ei72NedOit7ZzuWAvgghyFmp7cEDVZjKoBXuGC/CzptvXuwPwSg4Ula9EULS2LZk
F87ubCLlozukddMgjmyw34i3RVS8JeuoLwrujjpI/9wv+m3ijx8KDVMX/cgv+AXj
gFhQrSwcYIK3vxxWUa/kLRnQcZRphRPcvOQM8bmoEYSZu0BjEG5kmMdNPSjNcZYG
2wztlCkefnHNFOIZSnfCkY8vVvi1LHLux1765nVkIZFMFDNMVNuURRgRnpO527Ry
HtnA7mZmoGhmmTktjah6pL83a29FNsUfBfZlLBo7E4N8dCJTQM1hgQIxnRX7wJ7n
pReXNflhd0XptH63Rxk8+X0uVSW1NklFVxESOjclqm82+a/200fB8snUxfgnmpVm
JBN4lgpXgyA3UPRpZjATqfA0DIP/NzXE9s0Y2ZaFpsQaYVMjg4+j8yZzbg7ttAqt
9ESsRC1ABaSCYkVIe+NCXJD18qlZCK+rISrKaBra6imsaGHUNEGce6Zuik/O3F/b
6nP+LQgOOjYpl0F9WtIajV4oR2IPTF0uC/z1EL8sPCJ8afKmXA9cjgmsEZLzLSwY
OZmE/Dv4nveipBLMGo/arIxUeXW19yWp7zz0/aqGcUKaM27KfkNkq91OJ4J1RTfp
zDu/uTNAZ2g7NnUd6flapgjiwD9NmkJDmTkeRdxBeOgSTZecu1Fa5+HW5CkGwqnD
d9dDTUWhO9dMsvFSmAhBLWbeqQIkQ/EtMdlGuGpCoFM1W1xyqvlJyrExKS//18oK
YwMfyxNxZclZuyf72g4mBfU3aMHsSeYauejPVbqRhTMcnsSHeeV/dd7n/dJWJ4u9
ss4YxlQhVpCiXe25CwU89SYbOHWWsSQRdNWLz8BeNZrYGhs9qqxjUcnbMNqEn2OA
wzFdx5WOy8PMYtHHLBDbPaLB/CM19rKlg840inuflYLuUUb9qrTZdxvwoHA/sGQS
fvFGJtdCRiemCwdcDS43tuXY3BijI4xNQSOet3sLEvtimXuUNqd+QCaODSQV/gbY
ro4JvIU5zFGXmKAysCJ3u7bBnM/YEG4RCw+ZCm43iLWi+eJfTswalci2kSB3TNrJ
1io/kbYmTXLn/RvQaftXWn/UDQ0GKfLptSt06Y2hGY4pyC55G/FkygrNhu4PPg1n
jDQlUkZkdupil5aDHd8vX5TLyrgjzd4iaXqej82ldu7CXmNlc+ATO/IIxWfOuI4V
OV8ajXKBMuWTdtZsMlekMt7HtJLhcsLxVahULS/9mH808ek2zMWjezTHlYFy1c/C
aYnipz1VrOq9oBtlZSRryxU6ZBfnBQqYDJK19WbBQBsbr40cm6nW2lSXPikQ8XLx
X3VdDmBwGPMRphSvURQddmqGAunwesl0Fg+5QG50T+N+LAxNLf2vZXouvhS/3IZC
Y7sRSH/xD6brEjfzZ7Xox9c7/ic5TeKHTOgfr/JRRN6SV9L3vFY5Ce/E7hjy3V7J
mLLAD7KIlBPgjQDVlzF9nv/2AV3yds5Zfy2+syA4eLJn1/UJU0zaKXzn7O7B0Qr6
E/V0EtoTh2NWsI0/42uT+2nVx5JzrTzE4yFrBNg4REfroT/S0AMBfBT9b5NDnvo6
YpKB6NH8s7oX4Solj/nhEYynfMewT1m5lEDlrckjBuiv47vdGVD9IPSLCdnGsKmA
DQ68i3MhRpHW2JDkOu3VitlJ8gsMCl59l5wSnnFC+P77DiKYbkZbP6rLAltW8hcA
NFB+3XA0o7vpK4oWliBHMnb2O+Z79N5R0lqim/ThiuPrGYeQV9whMWL3Ez21r476
l6nINYRrA5+/y2Z7NRh2XI6FiiLpZ38xY0no8228RpHmWRN/XU2Gp8/E6DT2gNW4
fpFDF9+JB2fYTmT+l+A8LaoFLuPwgSQ9ySmIbYo57T/g/FO9IHQokc2vP7JexsTA
tLFI/O58T9dpfo2Ay1hG6IGqklPkQIQPwd8dWby0emyoVE5I29iEjjvEKmpC5s6p
XG+vHHlxRGnLiPhlL5sXU14N4iYA8XUgXOyYVTVhZ4yKlePZ+AS86Bc4W0tFJMn/
kVP/DUMUELXWqXb+/1zcKFhUOvF9NcHNpFPKJVfelQfHdn8FrMY9o28ykT1mh58P
xc3RWaE6Ic2ddXopv/TIzOgBJoO7ENYcsm/B1EoB/nUgPUqsnN2cOh/HKb5jZYtI
lWpH6ZHLjU1T43Q3aimMBqNAkDrhsfpmJruGe1+8pgLHPqIUeyVyjvWMZ1mGZMlO
i2hOlvuxLxB/pFBZQrJY76vedKge5qKRMpfe408mW7+bIiwef7ZOYhB7I6GXe1Le
ciwjmCfvTLbauaUrqlojPZA4JO4nkC4Tu+0Yr+O3zG1QMegrHTlOMmTyLSSAtwUg
AR1QU+Pw4dJXZuU+5ucB/cxZNRumKYs2UBj1J+DHfwRLQO268UKS2XLQKuR1YtcK
bOl3DG14Muxn+WKa4mFIF2fjzzorAHQsNmiimmb6WUS0B7PyED3KJIAWSEm4JpdB
HKk6eVbfFL4IHCiTVtcQSkBqQkpzwn/xOR7vVRORsNKj5IUGUbd26TZ8VzycXm2U
R6J/RsiJm2sthTmfSkq/dQ==
`protect END_PROTECTED
