`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9c7ule+rNlQGDt85K3ZjPGqwjjVBuZjVuhuciblL4gvWpZ9554wSTWCo2TQDxDoj
9FUrEBmn8gM+nqUqpo60qcxWyvmKoBfXJPIg3rj1lXqoHKKNjv+AGA3n9DfVbLOd
x8xejQgkEdAHVMb6wL3pN/7QQ1RwH/pStcsqNPSi0jk2k7H1Phx7FGQ2VGFqFH1v
2FTWizBBhW+sP3sJJi82Y/bJzWg4H5QD+N6eCPb3lzoQLaXycuKGrJ694/UZ1DpD
I7nb0NHAq6RmpZB+PZzAUphkk/Rg5KkqmkolOHij875elOpIzcUb7erGPhQh1VSh
oXXZr692jxl2NiV64XRn0K5tmU3EdjuszdAJqB9TNuxjjTBkN2aV45tCbKDx+lVI
4tI7NcaO+OdqwZf1FakE71WbCUqNdjV22zC/9QPDqsTI/AhJMkucW6dWx1cjsk2B
m5xMSRPhH2bridwaScrtUwLqUfCQWvnsggv7e5rPn79bm7P8V78/nWfjfXkQdArk
Q/9d0Ppo93ypzJuKUEevcfZiuiqIDiJPyjy4G2err+2J4Kzuxr816k7KT3TgA78T
cWsZOOqniiNeySlJFxDAeSD53zbTnT9FpNSGxKZK0cXYnOLWdJGvl88PdqlQWbIi
/4auAPgHCx5kLx0Ft3xkd1DsABJrvfPbP4qrSX+1/lcYUNhDvwHqPsAkevYdETLG
/6x8a+Lt9jL2cvZlHayOCbZe+pw3TumJrdMAq13AqPE/88P6Olrv5f8VL5GHynNp
Ob9Bu1/nA6tKhqvQAkUFLuJSFm27wq6oG2FKbPqU0dlYvK3mfQmA4Kvxfve1SYRg
RsarBWaVyGWQWKS4pPFXaq76jQ4Zj4BY9+BezCO29gMjaEFmcaN1fie2CcQFlVyS
yHvECxkRsCiyNpORnifBcc8eaePdUXbjfOrr9a5MesreqRhrzvQ6V9VXyhYr/+ip
dQ8sHb1lURKg+ZcFWUy1Zm4nkiYPVzkrFVrS/rkw392vhK2w36IxNV4Jk+azpXLt
zaTkZ7ur8EIC7hzYoRD4e8+AuYte7tb6yztgeIamaVKJSoHzQkxDwVBt5BF9t4eN
sdP8r0T+c1BSYya0wLr14xejXgu2YUOG2H2142B0DKiXp9gOaHmEOPoo33YOzSUr
Zgs6w0aN8QLA2VCVG3v2tESzCSsL4u+q8Irrb/gZgFDEluRZLyOKGDvekBrYok8z
oXbaISBuVwxf5ySWkuR1nXDQoRgCOsxKahP5h2Z2JkCcHrNbfu62l2/o8ckJvycw
9XKtAkIQ9U6TM0KPp0ceDNqs8Oi7BCMnx9LMIUa5STuuu18aJhKI+pCqmkb44/Yq
dx91yrLztoTbzpvR1GRY7rpoK1JcDIepA+k5sahy0BkbNNDL95t2kqllyS4E6HCm
URBaRi6brvblwyatKy9Ulxevm27oTzhpz5ekiCfsb/jLoe+w7JmgtAEz9/2zs98f
mbcOHwZFhTdDPLuniR2pce8puIyZiq3i8MYc3XmvFsovYlNkDHQNh9dgDmvzyWvm
7jh/KOpXuULtEl55qp4OCIYjLqBsP0kgQ4vFHlp2jJpZQnohomVvhEcX1XSolawb
Fg3DxLQHeHP9KV4QCjLSOw1ATGbYYRQye+7G79uRDtJAS5JvIg1R0sAHukr4xPBu
sPAq30J18EZjwvNE0QXZZwCK7dgAzqAL92xVN/U2YuZJEHZxPcMkPiDoQdMnW0AF
+v69Pm+0WDJWQfSD/vKJw7QNDe89q28B62EDTYL6OkZ7nlMwZivZ6VbZZ7oIwh4J
cWQmO18/dx+biYSOd2bYVgGOqWDr7mfnZYp2ZSwBJNqjnfsw4NYhXWznY1L6glYX
OeSdY/ZWH/r2/vj3tZk4aGn+TrsEdORN6xVnutxnwalhQHhl20ThQpBr9U/hB1Ku
Og986m85lcO7TxdYuzBWHMiWG12RawhuUqUiUDAI3GWsY6hZuanrZwB74W5rDODe
YH3XV0uHO+JaLquPChIFiKKwkU9BHSCKDR9Um9gJL9eic3bqpTDftWpd5vQ+SsWi
KtktV4RqFtLQ7Mv6uQU8bwBERModRJPXf+sknRhZskNiRE7+TWmylj6iWQXi1qAy
L/oVYgsWy0rCzDH4zTcNKYSBhwwPH7aGhMtplwSkO45ejuCKl5ceWVwMsAAblRTC
nV6slO4rupt+IJssFmejzD7GgIeLWBVq1t/GGAi8NkbL7JiKmH9VQWO7GH/84dat
Gra/eeTHw5Vsb2Iz3SQhisHygxEyp1v5NnrBVH9hJvqLM6QHedAOBxjdmcYfHdo2
OsZXNxCa9U3dVmuYLwRNZXNaLn4qi82nYcB+ldK8H6A+A7DHuO8Lx6cJuokpytCR
WjPN3e2jkSDRfYfPZr4Uq76jx1Xn8PbeEa7693YZemYtUdZ6nzTE3bb53AqPWwm5
Y1x/AfSMwJEyym1jhOl//Ujln3XB9oo65VFpoEnbwYTm/vHwJkZZn49X1UpkTYz9
1693LbXYKBmH5LqNyyJcZTdHwRlMkWswud2P8wPOdzz3odUmU7mwHcfesI/jmSKV
HumZTTUk80HaaeVbbFas9A2Yj3kHsDSSQdCpihz03AC3F7VDpAlAj66JzQLZAL2B
h9ZKtdmT1Kj9N2kXhgydL6AysgiyBP7XPjB59e2av/mxTDZGaqJgCZzxixPNxe7P
AJajCGJPvYwArB4U/BG/H3o9y9K5Knwk+sUlzp3nfIrj7V/DNjoumws9VzAR3juZ
S56Erg4x7D4mMRSwCAJx2t/ZCIFszs97HioPHYjYE5zbJ5R9LH9Bp+WqSOnht+3c
c1xUFtcqlb3o6FDChc5igDi2h/h2jgej+e8VrU6ZluN1yZ241HOlSe/U1/6i0Vci
+z9jBiaFZMg2e4Z5qaR7On3vMNmduVpBJxOE/q9d2Syapy4LwNfflsPU+o3BnNhc
tdvljBWf7EBa0btrbylQ8i6jmGvz+49S2HluNCpO4kwsIqovsxhd5cNodhspfuWz
YkxWc9RaTfSaESNk0w6fFYAjNYkAcZ5/t6HJ6flo3QPBLkkRfrzYotfrIWleCmeK
kdjNwR5An6+z1y8651slXuzy7pOL8bsvvuGFeCjE8Ljfwr12fQ7bUf/7X89Ujd9Z
1misA1pwbASD4dGcPV3r41OnuvuA1JadbHxieR+yoXPXdBiQRsW6GDHBGmyFWJfS
TxP1ahjkjnsPUaHk2xaoUYm9yt6niYbYxAc4R37e6x1KWJtlX/QOsfqjsXYo7mFw
kE6i5m6dP5BhlenRlH7Mk9CabandCmJHMcKiwck/gAsnC+6/jy2kCycBFYp4sV/6
oUFBEvroYALEyNacCethOlLRZoxZKbVyq882B9FEPlrrD7wTF4YlZNZiDaYuKIEJ
7+rVqdm1DHSYXJTdOs0jhoDUebIQItaawt6yBQlZjafeJBv1QRGUmxiKVpChTIwb
E6ABDbkBrYml1HFwdYNpgo55g3MYHI7o7Uhcd8YS+AJ4Mr5AE7IRPQLqpRfNG2CW
2ZbADAwlE5fNiq8TCqKEYbmcg2enfEDoRsLkxUFAui3ACQLGlre86DQpOFdwGxAe
IIWDtME7wqeJOoLHiIhRL2SfvegakYpU8V6To2qDQ9LYJ7d0/uo1ZLjouYFklk05
9gvK/v0eW8fQLZ3VjEAFCNVZVxrIbAqzsvl7WNdKCGk1vOG69ALm17WmTlRoYW0W
Ua4niiUt4fOs3eA5my7jRKHBUmr/SUjKKitHTZBaw4I0Dqd7zvMT4dhYFZw/x2n6
zsONloaM5ufgXVxhruUfKF+aRcj3kftHAQOLoPFKHCOPFC1GP3a1nLNs5feLKj6t
RKLcx4qJR+vpFqfc4HCt5GkW+Hyb81XUYSncvylvF2AFXGPZl2/Y32cknweep4zO
r7wUYYx3sS82h0GJKk7oKcTdt2shU29cfNns5hbNJKNKLC6mQVpD93UH7iBmaXT7
xHBO+PYb9JyHDWIk/VFCLctLSjZ2/WH0j5/U3HggcGNpaqOeEyr2atpKXKCIBcG3
eRokhorBVcl353gZh+e1ngw27JzGRsSH+ZznCn/YTVteV6uIqqTI2wUocq2V2l+i
CVJIIwPbYiWyiVrjPHtW4yPwUM1u+BL900kbUpIZ1v/jVxsYoGKi+GjDcikkGfoR
ZYBNUlJPFj3e9YnY4T8cScORLCEFF1/7Rzx6/cJ+rZlXqVUNkrQqO0A5d+bCJc9t
uC6La9bu8FoVPRuWsekOfu4yW0oEHWq5SNWijb5SLYOnXqJQSqoUelV6S/yZzY4z
jb7JQvu+P6c9kr5KZDfbjGibBeOIWBDqo9xX46PwBjvU/3QnpMUeJPSIwlKcWIyy
OZ+1ABv5aQ5VFvEMTZuydIIg1mSYTiRunmf2UwEArkc=
`protect END_PROTECTED
