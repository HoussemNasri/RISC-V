`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VRSQ5fnZKAdSfc2vX9WTth5E773w2xRPc5OZKXuZLeSoeax/yp02LihA5gdrUjj5
XTiAgpCR2u6//HY498qMsTnEt3sbW8LpiD6npiFlE86eC9emkn7Hoc6ddwZG+YIy
EHQ6hayF+IXJWWj8I2Qdnm0wzh4fouRpCKYsm7Z6FYK0KfDOoyLmcVgqrWkgHnA9
K+i9zuZrsEVZBs8ONJ2ZtIIhdC7EhTWcVej3hY8aAHIXOeLGnkKR3vQptPMtnshH
kZrupeKbtdZRsDV7hZ2XH+DTyOUy/rxZYoJwXAEw+SmcVoe7mC15HGO63eVU55rw
hGIVsIHC/dclERhJL1AkDSdmeJ0jGNkFw02GobAA5IYXNoOAuVUwUPYB3Z3b7TBr
WUXdasCrhitC9+SU2LAsXr6MQo8AaLCXD/DB8lCc5hagdvck3moI8ccwO15pcB3y
SrjSScZnW9seA4GjDG/KI5MxtuANSkyUayFWHZMhYNRRVMSdcSkdfrt4CxJfH5YG
avOw/YtGbl39Brncaqu+LMzZZJjMqQrYP+riFOgDubS9vEdf08qkSIhiBwDg9W9n
68pgZaIp9jewgtby5oX+z0vcQbqYZN/CrnAITAdP31FgPopmeZzvlyB7uxhCz5JR
DZrud8NwP5wvWf5M7X4PhW9+vi1xidClbGiffMmTZvqdsE+YTwU/D27FZnnJVsb6
DL7OYLtnFZ7Th4flZsbUPe+jTf4VjwPprHiPANZqyJ3KB20ShHWAzaI4/e3v6w9l
ukn4T2DlN7mstnEt6ECoTvblZSDoWI1hudNZQJlneTB3xXsiV/SeL/+k3lItVX8L
kIRzfDuA9qcjK4dVcQk0uADdHELAs/e5my/i5OtCqt4=
`protect END_PROTECTED
