`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHNT7980HN+vBoU6Oz4zXNURstCeRHIKKYFXeVVM+GbFs5oylq5w2Dqewe6aVLYK
SlsVYAveY8Jy99Q6tIP0xuaPZt35nz6X2Sj8zP9C6QWgyySfpY1Jy3Urlyt/vDvO
G2ksBtNBCt8JTaMfWhf8KcTUaA2EQoUKzo33LPYQ09eQHf6ma0qEHvjgZMXdv3g5
kFFtu+QXFtHUqIWH2/SwMu1Tg5N1SKCb+XuEQzESRhT42MjzwSERGDSCD+ezgcbw
lXDdgr1+OCi9SyIJE5/UWMZW7qE8BPCwTKhoJfDdBV4mHoQdGratHtqrM6O0BoQJ
vMsW4/6rD7T4W5jTGqA61PeVluQwCOvYkx4gCPrdDT6twFgSJWvQfMdM87DFdXir
y5zPnT9rT/2QkC0uEzIJVWFZxOEWmHRPGScKKi85l9AXknhVAIfhol8T29x7O3Qp
At59QD2TiBKVFhFPr8fDqNOcyZDpfHTVFHkSxS3aI9TUwmk+xDKVXA0NzBoGFYiH
nhafTS9SJ06pbaPgl6OnuuKhglwBmHymgd+vcFVeTv7CtxouJ/QvS2uYoPlnGSU6
h0UmRMa2/AoEKyMaeHd8wkJOVItQXvdcFDYdHhOJLNxR9D9sUXpeP15LfqnRAUh+
1jksN/Pwa6asgxxojg7rLoGQ1IqyEL4HR6EWxxcwput+fdl15RjXklAf4FcYc5fJ
9MA8svk05K/Kmxac//YaiTMatJ9lzkDeqJH7bceL3ppUBEbCtIBuJG/CW94Ik+ix
W6n89STm+kaa15OZkRsYHRh3r4CfelWupB8KtXSOdNRAUWSCy3zpWTwEteBn7kTT
s6yUhufYKkZEpUpTcF1bAlSGkAL7vCU+eIJnJnEdJhMPFZmhldWAWO0dL8cIVBrw
Ls8r91dp7KBZNvzrN7um2gpJvTOFetMKDrB5YPBerwC4h/l/5w1GxOjS0YOW+s9U
Bh0gH42tyBq1anmy544fB6dS8z5tcamZeCudwx2cq5kgK70exyCy0dd2Ntd+e4I0
83z0L1NA27Ojlbz7n8JUlnDD5ILHwVTJpDpKjruGyGg5/SedwtY1qQJnZ0dmh8vQ
DhQr1TqJorrPDFJmYP2l/Fw+d0EtxNarcerq25Wa03yNPwgWoOjhs+DFgfmP4N83
RT5Bvs5553wrFGwBfQcJDR8H3AAt8KTNk4Sn3pOJI+6bVTM0TNseQTrtK9PRjKJ7
QAqfN6K/IDEYtQr987zhpZJRAhgJUim+6cwSEpLUH9ygv2vcH66H+qzThj3YO907
DfziNV6hNTSTrrXyHH+r7O370eOEwrNvf82ad1s0u1b0xfCBycgtrxPoiCjHln8+
XJSBoV5myMyk2q0beFiMBJqvBnhd0zw9jnigOeqTdksGUZac5VB/XlttOv4XUyug
OODYVyWluA6P8q2BPGTyo7u8M2T57K2RAYibP6Qci0OXkklySRi6aMHMlpQruJ1H
v7lCoqusNmfBWfqmjxqnqjUO8MLokgAYBUgZB98fBxGrn9jbQJ1GzjQkcgpKur7Y
X//RgkvECfYyAATSvcUIySxz1KlyV3Qt/uZxpuuJOrDoGSyqHfpz9uwO5JLat57J
ReiPXyBoChFsadtygCw+ZljqnfwnAoLlhg+bfSg19C7xRlQ+UgGKJqJjI88pbmR3
DUfbYhRQnYEwS6GgbUMI/8ZDu6fGeqprb3Q5QGlY002gdTVyKfpPJvjG7LfIGRGa
U+rcQtTXFXoDWCQHroEGV2uDEonuAt/jNHEEwTIiJl2J59VEh+WGTDluzpgDdu4X
1iXQ9xwhCkpa//0mZHMsuQm13CIvxtX10QlwbFcjpstWbhbcIow2Wu6wNjB53PXZ
yNW0O4DOZUbM+KcpN/WYUdxKST7LBKU+nGeCgsQviRfIv5iIKKff7+12AghtaiPM
uNwy00eqBW+YwHOTQTcoUjHxHIzPPR6dL8NnApdjlTl/Z4Inwqyxi1PoAJ1tXpQE
37JApYOiNHOWXnr8nFhjotcDDmMB+Jo4wPoj1GiOi7+weXiPSYTLgprC3N1ZK1sQ
8MDphfmOFIAwsjhrCf1JHIt5LjjAYN4f8r69eaSiKZPJQRCo3B+jEYmDz3d9USEX
ExmZrEvQR3VTjBbOjK0H9QHfwo2GR/elu6+8DrPnhtVkjQvEkh7wvG+/Ws1F5nQA
gbjB9xosd99jaooQv4CoN2IbtXtPaqNa8zkEy8qGy72sNTvaqz8KNbYfFRyvtJO4
IU6l4VRSJAK4HSt2LSW2b6DBpwFYmLtLtI+RKD0RSf2gkjbJ5mSUS3ZuK0sSAU9k
hKGDMEdnOrlsl1KQESiWIpWqm9fZc8o/7VaxrYqRHyZY59Cmq7JgaC2Hz/+v6TOM
BnO1/QxukS726G8JnxOTOQ==
`protect END_PROTECTED
