`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFaBhfoYgzUx8rTh540hJAIaAU8LxVwpDOLiD9RkhT8PgedP394q6DBPfpprhfFA
UWk6guvrPwsxJuuvexGiBqSf2QsMDwVRQ+mTrAzJ1n9Xr6zR5zimhcZGJfvk2Np4
CAcEVSmqqa0mRXCiaFj46glpfq4zQDgielJToTcidTEjcb/8nTVc37iperjk2zRf
oHNhIbMICxguKvwBOM48jKCJJiJZSTJ133X4PFA5CNvCTCg59DIGy/WdIQm/xFG1
qG8LxKpmuMJoMc4z2ezeV6sJL8JQJn0M6ur0LeZx8FkqWEQIafAGAqMTsm9GcyVD
MedqsVlaHytGNZaY5MVPnlOeeuO3CsXco9oXGCmpiOpqyyY4Aqr3ySKqpi6OgnEk
dswOltaGQzeqpJyfmRQEWLJ8uRBsBDmD2cfkZ2nlRNl9Hm5gGxmBYPvUtBZj6Qq5
PL2JzItKpQME5Jf2r0YZ6oovLymNzPXHtA1PWgIY2muwzAnVrlBJlEnye2ZODMWe
RXW6dMJ4LSW/kCsHF1KRtlMgkTFA6yRWDrK2UqUhEqBRe1SHyZWjZhUJvPPBwPvi
MjhSY5c3dQHTrp5iDjkxE29lkPVV4eD5jaD8t9AM/QnQiHuy8vHCMiKy7241TCzT
60XD5f7hheG6boN89gzaU3o162kV4QMp3EQ8V4vm8s+5dvVatB5TM7Knwb9pfRM2
pj6XsQc/T5rvrG2TrGPmUdn6efmvTtsqi0fjDpz2Pgb2ipga+gPNY7YW9XMJJZ0i
yI5P5Y3dFT3drtpoo5dv8hSJdjaGHkXEGsOeovgVdfUQ1M3wD6N18mg96krH7lRr
pmIkqhhRXfZYXc8umgEgwHhWseinnnShPEuLcRuwMSvxHU7xmNxCh2yb2newpWFV
4hzkNekGMXLqvhmFUKZQqyjZUwBoPUG8LL5Clxdsocewiiwo/ZEx3GTu0LpLbFhI
+HrKJ5AQf7sfybFA3m9cnlZ+pTH9RTg72Q8evzAp4sORnYw4OZ5QpIs8MLEtK+rw
pYvtTl0HO/n0P5jhDjHzfb+g/cld5bMib8/aTR8eqsvgP5d45aQu+NRtckfcsvtu
7LKG1BoChq3j2Lm6wV5yXdrbkbJo+X4eG/UDvLUseBrsECqQlOd0fh23KHJZJrJN
pVbk6xoVf3zz4DaCkIRmKaR6j35e9F0i6iYfqRuHeZNr4lYziBlcKNtZ+ZK9i3kf
m28fSzUwGKQ5Z8l9t6PIjbFbOdoZQricBzsDtJWHBBI0GJSJg7BGCU4jAd2vb7Dp
BHyd4Gc4hCQVjzpwL0GILO7Go5p8tyAjswbG1PLVTXRbXAxlvwFYAa3C9bKnvJX0
vi3WRtzo9DxF6ES9JVzBw+6j2Ojir+CHPs8QnUdS9JTb1Sou9V9haawMVgEda+R8
TTb6v3qbGsaEBmACVoKLZn6s9je3e62wSc4/MWvIznlHj/285BqKSeFn4nsIk8PX
M0JX5ItGyZ4QCr7yby14IAX1wg2DDVriUYB4+W5A+8WNzGORSSlWybHkrXeUkzA0
/rrIEZDi/Wz/WWimljoeTELcBPrbaGlHJwdvhYgS9BCjE19vSmACTfBY2NcFd5gQ
NrPB6AsLvsejNvh3BK04ILQy4a+ftxq953a1bAfv2tNu89W+VplDe6+Wh/N8rjRA
WmRmWa2YfF06NeIFyWF345zdesNa5AG2vLo37euXy0B30J4CTBT77imq4lsC3zc2
f9d1yo6dNBCe+0v09iIO9j7yyC5RWoGtvkQukLudrmVdVMuW3FDLS+lAWurQoGSE
A7ujajOGIzovkuNUEgnT8BJkGxNT0UlTJieVWUqoWUzo0VxQeSccz4VaauA/sfPg
Oa5/+6FxOQl1WeoM9T6HsSp5HNZZ+0zvtlkw5wbvSyql7rqlUTJqZH4SGedwQtmP
sPLE6ilZlxnPRfY7+QGcX+dZp+FyKLcgYtWoHL+TJKtRcZzsBL9P6Eca3R1kLWbh
3eHKy/L94hjx8jnSfM+Y2wnf/8wVPBq+6ezNSVRhZmSSWXFihdmyKYt9FfZjj3Q8
9iZ7Oz7QJCJdNfeYMPNv870F+VXf13ZnerOZQIsYwVd3uZx5FnkhosgVDNquQa6V
PExpBmrT9EjLSo8KOrYDR/oE7DgLXzGbuCHPmyWNBbhKuWDDJKTiKaRE5S7garSz
+T+BEiAC/YVFRsWSCHfffcdSlx9t2lu4/wFGuPO+RV8hAzmU90W4PFuR98Il+Hbs
317OV/LJykzYOTYOUix/0LQThOmUwsCY4WStPzVteG8J80fK/ezh1mnuwC2kVMJ9
xu1Iv44PiKtLP/69ppn+IgOOeWxf6pIZnc+ZRO2pRx1t7CyrnHve32YF77QQmDS5
bSZZOS3rzIidJ4TvxAn9x9Vr8K8vIfnXSdl+Ga6ybDxCzPyhBl9+zAz1VNYVTtmt
YkDN4sEsdHx3KWlunlKOLIokJCHdOQGJKyvXrztbGXc3usRisXLHXAUr3ESJg+4h
pAyJ4AkedTWzlIcl4EmF38p1TmzTJUL7ge5yqk3gxsaXrSzeV56lZRIiHlVqffxS
AulFvI7iYHXeyWCCwMbw0QfX7mwpWlQ6dQhQKy1ubMW6CA5zBQvPhZ/pP/C8Nix8
brUupiyVM1FHnuDNNnY4pdfKCwqUmO1ev3Mqw2Mv56vG39NiCDfw5sXK5no+c2lP
nxy05piNGDy4TQZZVdpHEpbxbQVyukXnCc4H9JDbHNJyobkoFwi+P4IZO2Gm7hQV
mY05vSratu/vRGnhegzYB20LGsY4yC27XrCvWij5Aabn9E5FJraYO9iOTGeBjVxI
vuXx6nN+TZl4JQ5FxfLjje8gw/PRK4+gp5WZTIPXTsawCmqOf3TxN1uQNmvnN7ZJ
PZg15605ZsfoUhqkc30wZ8BegGzb5YxLFUoTBhVpqTayO0SmW3MAbL2hwyxaVM6v
2Zptkr1kwzUkw5viHXNwDuDwshfQ6CkZEnSYgPWgYwkOFOcYEVt5jIjLroOh/DHw
oYYtsLgFUdkXFIW8K+KnzlgeM8JvwyrQ3ddlIdA6j/WnvQD6e/uj8HIddQKscQEv
zPMMnjC0L0oj0tAz6JT3tYWCa7E2bUN053MIwocU3WMsiSim9RojWZh5q5DlpjQ8
rDGeP6XcEpVwtP5cLyEqcAVtQDECc82A3QjgkoMGHy2wx6s9RvuEkDCFi2cXky9z
JiEAAOF/J4066nI6IDVOK6YO6zWkSqWr9A3ra4hO8GitzYaS+8ZYuEoaEhtD5VIB
UEtPBdjZozKwxratWJ5rLgFff+xVPCGC/WU7e8JGx+UwXeuU1+RD5OVxgrGarM+h
vo24EG4NIu3F3HxBzvglrELIvkxnvcaNZYKPrW/I2ZNBm0GLTzwEvOaFJhUrgOD0
lf+r65QzPw9rwHD0LHMouZluxxO0S9eD/mYIFYG1nk5TsN1LeGur50MpTqIkYGWh
G0jme8AIRs+eM8fYd670q4uP0aExqGjWNzQJrXyhjCURKduJ2JCZxVq03qFrbuBx
/6h7ghpCsMBjmmJXXzUsb1qYiCPMJyUy/URO4rUCCyIuJssRBJe8iaHbWa4GRl3p
Pa72LLaV8B/lRiCNLHHoOEdNqdhvg48L/j8m9mJDK8Xe7ZX/DpVFrX2DtiBx4LvT
f5RPWu3ff4aqVFOvjHc6fxSuxwygZMdoj8jVUAx7NeHGuWfUjOaH8py/6hcu6zpq
DPN6nEFKUWeV1EfXKwgqQd40yNyvxY9GINB88Tl2HobGBTo+gHN6K1kVoO8s8qTn
LqEvqlZmq8w4qg0TGRBH4E4rw0iqYK+J8Jj2aRGKuSyF9mP/aelT7JzZpP4ziTuB
h/zacUxJDgwtc052nN/vkOf7k0+DrVwoqCoH7HE84aaNPaD7Xsnx4hIw8zKOuKye
0G76UX5fkKjsGPDjAiU8UjMIK5jXhouY6DL5FDhJHk5cD3fYK302ORYFz4qpCnTE
zBmLxqaONySti93WkI62EOBqFujIuMmSTBN02bRnsmEkCXt+hMpAPgEMQXNII54Z
WKZUPUfPKEbWxKTd4SXH/vLTfLmw5QaU7KPsEuTpzre6LT3r8Ylnf6ra9eq4uN4v
MfFaaHF+bhXgkh4InyN3xj3N5shkwuYyJPoXfh2Aa6tawA/dPHrbdg4obtRyHBWD
HrHZKINJzOVjzE123X7Mkfo/Oyzxm0qO8uLsZt+YqxaYH4w7ZRXrASxeooe4W90Z
EtyOjfr4fPXUW0T9kOVBtUyaK6U431KF2+RMKu81EEwcp2k82PpjsIPZZwo0yC9t
RlJLWkrzvl+Fyrul/0BMdzjeOsh9bJB64oD/q8NJILQLzHCj6qOozqWP35kRB05A
/M3ferGBVq59oItkAn+3sNkXrbmkTc8zluSz3TImyDuJhc9e4UZH28/U2NEQnS+v
rUADJXOOwSqtdAJz+UeJaACAEYxDWLq2thLWbj5MOFVD3T/i7GG8cqzx0rKi4pWD
7CBTpVIl29tPIhm11tplYidBAC4oT/CSw/QLbxEmvNxGwnlaaV4sn3keAtFYdNIA
fBY20nuxPlvx3c5Xx+hK/LyHbgXJZ6O3gbawTmd/CgCsxbhmaHqioEoZLUJkXj3B
Waisb/BwCBmwRflSN7EvW0zzwdwGIWkBkwiTOuNclUF1PYkVQj7B9GWcVy6vO4ga
okKTtfcZUSgDX0WrZ4k2p1/JNhhnWNei8yo3Rs549i+4gI64sYV4cRbamStPq3Yw
6T4KvW0d1IBjY2SbsOEmBAygIbtPDXHnlGa00FckouXS/4BiW+pG4meB3FMRHhzW
Y1qjcJz/i3+/r73MMHR9/McLVaq3Mq4ee5LGpSCWEqfi8CkAVLFFFbDDJrrwztgK
FZQW+Y2hWfeUZ7vkWJ+lcMGUp+rDNBFbvkIxlF2mrzXnzWfvEs3ZThOyY7Ekc4ph
2KqMA5fFLcDrJXcl8MO0VGb/PugEoQ+kh6HUbnaXszk5QLd6aHlGg6kb1EpJMoCl
u12KIHXVYxyO8hy7NgC8tDDoz1zD3SLyXa4PEzPgH9rYXBCY6V3o4Dc4LaswVjOS
F7UuxUlnC3a9mZPm93gF6SCmiy8WVa1TLYtMX3S/6cI2BHmQf4JpaCchFgAkSYJo
W27Q5gBtDDtyCyqfePhiCbEtALk9hTBI6TN5dQOjTmhFW/xR+F4p5yM5DqLMjKOG
W74nY/gojQx3c0L8uaBW+KvW/cpmRxK8p9xvHSyJGJprlkQDssUNepQGjrm4XwTP
W8yaNm0NS1agjCYg5uGIEwRwIqLd93vYAAKAsRfnOZqBVVKCpO/QwfEJotbYXZ/k
W7stXgaDlERu661kPZ/AVKt5zUNM6bC6X2t4BruY8H6SxuVpFexOFdlk/NffgYq/
hWrLN6Q5QghzBMG2M7XMSy6qqyZmqs4X2J0MTp0Ao35bdrl+IzEqitdeCiCJgIE+
AnRD4rZhaA+bPA9H3//WuuMgE3GfFIWksXMVggW/c+W98Kon/cZ95EMLwRd7+LZz
sz3sUQU8mvtjFaDEJ5oKmHPlN7jHk4aWUCFHim+5oFVsS8TGWnm1URDwvM7yu5Mn
20+BsvxTxdWH8yHOc+uM77+yXPAOYbTZiKVNigH9/ZjjZa3x1IFrN+LVyhXBz/1v
QTq0v1ILZFRgkFYhlam2mxEYZqwwYc+OCyUKqy6fViLJi3lhSRUnE15rSPJhdR+/
hHY4heQyrEc0WLYq26LuvxaSkXB+k9MRy6/wBpkfF9WzUlUWTyQLAxfnhnlbuh16
QAvqc0QyAtAP+vJ9UjMkFoYaxxE2xlVFU+y/Evg/wQj2CitjNJhjLFyqnQDdkSfs
//sHCvSyomm8VzvR39VShp/q14zhzfSFLwYsxIrrQiv9L4WNr9XIIlo+CtTWxAdi
/j2+rpMNCWJUVYYc02Ypi7ya1acUAQ+soBRkTf9nyG8WY1LEhk4rX/Cm8S30iUDC
S87aXI8ew/d+pYDNpEf6eMiQr2B18iuu1jilOx/SkDL/plE4FZi81Q8DtBv/FSOq
O+cAtVK8r2quWrgRpThmpJQpVxPHaRfFCn6TCuqTRpiaeRKhxMQUW/O7XrN7mN1m
f9A6fGGFeHpdFbNrtJXSUSxNSDj+6yJfo+5ECL+tfmZQTpAuLMKvkmAMpUlZzlym
4c/OjyJBO8ntZ7XpMlUhDnIpXXXI6xXBs9WlMQ/mUAjYPP41GSBKOpWcRCr5jrbc
lI2jeUqGEeK+YVqC5e3V/vBx89m94WeiND+T2xonY1IJTfMEMRA6AY0g4DqZ6eB+
I3DpyYofIASL7gdZ5fLzK3cDqqEubo7dfHX3GlIk1V5dt9L6pvclKRFm3c23D0RA
TPa2TbdYPi82YN14R0cz9lDs9UWPfcD84Exbagh17h8CLBtKjrIgGyjy9kGlrLDa
qGpndFOBoTQCLWw52F4XaFmp+7dGhr4H9FCLnz3S8WqpUTSMEbvwxC+QHYVUi4ty
RJY0PBgqvu0dgQTJkfo82AXP2vV4Wv9GnX9b+jqN1oESUrMN6FWXmz7ZGHDBzIA9
gjjhcrKXGz/CcP/6XwTbK41SQPo73o7YY1ryLlL6jdwXHpygFS3A70kBAqbgAFUX
LvkbG2QM5acKTXAKpgSEeDwApu6Mx5H/b+1wsSZjvSVccIM+2gjVrshUI6VTJ9wr
osT32YxcOg9gk7UpR85Jb6yCzIXS4qtIpR8XGNnHeiT2anClzSkk9GkcnWfDy5+S
08XY2qQFserIg84F5RRm4vb0Ss4XB9DH8Fc64RSpEkNZGHcjSUOcCxmmVyk0LhEs
ntFtwRnRBVBR2T6tXlxJVbidn/nTQFinB7ygTQauMub6lkOUPGadpFha2z5L47+C
0arcQnPXkVFL9ZE/kSN44p1v9rLLj6sepRtKyBpkZi56Ab8w1ISf1Zq2+n/YeQ3Y
UvB4girvxvEmOyqtFaE2HOgGeyMZd0LvX9mlQ6mfPop1HaCcs2vVG0m2Crzi2RU4
cdpPI69M5b2ZhbgkACKCbhy2G98iqiY9yt07Z1WGvcVGDKBgmxce/huZLr9pItRC
9pB/gvmX7OYYNcW35QO6KkvGu0Yo/JerC9OhYw8xCYEGMmO94scxJnw5qw+CTCaT
6oYYaTRkvmZgECbl9sRzmTqJREZok7j6nPRSWGBeIdyAsN6ghFF0/IYOK5wEcsho
vcuArYAG1EwjjygnFmnUCjLa1S+XerSwzmPlSxQbw42hHD5vedJntEQLl9xCe7vN
WF0qUh0oi9V7KpKsUiSh37kzDCebjP6Q/DmXu56F3qcGrsoqBS0E8VHYxDelnJWT
TuYWM00nuESuszbR4YVbBWO2t7d6f/1e2x/7Y01W0frsP6J8plU8ClVIKzUamRSI
iXLSSCBGeKQdAt0JzhdJ6KLMh/UZuhWhyCkpWXFIM02zy489B2GyRFuK1DRzyMxz
+EfQYN5itP7Mi9XvXfA4L2im3Bcq6Tlrk035MUQ/L92TLFZKynT9zUyiBKLmyaoh
TtgkoXUwc3On9pCF4ndrLsSBWs61+/glpXF/su1oxqh9j1RyxbrlVwKu/eF9zzj1
m4KUfbg1LHJGNSKXt9Dxs4WCcKASs/hS7q7apx87Hx4tBWi/tujTHn7d4AApNJnA
/0EV74Ko5+Pb2SzrOmo4XkpyIDPLU9ZDbsnKXOzO5RRg88yu9NUDJgkDGFeM+RLZ
f7kh7Mk3OGQrsUhi9VWyE+mGLUSMFqkmx6hJa6LZLRhJKGSB5jTSWOx11EtChmpY
Nruns5qudb4P080eT/ypQYdBLrZHtvQ7/U5fLjjdkVCHSeXTbmE+PLRiD0utXDSJ
XDhsRE4/vFoby2uX82uvAO91Etnj3wlAIjenxFV53Sz7WCWOBbO5tXqlV5PgV+ir
+HYp5aur+17XVQZfd5vQn3EwPuhq4rNQZsp6TMco25C3Zh30H0dPVbOriZuppJKw
Sd/IgxcsiZeNuz731hpk1CcZEEICfxRP4lduRTGmlzwn2XAGzCwL3XmMN4NUTR6n
uYuxJSFRYKMFFl/NjDA1pjhKL9enfYTsO0qeNKBkTIEBBRA2ETObbryAgG48YGfZ
+/9PGwhVPtNAEEqGT1YtSw3MLpFT6Pbbv1zi0CTvzODOnKMN5+BNcjMPENfiwN6N
LosWSzLbp0a8+to4SFtQ70/Ex5B2GiuEbgNPDXfjWTAnha7qD0dNp2qw+Mtsd/sK
q5pbOKtuJnrGBuzFYxuem8h0FMBfnCrZHvo8CgAikDcBmdVbWQ5oXHG1oajdWv5t
OUoeRJWYAmJdTj17eBsWtJE4o3IGyDyyUP9InfYgCK0C6lYVjfARPu/zVROLTI7C
HCZJ8oU0yfTEzQaxmKbrAEXCFoCxcpJKurZCmvVTdeWcQuLOO5NVNDvR1CrOM1UC
PL6EVf2s7qY9ILVPerSsUVxg/FwZioWzTC9c3Wd5PxJrRDHxTi/dFlbH/sFQX2yA
SsM0zcmvND/OG4ApskpT+M0Dx3WtPD4iW4D3Cs3IJi56RWoHrH1H9mxXMaVqdqSh
1AmY1U+yPXgxZCGGc6eDhSAZSKEZ7/U7wWFxbI4IxmLlObQ95a/H+jHuUp+AUtW1
R4q3lgRDF5B8xfv9FIPiSYDipC/46j8o0RsKpMFWDawNSOSPx0v7OHC50x3IWJDx
VoZDoX0WVGshiR+rOjLdqGdP1iAFAN1vqHU7Idy8pA4yafNihg0+9leAKLfU2OSg
6pspZfVe+qej83mfvQBYYt3U1r6QXKmExJD0oEECWNRU34uCjVMiN623LqA+UcQU
P8J6ZpAvqGvvvxCcUZojF1alBV9ngzp2Tr/GLT/C40b5lTuxcelUDK7xx+P5QkH0
XJfSoNP+01um8RvrGlYeHXftQJs4XGEzIrvg7mHMKvNiTDY2Y9ASiKDVIgUcVSgS
G2GRQ3akq3o1dgGLs/vd5jkJ2KoJ4HxquHi0bkVg2c/kdOjCWnyUqslHEhtzkF6t
zuxu4MWGoIF6zy5Fk4mkxRrnrx4HrgbOLS+dpbz1yHzVsa1Y5lYvQVy4g0/3RufU
im9S3mZCTMMsoErOesvMrFr0KFHCUxLYgXHkp6YF4hnnz/aiJ8+pSQsGKx4mNKHp
lMdAkxhZkcgFsyCRbL/FV0ScT6RbwCD+JXum0/PXEUsBe5gcL/QkfUZRA2WnuZVL
sCFl/D6fHrrI9rQNTM8X9CyL/tw7h3riD5JYstMldBrt7/4FppqpUGk05T+y8b94
hznaWt1Z52riUuOWDs0LLRTVKX5KD2k+xqm80m6FKrx6lT4Soqq69oYbyoHUJz1E
LpHzHqQWSGTRR8IRjxMoL1UD8WXhg/MReuARvodkOgQMbiSi+k3/LIHp6wSrHS+g
UxH2HQvIexEuUMddJaJwwiPpkV103ru99TPH7XOfhDAPK+M1RUVX6Ww0TouXpCvS
+GAXIBjtw38dGNLXk0wfCCH8vvLsupf8apNUXSxYrTFDBVnGbF5dbGnhnjGJrvhT
yQjkLClGDUIRaKSyfncmBNDbzPIMiyEWkJBmOGPS1P3DFS792sQSX53sgtIaFiK/
Tvco420E7H6zayKtTXYyHFQ7bWiKqCOEgEk9pNcxwZeFbXQE2fyZEmAzCUiFY5TH
vWDgsn7F/5B+lKGKmzC/Hdm2xJTO+/DNoF3jOwIw0P3bLB9vCpGEOiMw0FzgfzZ0
ruUZARw193t8GPUFrGnB6H/cSVslahQFaxHECiw/a+d+a8ZAjmcR/iRZjfejrEIU
DPUUbKOgjI9ovyR0bhkn4z7ppXLi7w98FNp8K/59wV5UTmPu7r/X308nLxj7QI0o
v/ZCo0Q+WKDaC8+Y11OufK+H6D7rltG8rzTf1SvDBCaB3l3a2k60R+5R1VPlF5N+
1dFCC0cOWCeDO6B1O5mdX7BCmw0HTsY22qz1eHFNFCEDvkmVbglsBh864LXk76Br
Q2BPYfqp8uZz4wOTIRNlLkv1+nboyZ5HVu9Ue7GzwunUa1sXV7XeWrLD1IYYOsS9
A6A6QjT2fZXuNj5AAG8AwzJRmHwnxnw9yvslcZzG7BHTEBr1U8x8qNStCh8+bZfA
Wov99rGgmBePEefV5z4lQttP52qbUVe+75QDEytEDVlyvGyXUAVVDGIhKsvjIbd8
1HPXLIPDb1bJvgR35/lMu2quzvs+azJbITvEpi4RNgIKnxowYK8UMTzCPFHPQkKj
DDv9u4/CMCd/XYFQtu5lpHKaa3091Ny3wEcl04qi1QdLhI+ksRohjtGRf9LQZaQG
Wqp7JzhE85kxRBOT6UYDkaeOyz8NwhINLeQAwLcyxLBgVdWhBcBbxxJem6k9ZpTW
UTqkhSIHwBLma5WmvY9s6ZsRwcol+uZwzz2UC4qQyWpY9O+aS22KXfLv57gX4I3/
u/k4O5HmdoombN/K5qflk+A4OiRkYNA1Rb942nlNSoDn6cD+TfsRFGta65GUjiQM
A97JaUn/SlMQRQnN3H796iV1h4oeIt4mIC/fhRp7OCJzzhihW8CsJMfbXyK0jrvx
jBBh619dHjOHlyOZNSa0s2+KBPSVbCWyfghVLIvXX0vAdNHBgsr6KM34W8lH9Dyl
MH2lf2EkRcGA161BZ8+fRMOdszdSJCUftvNo5WxMEHOGWItD1H4iupVG9Dlv+KDc
NE1ASwc1tc1X6XagNKKrZdKkLr8XacnKE7ovl7ThQWAxncospNpG37hoocSIdWNd
FpfJDm/8EePnOrKkiSTR7N/Wgyzoeejbi0Fwp9UegUu9Ez+hv+sS6XXtImLL88bs
ynsDwE8jMLQMxl0cKYSv6fXqKSElRTKdi0Pr2OYUQknZDi8CO447uwPgDHgiv2Ja
SBvNqiDdSImiaIrXF3auKmF6m3Q7mmgm6dMz0fFHIvjAI7hGWVrJ7/oo6YRFD5tD
TiF202OqnebOV+SRkDmBCasphCr9leHpcgKlAgSzPFBB/PFZ0IjB9WUr2sDUNo6U
BmWXviyiGRNN52AApv2tLPAlogTHf8Neug/fWUJzirWBchSKTJ8GVRC8L0V7x0Lq
AJSgt2UxU92WaBp9wDS3orygRH5EmX1VXu+u6G9Hz73Qf5uWz82in5RM4k8xdF/8
hOdCquWhB2DGVISd06okibkvQEZc1hQpV9ItSz9wkWz6g2z1JS3R0IkhIZUWXo9y
sCtDUE1k6aFK6aa87BJf52tXnt7EQNz+S0/iLXPsvBydMjG9VFKTFOqZpPTOjJZx
PUPJQ0lJe9zmFO3PFE97dvaFX7sesWQq2S22zVN9+c8wdminKzoiWMhXyFEsJMA9
xwF0tGiPbfJLlQCF3Qp/Bq1dNQJpcTKjsN3gIQkAk0DTEd07VvAd2pdn+StF5C85
uwW8l4uX5fVIE6IeZfQQA2lynaBpFiRIgYWhMokSkCFOhq8prMdFDSpLnaq3Vj++
2cI5HpBUS5DIHxu2qjzQpzddCbSZurtH6QD0undy7sGIGnCEpa0WdDiWIgo2f/if
zMnLXx66mUX+U2lCg6C+qO3WD4NZ/FOc+v/PvG4LPqYDFe/7fN1CH0vYYHBk59W6
lFl54E1UBw2EwlexDiKOK2kBcQZu9pswAkcVRhQLIBl1il23ZTKgqh/GqhdOLOjt
LL+/FevGfKTNLPZU+PPY9NclJaFA+enmqXEe1cYOWr61wtFGamSc58VFXUAoZOAp
4uo+SKV9Peqb5E4DDD2mDylNEv7jcbIDJiX/kE8aWr5ckMu4v4DDdYZpFwQWxTT/
2maXYmFUdUP5q4IqJZ0xOg1NO6ubK8wA52TJ6QVls3/wcDvo5WMyH34xtzVDI9I5
rdfy+sisMUXMzQdRaM+iopqlQuqQvfl4W6k1Y8yKX+btkM0uRE8ARPPrMl0YrBx4
CL8MFkYF8lWQDG4I80ZVK5YirWEAIRhUfRa3Qgj+xXs4Fpi+9tLOQxHs09ErUAkz
lTj9tGDGbnvz+7R2W4WryKWTjiHQEfnzggwk4oP6QI1eyuM4GdI5nQR4P6BLf2U1
9/UqDnC5Ke89Wf7XBgijleztKEigYuK/I/WKeky3Gscv5Fu5V3jpvm0Gzcc4p7rN
35MbXARTjf7cP1CXVhqTBKsfcIdWaZh/RR4JneY4vQhIeGggUkxNJBuwoOu+Ue4V
+yiEsvMoWVaL3FBDM4+krMhTZzw5UHCzb9/EYIxUjo3hYgrO6E5LFQ4sKlvzODVl
K9OcyHPA/Y4UX63ib4LiW4O5j9jXX/5B+5KGwQCarGE4eXSjJMlqgjKboaxktZ5R
gSCkQJPOY5SNATuIsG7oqK/BRswI+2CD7lPDwHJ+C7rX5ksVFT2cOjhnieeWU58U
jxGUaq6bTqbtqTePbojcanHe/sXgEDpKn70KqSNfGCdXtIs9l6Fef6o86XUyZmHC
ZtL+7dGyMPG7eD0Ny74CpywuXKYkH/nuO7MOT+Keq7uelBGMa9mDXi1rJQS7DMtM
9ROpJ3AF9fDaG4YIP8Gjfp/UY9/owWSl62/WVOXID/dcwLUWPWBrjlwyzcVhcbCs
GNUiAwkCaYeyTnkZF+KVnyTTGjeY1Fn5kMdKEtAcbxM7k3x7gYifSJF23gEaWg5D
kNozXrqy3q0UiSIooqZwgBH6HpHkktp3D5DqLU6HaXxqOVj8Y9uYXNxobhLDDEWy
OFck86J84qh/v8iAQ3JsDNPnMYh2O8v7v+ZhYNr5lmEPuiefnfhFLosVb7QtPEcL
ipnGK4Yf4KdNX0sJOl2mm2v22dSZC8Wi01ugz/7hFQ3T4uFrYNd+kb0RyRRsgvfv
gtTi1JwxoatEvHuCqrW5CRwCc7mW9s9L+TgBb/3Nfk4xGCnNhL1uSGDPWDuVuBqp
Dh1FHtV9seV8Ez+6R0bC+mvda9DUaqXqJcTcSwkyzv1M/no2X+kqclRpuenYketW
JP0w54+cNCPYeBlUBtDqCBKlClDHVgrHTN/h3O3v07TlZJnvVM8kBujXSI1RHMSG
MRgj5MTBhrlAv0L4MjzmTYc6JmF+f0bVxubusKQyi/8rdxRM5c76raD20ysc2Mro
kTy8aE0seRr0KMx+HzOQC7vBP/bdnuDz7OkG86sa1Nss0bTInwdBVh7Lv5g0+T6m
u6mB1O7VpeABKl2YSLOq+Zcy1M1cOZK7uBjZpj6yZFZlzH6HmfZSCmp4eUD5Y8Oh
7H7zvjVFUzJXDCZVeAeWZU5WBXDbc0dp8NKKb0LZgTzhvTxZv1gXjwDZ2ho2LTr/
wxeQY1zNstQR3bUcuWURTlfX874W9SK8UaazQWzXnB0fjaLtXfN6pscT4ucNBhV8
qihsRsGC8CS2Fx+GKcvCF3n58Jfg8WouP7wXj01RR607dSKVZl8HhsMSRpY4FyVn
/J5m8BB8kuhW8lhII+X9JTByYWXtFaN/8RE8Ya+2RwzVHCyuBQVqxVJhR2mL9ndq
J5Gmbs8Qc8fT5Ckx9G/3Jb118aLhL0BdqY9PScYVYfU3Fo9g5Cu1pOex718XkEej
jYVkxwDCgZ8Ik3+kEoEE+kD6TqrbCV9Ka98RqLTXrokO+iJsIkX0svm92RJ6yMiW
T2zd7DZZaXaynjzpFfPP4i00BUU+h/op2socz2WQdZZc/5rH8aePYOGpIpkJiuLG
SDjoCZrUNNIbL1pac6rVT49lSr7aEWJxJeg8GPEPkrXTVjGH+R8Ok/SkGlALEJGP
CVABP16EekKDRahJjWbit2YTvKnlkWyXLap4+m7P4XPLvDy/0Vqztye3MdgWwGQK
sj1y8XnIKwIyQuhgAaICrvcdxi+Zpj32fF7OUGvPHUo7kyNlW5VwA1uMAq7ua0Wf
7+LHUhgu1zHUIDaMAFH8MSBiyrXt1FUSXyGevxuizpIfty1H8ilseXCvpHu0dJQf
mNYHNPV69Zo//ZqZ1elJrFP/bHxZEC8kqJrEO4YIKi4Rp08gX0Bc7rj0DmqibHZC
h5adXHkkszfOb2Cwh5g26SoEkDBKIDcsQRPZeuBlr9l9biMGFAkFDVIIqaxZPW/7
O7skNASEY/5igg8T4X5QWAahcXjP86fU6kAnfTQnKXFdEr4FWlV07Eoygl6FQX+7
KeZs1ZHlYFq+YRGZGL+LNXFfy6FQpoggxIBBBQl2W+3UovWQ5iIrDChc6c3EB162
3j9M/nv51M+ilI9QlK09531UvBvq3WYALtzef0reTuD76SDwVZJqd17n8yUkYlOD
hLiVnjuDj8xQm7TgIuOTG1tO2A+L5UPuCVPp7oPJDZHY4kEoPOZ2KUa3dvZ9F4wM
CnniQg/imq6mG4AiyWXzS5zAhJdsOEegKrKe2euqr89nT5DxdSTxYqSXx2MqQIAm
bDdIKUg+QwELO7ModXhi8wx0FXNJXsko1GNJFQEczdTeGDXDVy7rVjxWyF+uzeZl
HSd1vMm/1k/bxnTJ0u+sNJguV8nLguXMOr007pOGBfwwumohdDLHnigJEnsVuKjp
YbC7HZz2bG7wRYWhIAg03ZogqT/2GdGa5LqYDuMbYxqlRMpUcLvWSQxZK3TcQy41
86K3JYEuR4mbkXxIhVK7r2nGRswAEgL4IGEfhwWdKhXcz+FsXQLu2S+IZiMIN0ho
ge7MrUbMIIAB+NONzQTdoUIweL1tZsf3bJFKFIiGCaSFQhuXGezOQLuAMjZw4S1R
ZxFOJlLi7IP5sb/kY5l7qRY7bfRAI/v1iICEDUAPwZjnl+9+IIb0lJlRLtCzvDtv
7Ggimf86nypmeG73iKZyqKLe7V+fj2PP7cXVNAB7FOYcLr1hpKpH7/snMnE425EU
lbxY3YeRUm2Z24Y+XuhHoLMdN+S/b1QoEkySBfD5Kphy5wgPjPbYWn5YqtbRYqcX
w+QNGV4FkY+WPS/ApgEcS0N3Fe+O1EgPnluT9oWDs+chQkX5JOapMXtu1upAdmTM
DmMIP7vbC9TpONConY8C7HAqU9VHmDlnPyKhuKxdBrZmNFyIMnPdhgAOlCrjSdr9
Tc3KaM+prWtVudSZsoNHe2xyA5FKVlcRtK8R5tDp1FzQ9+f46FYb7glKfdJux3ts
NML5xVSumx4ls3FDorJYGKaZaTk7a/A/zht0N7oyeLaBO4nrtF4E5U21UKMOm8mf
T3NwTmjftFHQdW7L/fjWiRO0HLSOeYC1bLCa/DMIfccyMSwI0eZweIJ3hAjhXSq5
WvP794NCjssneN8fDLc/AiVm8gSff0DUjs0fVV7j5Mr/cXWlJNs8e90jzyJPdrVI
KqLI9+AnWuspvHN9PUdK7TZL2xkWGGe9our6ug3sB83NQUBfn6UpqmvbzqA7y/km
N7FX4HWBW9N/gUVZh7GyU2Vvgsg93SlaMMOnOqWN/TOhpL/W7NBD5+4D/SFIfEZ5
2dZnN0P7wfqQmoCJ7BLfJiI12TyUUEP+rVQkO1nvW+EWTkp/nB3/+2sLOeArhjct
UkcgMGD9IZ4zaOk07R+s+fGCgzka6ORMlKjdUTEQLz2aRBDGxahmqKwvwj7BFy4X
yBthcuJkKJiHoY5ZP4tt4gebpLJcQYqfvBFMQNfE2Dks9tFXARv3RSaqoORJm+AW
qECmIQx/dBAnrrLMiKeWb8MW6theDD0c6TbRfGxsDH5YPOfxIvURqF4xONAL5xQS
RiNWDAL8Ar0wBDXEcNNKepZaCh2meFdEozvDgbJJ+vuCgXLCz/82dsCjVZLevpt6
2Is6MjqxtJjF0N3uoWzu3eiNEX6M48xcdfUOAH3rN7ggu7buxz6n8Rj7wpElsTIm
8sg3nvJFUWB0rkggi7olmyGcon1LBBY1jYDK5M09F0tZIEm0wCqztTGlS8DwQQSQ
6gp21h3qtYq+je3O9GQZNzjiPiKK4VjDDTN6tbDb0q6Bh0MVo58d978WEbdP9loC
Dx5FBWo7jYMZPDWLLDAU3BEJjmAObAoH8n88FcbQkS1ttnmbp6ces4BEEmgtDxa5
9dHvAW5yEB/xmw8ijLrqy/M1mvcOCww9zFnmi24fMqHCK4n9i7KaPI7jZYz6blrt
cTbRBnmybygtvWi2rHjig2T+NywhukK7tai5SVciYU5LNdkxeYgHflj9oL7UZkNS
qjQq9gvQI1xLW+jfoA1gY0F58rlUeB45DzgEDmt80EY6DNP7s25TgN252uj5tRk5
BCuJnGxkivK2cV5CuHnIEgjFR2/YA5s+I+CPk6c/QEgh5nLz1mIPYNJ15xiONTKq
KuQioO7SSRXBRbvg/adiK2v1iI3QHeFjQ2rqq+f1ZE4q75slz4oqrCGxAjn1oony
Do2+wSWyiVRoruTOeqM7abZmC0rYHdwubIpi7VDMqIUaFK/cADBDyZPR+WUNmwtp
ktqfVEiWC/LMxVMv9J3rXiDjLJNVlYiqH45X2+pvsN9QAYTbKveMbK7yI+/nWC14
+ZIULAKswMn2l9lKiDri5bW5IZfmqOTcscJyOb6D2RU6XnLik9fgs/4daEBrxTTJ
Fa9527LuVKYVPUW+5NVYyCnxB92wrbSQODyiQE+PcteYPFNInntcQVGbK2sRppej
TNX+5A5Jk3tUXY916m8xPJ+Xb0THeRaX0uAWMKGL8JlyLVR56nWRkHSUd9hAEvP4
2WWQ9kAnd3H7vw8yIBcxAjiy2l6y6UjelFa/lTbipERGXC3ftpD9wqawHWFywXvu
V1cPofPjgBHzJKPT8niYOCr3EXnEnfFj+VijX9KTuTcuP+JsQ3wPILxRFmZ2UDEN
0c8SZG3SAh9+s1SENnRl2Xxd8nPd+kV6R+yMElYd2voJfmCWrBPRVffFxAi/Wxzu
3yMcFte1E4txH9kydoMcNmpON7RM/JRyr7gAYvkyyD4ggWDJTMPQOvfiKLTZF2Tp
fXvCJJuTAmenN1BHqG3nBABHsZOYMD7jYWeqPJA2/xBtOa+cRScBZ40t3/ivNIbi
zGBkMSAIr4V/2KoTNARpdP3l4lP+YfB3uSUCMlxNBrf44uhPxLU6IMO5bITSpfk8
G88OTEExbgDLf/MtRv8sfCQb4F1EeMUnzKc1K5Ep3y1o4Dm1dbC8WEi6aZP0rbRa
0bkG84wgH/pixWQgciVW4RYPSbVdUi2CWrV2wIHAvVbhw4sKmcTtwGUbZTVkv4vX
6GYDDp/D2PaFUY0AVP5/T0pc65jjVhSuX63PMdS5cy63Tm9TR7tLRdSnyvvBFEoM
znmNV1nSzfe8do3H3IPzt5PBpU/LURXtviyghzT2q2A4sK7kTu5i4IaAZ0099mmw
kCIFXNWh4eZppRFs7ejqtA6I8o6Opk68LyFSLiefrSMm+7R18ljfV8IJXGzHXxyl
VNbItQjnyWU8C0qn+Wps50d4Iq+p2N+BguUq+huYRRK31MqV6JcJmyMeVlHk5oCX
ZyNWodTYotG2gtmBmoBX/EyEJh0DuQ4YHUuCfyAXnDCvUyDULlzvz+fXytrDfyvT
stdnOKnMEwPw1kTk56t37/gI90IIS3iOQUFyMBDappQbrmATtWQKxWu+vETIw08d
wcWWYt6Sv0mnyareyYThX32PTwUv+sSCVBBVSiH6sZilw+mfS+o0ZTPO2RSH77TV
SaetTFH1XiNJBElOCsV1FEzb/Nn1cH30CwU4OdoyNfuLszlohEuUn2sxDDH8F7zj
GJ9JBWGWuFruKvNBVnRxTsEUu29Wlo5KMtXo4fL8N60nxS/plpDyIZSyqxMURTPw
USB06bNzYZF4OahEjSQ3N7TQH2UjUuvKA545OVF0MihImf4C9s/RImOC3LlMfOnd
txUhvqbw/C5+9oMvS56d3N/xjMpqERctRhZowh4732lNyNqO099Qaok4Uuoq3h5x
t1P0x3QKJJHHbiZrhZLKeDdv1StReMLRiSx/tTG9B3pLRMPxahp0UvtFLnwPJO6C
3dEHBbINj5fEz8zseSQ4QlBOfaQdZX2KSss0utWv+KwJHlS0ArBCS3iFT40wgspm
CZqQP6mn6v0ozM0PqZx7Po+6yHWmKFnwnVHvkSP+0GsPhYqvgdpfB2nRbeqkjpFx
llwE792UdOWEq+2kuZHlRGO2VVqC2B31YV6FMIPAxKDTI5Qa+hh9V1JcmnSl9dlB
K6OKfYz/JcOX89Fk2GRYDwii/dtZQZhhbNkwPeM1XWq2c+nqjIGQ4SXTBq4yEfBa
sLKOQEuHfW7hn+EYTxhEKr51ScSMvPjXB5YclEMqMmCadQhwnX4TnSdGgj6sX9U9
om6Y9KcVOHLA++jvBexSaQ4GucJlE7Np22pTiQ+e5NGlZ+Owgg7pSmSoSV2sRGWA
49gDGz7BUx7TngCPlTkh0F5rEwbw0zVJst9wHqVh12NniZRvVfkaqQD5L8b2I+80
Dmvu5HoC4kpNL24/mgsDJ+lbXYLvAQu0S3buh+tzzQwmRsS3EbmlSaUfyO2EBHiO
CH384KXcCAFmFBB70kR9EQZShUhN9jbHJBkobyrDrrMRE17i36AKYvMudcLOFSsz
YbmmUeGknEI3hsFuihVWeoYgFUPhBpNagCb0gCAIqFEY9/yew9pQbxloJH8s33t2
yTLCOsgO+nizOMH9BXRmBbXL0sLR2fKzg8oNA1X93xwixZTPWsjsepv+ozF99J90
kKPRwtaKiTLTtU244tB614jD++iUuTS3Pv+qsnph67Sek/m1Uw1K5lGRh2ysV4Ks
l7xIeEt32uNvD8j39q+NgOAuESIamQvsurlY6I+ELKjlEfIEehp9tGA8O2f0N/sv
/M0rc7yhAxuH43YxUe9KLzmXusDsOy8mAXmEBQeblLwi9pIHFihBGzABW8cBZMi1
J7TXE6A7cqJ48RcNdlec/eYkkYoCKWGLPtPWfl9UEhcju9bW3s5swapLOkhaFgqM
P0TG0156yipVoXNgQ9M4FRos4opnAo3JP65EvNIINsshp2hzvPPLdUjrGxmPQhNz
gOaxtx1z3VZ+1XfTx/cyaMzLI/pyvK0rdwLPd2flD8PriQGKB+x0NhifSCJ0iWON
tlvLp/SFb2tQ6N/bvGTshxbgYqos103QpxbyzUMBU3HI1qZZ8TPIr0i10IYj8IwY
naWlu7ZctxDTR+ZhpXD24OJ850cX12fOlRAK3V6fXS1h4IbtguNGMKAbUe0ku883
fQQnlT3R2HVTrQZiLPTfYyz5+gDVZQhX/du4dztv3mtUhq13RcyGIK1WmEUq2Wz9
L383m1R4Ci0WZ+2ONc5kVWER5hkHo9f46tG7eBn8dxriaIFopENpfogzYPz4r/Tn
q1JKzm4qpACz99DTD3tAnS0BtuX79W8KGXBVaoisv/b9qI8LTm2OZVt2vTLvq2si
9D9HBpq6hInm6GVw2pXSRZglXufi9RfrZSB2yIetOPiX+vT8vTvrjk2IYXaX42Ds
D8+RZM5odHqRYyeR0t26rqB3RWKAl280fjivnb23ID28xlSXI65BAdYoNONz5oVb
eUzAKmeoPurlzAVnn54CnX3eio4I/3D4w87BCkqm1sJ8eJFc4S+6wrYj4uX2YGY/
HmiM4R+ONjMhM5mEPeEf415Al3IRpfCz3XR8T9Hue44RfMf/VOStElk1geZZ/ioD
LQDHfRuXUN596zoKBSUF4gvX2+gBfJE+wxT95D39aQLeOe7EAOikfhen5Z/pCPH8
fFSUnJNoHNFL9j4dNb4Sc1WF84dUIN/QX7fXsPIkqjFH8Ht5cK6jYmtUIF94Gb/G
TmzHgGv/jr0lnMKZKF+mKbywpvJUi0E+l2ats3WAX5QQ3dopXD+15+wkG8tHOlXr
dmaxWn6LIw2/hEx8g3+j2SMYTAiFvfPZ/ZwKEseSkLw8FZl3xidC9FV31wAd7vuK
Lvvj+/zo44MNHOgCV7IEGks1Nrntb4mc3gKtLO/7a2tyJ9ZB1h9W1jqHt+Genc2X
t65hjPbOEfQf9fEltaOxVcdyFBM4OM8LLo3Z5S983t+tGA/htu+z8HwFs9S6ANGS
0c4kxoP0AEhr4laY5idY7c3jlJwp34qe/aKmcT0guQZS4sPLOMxUnLZxPKOkuhMl
Feh4+XpyB5Zo2Lomx4QfMTX0Kk1xO9ZqwLP4EgWmop/SmhF6uursul/Nd9m6b7hL
OJB0RycQ4eFAn8T7eGkVh5DQo36snd35YKq5ZHRDk0Za/+oDJRekDNdtFvHJPp7P
ETErRtgJI706DT9JTtIc3QZTYA/32QmckXpjNxvsxJidRvTMm/PLzM6vOFXB1GbM
cVMJmHpVrYC7/x37DcKUA2PAZDchIyNIgr2ZmHFO747U//3cbdJQp5K0/epVS+vu
lapIRLU4NnC6cAhdCXF73NVye4c1xDwt9V3/lMpAtM1rthIK5ktqZBa6d77pcxj9
t1aRQB5BBjER6CVfOAqkIm/U5W6Wu4fSfx3SFk8jFiBJHTWeaOmC9WlzuHs/AMt9
1n65hhvQbognTOEW4k61w/i7earK+pe56ERbNtTlPX23TV9aOp17VK9rDUiVdb8l
q+AktDeSQ0dISDjhDB7f6slCBNFYs2KR0hu8sAGfyn+0sw9r0UTRk2rcarxT6ejl
RmoXmTODmnE/ntdX3kFVM2jjad0QtvTo0M7Rd0F1EQb/e9Ot50kBD5i56CP23fzE
QHmVAg+WBCKWlu+q9fGegLiIKN1Q+0RR+u4xeEDA1OdFX0J94igymnfAmAaZLzgV
DC57uBiFLewdJpIVKjEUeq5DHOpVWVHPG1DNn6aVpFM5oltsUGszJsrThVjfKYau
fB5TU7RhG72F4CNd4oujOONJZUSTb0w/paFXE6cVZvZN7mszLcAoXWQruMR5CysF
sZwYQx+4cV91Sxggj/7pZKFJZQwEWaTFT0Ljt1OjIio2qFHEhcpzQ9NeOmvnlVEk
Asz9R3v+X0hYjeLsU5eOorMhQ8u5V4laYcbslef3gKE4AN5GjHGiI8QFx8Q6wToj
CItCK5FsyS3O8SvGx4xQ2D6Ij9yG+KpqDiJL7XT5BA90YkgXoe4LoLsiAhm/0obP
ZEfVeeKJzxxfhyjZ02DejBCZUNadTH9misZ4rcN2hHtpWtSpmxVda9oZ7dvsgsow
U/uKWP5PICiIzUL0vWWjJfO9adEZhHddq4W6+dbWaJGsK1fX6G1y6Rcx0uf0vHcn
S7kJVN7z0+0K7aUycWeoVMcVjYHpDihBVhtyDqgh5U7/9od23CkatZ/NKWvGAxqM
TRaRKzsVq4fmoejOQMpHr4tmjnEefW717TPGDdNJ5GVDQK7soJnu2OuIK1lKfY7f
hwFJlCh4IC7PjzRTHS0sFdtXgahtnuCvdsSrhZAOBZVW4jc+jMwTDxPgbRmEK7hY
dVriDSZwFOIipmlWD6xRTnJ3OUuZaWxmwEZRcfIB6R07v8huz7qB8SCgFMsYB0nw
NXUCDlO+B4R0DpUx/ZZUgdf26rcIdb23iGqydBpSTUXd2c7zVwWIYcynPg5dt2Oo
+l5yCOYJQzqF1dEtPr+MzRq08kSAm7k7BnupEPwpwHrhRyF6hE6gtkD3+WaVKRX4
I54py0+tkU0sYWz+JGd9NZd+k4jf5Th8meqc4ghwLYmjvQYTVfE1kwo8Vvt+dCjF
wZAFUsquRVJl+KAg1SPvA+oKCKtP/9zhdCXRyHl1b9jWUpyglC5SmYukgCI+RRms
yN49tlp4oxat8CvIcmgQ9fMDMGA0bl6PrR3rJWB9YlJKZzrLiG9cO77pMubsNatt
L14T/EEmNA1t3Zknk+iCyu7HktQAi0oZurZ6pR+dNTR2lGLq4NXAL1dqF0/jPEX0
Yli1xqavQ1+izfUMbHH4EYZrw8e8HZ0TxK2mZGrAwqAK5pqp+dZCzTRn0M3jMFJc
7zOvDY4Gqx5CRDTUXsFIxj6Xpx5rbMebkmUbNxvPneDH9hMuDa15q/4lsuQyYZyW
G6YOec9SjAra8eZlh+BkLmAI5koNC215aeOh+s/MKrCo2DDWovqX8t/eoGSrRqWZ
6qHq/nuD6peqqFfoVHWyZDE5ZRUceHYM5m9V5J772AeOYFXB3rQk6JBJgrAPkxlW
SXs5e/gUCoeGkKVc0U1Imt4saEym38ndb2uic0OolvGS0qNz3K5umu75hZzoebg/
38yf6znLrIq6ql5TSLkbEJP4IN83fi+QkM3RK0oYY+Bne49mY9tWuj09KO0/lh+O
j8sz3Qg1J5NJIpsyiwTkLPsO5/2r1/JP3coMCGUzMOwBNDjEYYh8B4vWmwKnivTI
Ia9jXDt9Tk9QFWSJiBz3j5CLpmBm3AQBbWFMEYTOTUVkZNUZQgoTJLKN5lF3rKAX
MUVltLH1J6SZJfck8cbW9xerU5kc1kpPbFjh5rtuBc8WvAMIji5/aZI7OLbq/zAu
t7BMqBejUqc/w5sBva6xMvV04lgmUg+hX2SlgjAI++s6adEg3jnEqdef/xgFQDzt
XGEWU2CcgTHXpw0c5krmKu5EAMWBlVeDyqYdHilpOTLdONcX6/vQUaKq5HB3wUb9
ZzdLfx05uuDOah3QM2iTjGYZ0le+sXvYpZykIgmxigN/aYGT+kh6aPn+i1IQ3VAD
DHvy33XoyParUxeFL4RTGuslZK65BZlY2NDqMHPa/RYkPMd+dhDO3wFtgmne9Ql9
6A+A9tpD2/itya33q1fQWyPmbKngrMpTfTdC0RlF8JMDcD/zPizVUp5y1bMaDl/3
dWXei6/ekhDT6TjR5KEMprBYwlaqnQICgeNVqQOb7+t8tRofQDsTz1W/OUIimFb/
UT+0SrNDYOhkAMjPV4n2KqiN9zjqYBmXlanZodUarviScmpCu9NbaKkw90AxmmZE
GAf2L0wqXgfsS0DQm1ry7EafKuAYkzp1iVLV9tM2YBWS0cK4WBSeZQt/IJjv6kgE
fKfCzjtZLixJlNgRutXd4pAU9+GpAttKs9EjIePdqqKD17jRpIDnFm2V9Xu4uM0j
MbKPg7yh8w2kQg35fuYNNOTKT1vU9Kp49Dje3VUm+TVf6VuTnPgnHSdlvHNm6mgU
/9YZW+EqWCrQguRE641eWGzkbhDKEboPS6Vuoza7nYsgcK/cs70SLl2IuRLQYP7Z
o9QxQ5Wq9bGmHAgozL+I/D0SSZbyXEw0Sczq/225b1enXJVjFRyUdXR0qFx2C+jj
GYrTUjGddJOvfrPBgu6rilJSfhrJOnOQ9/zURhIOpKTYkpe66DJiD5tJXoONF2UR
Jm9giRdhl9+ntFXESjC6Y8ilLuehOKGoA/7drkIxW8pEXqNDuS+ZDS/NwsHcSQTa
396sFwnG0JNScZNAhmpQmkA4J05QNHZpX2Uza16dTZB0YIZsvcL8aiDEE1cdR0Dd
1igcHufooxBUsTtLcScP2WyZftqjQfB+Eh+1yyfnyVM/7/NUz2MagIqydYwDY49M
VL5/X26ioEFLyUjNSLv5yBpXKUY6VoK/a7GizaKz8jH/vhTXoFacMhyIHXW2+Bg4
8akbWpQqvrfa+XfMyMMLe86fJD/zlltRyVObx64KKhE/lgH7lE0PsZ+1zBIT4NcQ
lGM8PDjxC9S69hRoI056zmLK+NrcqRQj3H2qkwdL5z6Hljfi0EOgsDrwPHOItEcq
c3Samr2X+1/UHszip8nnmWONeir/Tx2LwOMdfpgOaMuL0wlcVm1PJ4jmz1+8XqV9
iimN0tafWETE5HkBBdY495LkYFmTxeqeWl9t9rrS6frXvR/cBweoVh9wNOl/b5Ei
8IflaYszCt5q/vDoPPjd7fORMlA02mc54Ici/OJAGVrKKqkpP9gniDaZJizjT0K6
uGDak8mwradIMQnni/r9PRxhAeNqwHG4xsd8sxYGzH0jyPl7068Yp/cLU5f0FSoh
DKVKGa8oY5vUtnLZj/9Arelhl0W4Um0Thhq7IVo4djTXdgwjpESQ/AHVO3ATt+5f
72RiOHywYJifmfKSh5jx7VGR/UcyRcM7jNfSyT3dtOhF/2+IZRZF7cklRlvhHd07
VpG2rPUlyTSEmhw1sTqO3BU2Dhw1SIDjzfzOMKsBkJouZxTEOGla9yYV6BeY8jbX
JgLT98huDgkCP8gQF9k67sC85vXODt8puAQV1jFZUuSoRKG5chYt0dLiol1xSOOb
0xqcpeDWHtGWpxgshiMBQEJ99cQUyKb/XKeXu3vYl1Loc+HrYEB+mQSyouNSO4++
H6NAfL7G1oRANaecAtJfHf2cbSw/5H89FPOhwlhSnk3slx1w/B/YZAtckmRiywuL
osUb28YOWziRQPnT+kLHCwOhoxAdAhsGt6EpYcVl/WYSuKzWvEFZkeorHrc8HndS
EgNVT3vI+kHuCXleY/rh/C1nK0JKT5Pj9Bsq6iVZPg+uItmuk2RFvlsFY/ARAAW/
eGpbWWnoP1EA7ZgqZGK1eH3lJsbYxsJTfT130xzpLYorAdqAiiKF2Jl0imP2c3Ku
50ifqT/OvfMssgZeOUnVBxfusc7aTzVdxiaQcVyP+4xgrtscNG8A/L4YJkgKK0/h
eb2siFbliwQdq4Nfj/DpbLoXrdfAwsybMNgl7l72CW/+KssQFevbaRm8CvDGoRZT
kOvqnCKtVvP2oFCGzRMqVXqPDc/gmmXdkPAzyb/XJI5Hr0rHje41nAWFRwPolg2S
EjIX2Og0dGM75AMvsN2kCB8Js2fTP+4+qQcu4T/shgLuhSOzPGa/DuuTNNwObKlJ
eRKaSi3JeeunYut3+EmbyffecPtgwtbQ3yHuaM7KUWFa0RP9zwFkLSMoXvdlbz93
79UwcDkqIZl22Idx8FvnedrTJIVuorhC0UwTqb9MNUQCAz0bkEEg88jZ/eglseue
mZP4KG4k1zmCnak/QnmCvhKSBSmit9VSB4ys2gF5q9JTro7ZNpNY0HrtKQO4t5o9
XP3uxElem1WUdwV47guLqf4coYWmjdvo0p8aCq89WdPZ0zKKn/oM7TWbQb1Q55HL
gvWloQ70ON0lLoInlf1ELtx4BTb1K9LFmN8AWQ5XonnZchIib1q1M7kPWaDR7OuN
BR6x4g7A4WB3xMwajDorH+PWqhCLCAPYcKuheN9W8f7IeQlEPJSXAwp2Ay3lmdcE
exSORCGOBoxCC44poDsKobCq7dgEfv3uVrfDyxU47lVofy3SSibacAEmUDaSR3kq
4MQbZYAbVVCqYo4WffodiiAxGcYsj/93yikeIK/VJgBVIbD4joZwHXYiRQ/yLuPf
vifaQuR6yMESYA4W1ll7EJFYJJiYbqV8OWzHm1Yb2uR/f1HjDtLP27khVWRjsO/0
j1k2q9EH/YKxyf6p6J+Ga/8SAc856lUqHOBt0m2Lqulnj3Oykp81hgg0aq/qlIaQ
wwLGEKJvYxhSnGOMqykzIhPrVS9AyCL7kL11eI8JvGMC1z0nTbbNUfVMsYmirvkq
k/1S1x5RDcpuuIqc5oIouT1n0bHso0Lx1vMCEo37OVAG7pEMkLKoS6r7sloTFB4z
YWREYoqGou19MC6anDsJk172b6ES+WgQlmqe3l0kgdqJV7Notv2uKuoeOKPVx/ov
gCENHAbXOTDey52Z0ILAomEuRme9zeYG2uDfcXGiqXApjxitmP128tV5/eEvAOYZ
gkVUlJMfMwoFGnto5Htn4DhyqV6Z0yuHfXxJ3FaosbBxBLz8yXq94KEkmqCbC0vh
SqDSwwNk6ZO0JiJww+usodcpFr2IGgEBGUUaZQ+nHEelQE6tJnizesrxp8fnVd1a
lUmEFLnt9WTbA+I6G9LOeCduSkXu0a/hCokxU8/1CkHHBt0YSXtgUgvZdMjmLD4v
rfe8R4bey1Yu/zubylhYc5ZOG6Wa5E0v72C4MQ1aEJ/JNJm7pVWni0KDyyJ+eQRt
EnvUr5Ti0SJfNMR3kM2eVwckxmlynPOgw7yDoXOPvMK1oVwjvlj42VADuSo8pcNy
J2HKmc225Gsvs95WWp39JMCAdy3zGEz2Eq6XPziRPrEIhBRorkRpHLj15ZihmEU/
larXWbRLbnERQGPkFEldITHYjwsxxKdZQ+fvKMv6sv9NWdMbtd249sHEydbBmuLe
KlPCwwKdtN4h72RIEzopc9Pv9epyOl4SmsHtCk0GLaj1WWFXWVE228oJfEHfP//k
RirXO78TX/X5/Y/ef5kDstNGVlgpM75GOhUEy1uIECbRErm8N9jOKGDRg1HNqD83
xTwAqSRBkWLixMMdHlziodmAaHy0cSQ3A2TZ1zzmpzNszQwfWNKzbj38c91jVZc+
d9NHfw7jy5089qiFNk15KM16NFk1fd/Si/Qn0jE2K6Nojv9Affe/267U94dQVHkS
FIJ37MqEA7NqRdEnWdz+KS4GfZxu6EwFmJ8cdisXoSHwNglGsu/xX2tIPH5M8TtG
3pA4ioo5hdU271y+0v051HYdwO+XXfcxXfRMEPlq/OJfTkpv4aYH9kOsJvC9j0rs
xh4ZZl7hWh4xX3gDuB5r2C2mM8wf2yXb4chl8TA83BvEniOoXi9yfJ+EXrLaK7mY
99kmG/OcR/P2PSGsbMtdU6oKYJTs2gNlIltjOH3v+u80DYtC2PPb+s8S36ncnj82
aMXu52s+TQl0ECYbbHwLv5E396ZYPJnijU/Q8pYlPhtnpMM5OqXMkbuVAh0PuyqT
kMWQ845gGzajorM1fVs+3wQSEYIKVa/HD8kAdreZtbfpt3RkdxcF8Esl7tzLBXJc
ruF+xk4esnEnnRUN/JcHKaZz9PUc0dD/efx/XEgTRjnRlBUJd9bSqdtCyKRlzNPL
a8dbV2WobVDW2YJ/pQw9n0poShmOhFW5moAsqw1XxkTfWtBHrcUYA1njaof9kSlJ
obO+rUmXFJQUkoe5iWaKnFnocMjSAYh4e56/z1zs5a83zXDujnAMcvNoMpWr4YAN
dldn/Z1mqp6IiviZ6+jGdqfFrSm+y3d04iD2azzl7pYZ1Uu85PvLwwFR9/qkoK4R
6LHPCzj6+ICHkoItMTX4yEM4Hhwvw/PNfuaD6l8CuonA6GfAviSu3l8l2gJl7CgG
hWgWcCJuUOaAiipEfgwFWzsMYbKufTkBRiUWP9hJe4GEH2FGqs+T7arzkIcsbpb+
7bNcPIV7l+pp0jLjc/dMDQbEJrHje3Osxijqv/wAOPwnPlr0TiQ+nE4spR8I+RwM
Sz55BIoon4AcumVWX1JcM6eD9fZ3z0fcStj3lWOhpeo6X+b+EJmsHN+1BaVvgjw5
MN3rVwvoR2GYJ79gOJP90U2gcOHVtG6N8stonxshCY6pN40NvoDDIcvjtI1NUTCM
+iG5vq8BSsFsLmTt8Ysvm6VmJIWaMNrk6q2Z9DGwW/mLnCyPhFvcmqNNS6/k3lC/
W538O0cau8bp5uRGXVQIjSv+ZnT9TsFcn5ltSCz8QO+7x7eVr7aOZDur9VPMBCJr
0Ro6pJE4vVPenrPx3NJ1cQsUaK4nuSkPBlhHVGm5kP9S7T1PuuBmyN71OtC0HuDe
cfDdF0odRL6aO469OqAo29i9RhwpuN6tFZy6QWLnqBuznezQezfotP0OZMcLjMNa
DNrPM+FkwKeIBVEKyG9EkUHDmbfjNAPEM+CfyNbs/1h6dNMkI+8Zpx7OBuZlwBY4
FicAlt8B0Iv+8p267/y96US7hpevDh9AAwRznzBE0MU0W6ABQYSCQG3UaaVkkZNQ
SHKSASy6WaRyec9uSoBFXKxLjwIBxJg6TDGwkDjdadN0yzppxWw5dk2jgaAwY03t
wN1RHvGnedszTbMfZWWJng/FUePxxJqXf5fYL9SoMHLEl7GeMWiV1ElKrkgS4gSt
R27bawqJQZd78IYIdZliAhlQG5CZBzpNJVhHd0DZyyM6BgXf4uYR1QADClcGDg2G
C26ByhaY4sMBVJmdSZJqyIZNTwZdeZMgYYHnTp1q/tgzzMZqlyHPHAQTwnYjY7Jo
uBGXfQytutGvrkUXIuupQcxJFYx34Om2poGTWiC4SjZt6LBCUxdC4ScPhZFmKygm
LlxLO/46JL3tUjUiskHxe9KkwJpyu7+gWYObvhHa/k0p6HMO4ZRXPyWeMj9snd/t
bC/WHZPf5Ysp4gXtxvR22z7/B/WUemr4+OHIk0oOjLjkBGtZXXvXXoupcjlmO1Gb
SknJmtYYxofYRu4HDP6NnLMD8K3NsOgnp3KQAbt696VOUXXNSg8C8r8QnuZO5ZMo
SqjBX/s2Ucs2P6z0GLug5vvbE/+te+LYnGIFrYotymHMKfREl1fSi++f7xGTpX9Z
9bxrQm3LN1VHAurTjfL6CnwsjpyRLF3B4bJdX64ASd9ivp7b+18sza0SOtXrq1Rc
Ypua2pPDS6oddR95+t5tny50CWfiUIvsIePdvsmiypbpNnMBQ0QZHZw+4FMh/WuF
WjUBLDTTWYu+Pq1UslVROOld1rQvlxYqX6UbLFHma0Rui2DtILPcTuQA120YOll4
ogH9wtJ8daPwZLZAI3fFu2lUMA5HzEebIUq4bN9W9srGSxMJ80ko5APg0LFWjemA
SU2XStSWdTn6GaPQPPgrFftIegXF2W4v6riYpJVS/m10SVIQqb3nRdZ1kLU7vs80
0G3B84288103xhmjwgook7V2pqt2dTcuqCHYvJl2AcqoP5oSc9W7FSSMOKhCDwPS
tPs1/PIvJ239nBIxrGNdzjd0Ze+4P3juqTcqcU0H/DvXo8qecF1aELQ4UQPcag8G
VWC5PbezzkBPjJJvbitjGgOO2totQRBplTAh23mPJY45h/jCiBO8WnNMixedVw64
9/vqMLiq+PdQqwyjoIA7OE4pSv9KI8Cq6g2vqRKr0Z9P/rdgrZehpXVH5BYubMyq
E7N1rRR6FbI1XMkvZ1piDyBvKSR5ZbRo0IpZf5HgggqMSX9lh7L9wi1lcOr5PXqT
L+44Op5mGIIpVP0ngf0u+mMu74C7EXgBC0RGjeuzohsqsjrF7heGHlNncdfHCSGv
IsVPsYiq3RdqWby062RK8cDtRqhOCaBX3JtF9yCaih4K9cWLyog4xPYfiYuVIga9
K0X1q8XUv2OGiDuobKykfwZ4Ud/Wx3lba4tlI11e4czWJ5ARt3oHyxqZV1sDhRWZ
SxOJ8SoSslzBAoEtzCrVL/AFQZfrSRPKzuQ7urUuP61qaMwtYYa3X9821b/Go4m/
Lr1Pyh++VqxEUxKuxBC9TkqeIVkvbYNoglk5IVyjZmCUoXR5669NNpets4TA1flo
2Fb+v3qyJYbc0nps88IE0MRBU713R77rsDOD8ePg6a+FwNCXbZYvy2vocgC67jt1
EV1SiaGNtO0xa3lHR2nY439S4CxIPLFmyjQh+Lg0uHCSdvbDSXw9x58z+m+1LoDR
BNxIyUUQvWTp48m2jptQ3VA/fJyUJfK8grM4eiRQk8NjBNShxbM7t6w/p9ILiPRb
FYz/E3q/xy2wJ02spBgZEFF62B+9TERCJwapoAPYKsT4pm5wbSdt5tqESs0FWIxt
5nSsVjAjcYA3tvY1llMHIL2sKbRkAR384kmD4cK4ee2Msc29/YHi4lBJW/s9iZ+w
+Ja0NQGgdgRRhJ27+x8rLLf/6YuleX9WkbUB9gUXXJLCHXAiHEo6+UxBN2bSJ9VQ
JW4G3DYxBvmdVoXvmcytUYjPKu3uR//spRE/xTlfGthtC3gEWSeKBlTg8f+7Jurx
S3kz8G4Qm9AWwb1me5GjhB5Tu3YU9X64Ge/eAly8fjElEQRNe8xRorJw3l3iuOGb
lJ/aTZvPOu4Ev8ouTkU/SzIrVgXi2+JcozNqFpEwuV9LTcJwxcGl8zJqYztRGbfd
IdVyIwDhjCsdpEE59Z+tsYZPLWbfPfzwsor8r3L3HfM4yJ6duvN2ROwUIY0Jwn1V
zDhTImKi2KNdY09MRtTgPN1+RxM/xLie0y+iL+cWp+ZfVYOQkDKmmSScYnc06wVQ
V1MgfZWT+Jw3Q6cbRLUGQSHrk508EQkwBCe1yZ8h19S2P+4MvZYZ+HMST6cZ/vgs
mCmwnTzVAYTIjJW4qV3fyA9Zd0CmZ0zVQ9b26+kBaECe3XGeZQVTwsOeNerdx7lx
zlnjlGMl0cJNn1Va24Ikg+L+9NeyVf+aFoDF+NGHbtufII0FmMacIjlszpywyjzx
9wfkOWevsP7qC3RFNocd+tKXM+h5QZiya8rbE6war6YaEH/1lCl9gUipoASI/tFf
yJvdb6ETRrendiuW+heoUHUYt594qT2L37JxsG/M5iT53AHNeg23XVNNwP52/ak3
25WfvfnapXNVazjf8tN1BYrnNrWHBWjf7jYMzvncrlmGGma8A/VsGLUAqa1Qi3LT
6UCzex4cfS0Vdlxf7EwIzsG2DVSq08PJtlsaqyUBpqkC7HubmZV1gvTfHWimIvJl
q5woWC9ADfYwp5aMUK278KgoIbuqzp95O+twP+y0944Rqu38nidSz3UQQDQjADYb
H2G/emR5xCv8WnyYuWN7XgAJSkFdfZLJiOBRoQ7sW1ClkSswmsYptKrt1PpXASg0
jw7nQphuCwTP+q7/S+jdXGYZvUWEiM24TAXvF8HSaBQOTQ8lPOSIk3iNTl50kISn
5gGxwVMwZYEsAHrnAN2PxZLyIEGX+4PpOtLlNdh7uwNI13Z7ENPdVs8JtQ8QmRbz
CTR1I9VEmm5Nm+aC+mcnuOnt2+OkB0BTVy8yCWejuh1D/UvrYUlcM1yfp62M0g0r
Ab+x1gzzGJVoF8gcZZiTzTe3XYzfmUkDcsVi3ksqRoMhhIFQIv0/uLx4vfFQljZS
o4cnspm5xKGlXiLXLm6armIoYMN+jNHgqS1z3aqtO/Lts3Fm2qO3zfdIbVTcvicB
9tUjMrMUMUBLuq+4CpujBn5XJuPkkatTyBMzNXah/19S0g+CsX3B+wJ9lK/vqMff
siGvb5ehwvNW2H7KIwxUo1di/ZX0sBK1zSF8ROcj5WYCMRJQlU98bSo4ak6V9Pe+
z5g3Rx4biPFbNZn5TbsuJeD1cMDfb8l/uTa58zOm7yC/Sr50aurDeYUtZrvAVcoC
eXojmqNwvPSPLl6R4iHSuVzv+idNNvGWSJ5Je4jOGvcyQQqGB5e0EVMk4BC+p6Z5
RvK8wKkvS+GIVmECq3Ol/8sHEe1xEC5I5T3VqJnjUYct5tzkqTaek3pfHEphXCO3
320IxCExU//RVRAiMk406fFF5D9va8s/FYw9SHSkQGc7uf2sWzv4dz8FkM7HC/Ko
dgPS7564cqJ/uyuYfuYF2x741lSGTa+VRlf2qJO2cbJS01p4R1F8OVIXdnhxCEgT
hfwUlTUwbo2Z8kK77P/GjKRvGYTLszjGXsYfY+QB2MosxOCtYGUPb4EqGuzH3KWJ
3DrlDhqDKT30S37C5Yr2JbRvVPYReXvkZ/5FuwSFgI7UXwXYVe/yKBFjPP/TWxPr
dkfw7r+8kEL8Hjc9kXI8XXjJKHOR/BCynE1aOfz3DYP1t3Y6TtVJzw0NlqJeAoAD
jGHBFdkjD4Y1IUyD864yzglaVrP1cgsaTLJMLy4KCrpj6mSD9fasNuLBQbYm7iLV
C1ogsASCYbyPZBlXzQ6joJ2co35Smzq3WiX2ipv6ppchj+HJ5WtxVqBFdjqJnCF1
N8Ss0Wjs0Q1ExkduxCQdBD1ffuGRwAEoZ6AxjEE1oK1GSinYbFjOCMMHtM4XbvUd
gyOa+LrTyNFgYuIKLnbuYJu73RpoeMuhI4iDYPwkojK1h1HMqdrFYjzxQkxkkxkJ
fsriqsa3uVQvH59sxRGqCZihNjUzga63bnT/V8SRglNRhvDFKWjtxqzkyOZvUawx
Cg86ms4dHjjadm1j7hgz5TkzmzmknKjaA3quHTxyMkdFCk97ko9h8VrIA3j2p6J3
GHcUIbVEVfnXx/Nt9Cbyf92Lw/7J2fIVG0nANL11pTwIczRo0eT02eSrXNaQrAse
EgKDjo92rwVrFltLiG99g7oycjKPmCIkpulvhxnrM/wgHmHGzkBoopnHf4pHrgmt
2q4CvU+5wp3C45D3YCqB8QmpUTNjc3tG2+Ugo4INn7Ns5cQxOiHy8P34dzJzZMJU
++i8A4TB9G75SAyM9gvt13jIxNEEO/Yu2/YZVbLqkWVoRJrY2mPbBN4TKHE2jyk/
jZozkMf6mHhRCSkQNcwZttIhHHXsxgku8MqZNXcXEMV5Mqvb+64DZVOPjulBn+tn
7YVE9et24/ojy3HJc+dV2Cq8QsiHxCdAn08BnAF/227jxanfB1hEZEIeuSLgFtJ7
HTC5FDFYoADSHUvYkDj+EV5D4r4RpoCGVrj3XgZpL/4qgJW7QHKdt/wJYNvkzmJA
rc4dbuxoSbOdgq8dZgMA335Z3mo80n+aJcu3TOnojqy8YakMRKliW/aog7DF055H
67ZdD4kFzltrHgNf8j0C9wXRrzt1A9takGm5kFr98i0UmRknVIG7I4WEWkpQDZs4
b/eyIFfH9Iv+dzBLLNlPg8AiukNwxbScETJviWZVoaZe41KUYSwrH/d1JCcL1yIX
lvIuqdPQzxeCpMC6sODwVLuqaDQhS4IjP5t/yPgzUZ5LJ20gu6bCxcyYI0nJjSIY
YHW0HtTAuJKW0z0+3Aa+w37M8ybXVs19J1RniASOyKo6s9yP8fmngHUUxCqEyydc
uydRvs7PbhLVVCDH6BL3gzibuvAwqhQhaMBNqso+xgc4JyzMY8ylyRRKwJRIxhfH
sU4uXDBrfBmRs7UD2xsUm8MwmceOgXLxnVCtbnFbBTPRxDL6Z1ZRZMYZmqS+ME38
rTgZxa9OhvFkSJ9QA8CmWvlOdwAK86ijmoAbvDRL2f63jGPlTWQ6qia+IRu7UrVY
nXDrbr3p9RoKjHaGsW3B8oEbUgZq5FwsqfEPrw9Wz6xo5cMbOvErPdJ8xx3UIN1H
Ob0bJq5IRWEEubeXpZLNiOZc0xauvNyNwLQzg3iRxrDfKCN5Z4sqbXaztxQPjZE7
Md3Jw+Tb4Q8OzdtedWqNYbX1KYw3o6CSQRlOVui8mTeqrWQ14kdr9j/wCL5GINps
NfHCRWkuYXqkeh5ZEGrEdHVD8OqFmNSguQwHJ86zCDaY4dfxYZbGa/O3ODKltvPV
Vbcc2MMbM+fZ9B8+ii5R8XNNqFKYNuQGF79kOxS9Snzcxw4VfKpp77+hagihtqLy
29T7JZveJpuUEgKoR2e10JnrH+ZhBCfpVWMPvta2Z7s7WTCg+t9b+krZiyvtGCly
r898XXWvt98qOA1WchlI2wPHTn+WhqKS2v8eOt7jKLHZ8pBt/P5M6280C2rcTOd1
uJQWnCCUXQ8KkAaZyvzK8gc5eGGqtFvxqSYxrF8rPPsIX4SxtMgUC67M5cCDlPDl
LgHwxtNTgdMcBQDRGaTauyfhXsLP33Utg7tXFuSU4X0XcoWEURxb8IlkJodVsyTq
rAade46vMnT18N7sOP2pT9F0Cq87EL5cZPa3DFFQW3Bd3wzo3s6Wwxs0f4P9CfYu
8ezcF6ZjPOCWds2VyolR+ALCuuhcegU9zIEwYm8sVAjvRURBq3qZDLFPA7GIMbu7
7eC6PGJyDsN2pFwW7xobqkqU2E1J1VRwOIX80z404saeKtF7J6zua7mxZinLDtLy
7MMdx4XJsr2F7QAvsyCc7GMOMhbE4e86wK4HV6qjuue2rnbe34tfO1kU8ti3Ha1Q
4ZsTCwOxaBaWMyK2RrDThm97swcbhMlE3c4mPW/teE3nVBnLfU4buSoIberQ9YB0
3lbstbGmVcfQqe8029SX13NPkw9NU0KaIGB6ypzwC9iBPSv9hE+/2oZOdzWFQCOA
+Rmt0f3vcePcX7XYJlXH1QaG+CSja6FW+ebtwE75zgXEN1nUqw1kRpyBdPn/e3eM
VoGV0Ty4KA9ztqh7uVwm6hiQahdquhQuIYe39ma1hF4vKZgs0MgPSJ42z1RjWs/A
6zvFCybVEvdgJgXV024GM/sveTA1f7onqLRmUurw7xzX8tZDrto814dSGcChlkhS
hWavSGQIAk/yFNp6nudk7jdC24CZfWxU12TpaFJd7vbPlJ43eYnFjlHWQkahFUqw
uKIsiMv3lg+BFublc1UtHKT5eox9qoNPMzr/Vbi04/wQOK+1agLVuiBDwbYfCBje
1jPkpkB9KE9UU8qBrXpxzjJybN3Jm34Qw5CbvLy2GAh1V5GiqvXW/ILAdgKJRN6y
JkfwP218yfb5er24163qS8uL80awgseGwH77M0vy4xcuDkpIVmiHJNkftwv3QSw9
3mrNndFC5QB+GHtp20kGABpCFuU0bZxPqnyqEzFk1TmrDAuRvVySX/DbIw9dqxwz
lHcjy3LKB2ASyZBD42UCaQXvJdemW9e/4qj2aogXSg8e5MmCePuavtsCANUcxYVQ
7qA7DROwdDVzDZYv6RkFuqLMO9/oDECJnUlGB9mgU5KtShwsqin0YQ1BpS07zePE
FsrMNMrWvrd1zy3WlDyCbWSrebmqt5fV3AdmZKf0ldpXgt7TnXeSapNQfI0Tg7MT
kNbEZnL2qVJNd/xKw3xhER0rFE2SX/uGA/eSLJvEVVux0bLzEgjOdkW8RyHLpL2l
MmwZuaSUSrfuye/8BPnZv1cGk1Mz3w/MwlL2Hh96ylI3pnzYlzo9xTNjUEvR/EAj
NVu+ipAbMVHvcDOwvWuYTBTOgfVX/9pCOLl5fNI++U9ztgpIZUsWggbmkwPTyhDA
vccSrQ4LxvDS2SHyxRi5votGjM6Mc4v/jja/APKIHWiAw3tPCvdvjQBSCaZ84QkQ
G710zl2vH7Lp8OgGwNWoX+yikDM4cdZix2k2qA7qcr1kY7vTDfdeEaE0EjQfqWHB
nRqL9kWcnymMFnoCcuyzNCjHg3xyMnpzwxt5Cm7bOOaLVZCfIsCXNK80UFmuanpJ
edJke/8j+stB0TPygjce7JXN7OfR2RvqeSES46JIBj5I3VJp+9MGOCX60mEDoRs+
QXyr8k6mFXhjSDPIKAdd9ISjkqQ+RjEQq83q2R1XOSVf0U3EO1DMREXLC96jiOhk
Ug5C06a3C0xD2DQHZtihd/eCmc4GCITvKjlLYFsUQlJQPUT+yNgji50OxvySBa5G
Ua2NSUowYzKY+4itPprGyx/8WGWdBK1mZYAyvDQ7bDT2jj84vUeM4tyJfTbKRr68
TWJeOAjdV7mzl8SPWmBD5ea/HTgjyKNT/VYoK8pRZLDNZ2+tKH+wBZQ25FH1nvAV
lMhDm1KumxfFz7xf9WJtrPOectn6ea4eLyxMmooLr2P3TzkEA0BqV3UWKdbo9caF
b23F66WZxqcJwFHYX3oMJp5K0rRjCi6uOlsSXg9Qsr6kW75AcdFRiLSCpnj4atwb
BkCTtvXum/of3gw38BAOZihhRwFjym/nDVrZkK7L0PRO787yA++rHR1gwh51C65u
h5e0MxGaIC1owgR+ODQ5o3Gcw/sQ5Tp2h3f6AcWRvNlvhanUY6OZcFjUrw6Efa1H
ZTpy4guARlaTeHwOrEZCAGuRSUFp31wzgF9bJQB3cNMQp9F0OJXhN3li485d99Zp
3do8sthcC0roO9CRQdb5Kj/1nlOZYF/oH3XWaoBG/A7BCLnoI5vWIeruNUqou4hR
fx75oEDjA1FCAV7ebsNao84UbRPXCSYXFVp5HjJs/O3KPvGGRpXU6B57rEmkN7t4
9KcvQdCv89sSbXKa8ha+AQCC4b7GlbOmDua6b0GqkCCF3ET8QUd+uPEHyPm/b1gS
9dPG/+6dUY7nkb5uk6W0MCrV6pp/1ZM3xckXucocOs/TolkeD6WkKmnlpssW+oo9
EqcyYzwIpGh6Eg5H4/4oOIB3c91rBrEkvgY0qPQVMRBi49gX98Nj9+jqoYSI9aGt
Uzbrh6TI1UBh+Y3M/vqbVjoB93LP5uiv1T8LgHlfGhRBgX1NuZhnP+pGHZp/5nYG
8bJJrn3yUQ2jDWqWlK6HzADO1HYLaYwXQh+JkRgXkb6lqXP07qM6EYLz1Vwmtqt8
DaPeoqpBHT6qWzStwpeW5mgh5kGqzwrpgfwklrUc7e/hkNIhkNix+LTrHgnNEMIZ
f/G9wMZuAzUC+2ot4uUgjAbK5meIc6jWEkTW+7wbBcuccjGigL6GjmmoPFLK7Hag
w+VKSG2yY0QwARGp4bZu68xCDh36spPaZdy4mjjzpaEiXaeKaYKmhAunQHCnVGAd
CrsnlhNse1Rlazg/ZHuwT45I1nKHh8N9V2ZRlLBb9/WvFTCv40MKS0r43mdb566h
YkmHxIzkjQk4HI1tNCRmjTX1Pjjj1oPH81vAxqH2HfnbPDptc/J5XQWzFDf1TpAJ
TH6MIGdy0zKFR42drDWa+lA83z1a/v4IasinqI17shPAkUcM9uc/IUXfkWXGsZDr
XgWkxgBvup6zZR2v8Kuwd0ExvVlq6O2Tsdiv4NTOupuY/cI7dP8X7GeAxhA2hSOe
qEXjKXQ8vm8Nd0Z8WSLjbgQIBuUhNGUuxzOZR/D2AIV/57MgzEAh5ZBMIapPbTAf
03hL94j9jcUGCNxejvEUGvxVPcMjDJNCm98PVNKYI8ItLy7OAmkLSCY9Cc19Ja/I
Js1hQuOszwfpmD1cqp46tez1byz9jt07b6b1xAFWi+pf/+XCCUfyBVXSo3ChYx7V
DkDv9wwSSKfGeWgzdOTHVI4QtmGbUD6XctcZ0Xuk852rgm3jGJ33oBbuZzcHurDp
O+mLInQo9VxqiDN/VoLWELevDzcpvwpKtgwcvbA7oL7SsqHVMkAuKk5XeLy9TiFe
FwaiNnqxox5FTVwb9vDVoRVJLB7smCu/2PBsSAOaBJcLHbRaL1nGHRW8GLVenOir
Xk4F76sdwp56Ynxh8UZaUTPNsfnVAJkaMYSlaJFc7j/Gq6erwlxpdXm5bIqSZUVf
5+jpygExf8rwEdmbm8lAb/jVwLMBA06eVFcHIhPcpcQ/Xrc6NOKEtYMmFsI7zKFe
TG9YGQEqmzv8FedeOfDCZ1HCy6lX2zSF3LdvxVVQCqhOysaBUajJzedjekzBATdz
Mi08GNZxIUtWmXbhfxIk2xR1I5oeAwqbAzbphAnTNFH0hTtBT131SkyldqgnLuZM
bq5xC5vBHbHM9fedHiyCNrN8ggxsVlKCu2VhVfVuAErXgrnT0S299sfeyR7hgRsM
aivZZA9lzYOi8SI0XuhGUZishjZxttDuOinXrePqFeMp3nRJvXe3KqA2Dy9aO3hI
WtYKEBiGrk++o2dRYP5qH0LDMAcf12p/nSGJVDv3YvgC4exHSd9yN9u20CuDAPOM
oKHjGFdkyaMTi7kI7cujlO2y93d2VyBRuu3rJKzr0nhuG1yl6aRozX7jvx+hqyba
WibYjm2j1+wt8bCzQaZkEUkNJwBtx6wPgVD+mQaQX1h3XHyaOZzh0Hm6eEveNpUE
zEmCvIBlELirkijQ9te0lwDV1O5JeAyTYmQd1H4oxcV9GbBVOUCvGuPfjEmS37QH
LZN4O8XciM0q6WEC7eecHr9FhVGaStn546eain1vHBtuEY5/M+J0c4aP4/kyTEiD
yBFg9ZElIip/x+cv5OTmxgb6U2V6oHaOkGJEhAg5+VKR4+p853+Vdqo/p95cax0o
WAFi9XnXAbwJI36SV4/2qaCM0hSmaLJisWKOqGfsUiawxoudxW9GyaqFrn0aj2DN
r/5XE2JXCcqBJjYc9w6SK/q6Qe3tCU0G5St+mtkedI30Ex8weMJmUioiuqaZqI1M
bfyRFzAPzlcKLQDWMPVknL7fkbHc8GAxKz5L6aQia8d5wi6FdABtMiGVsOkIZp/c
zLuvFFoWV6EI+VPNDoSTk+GR36+HxKYqoCZ6I5WlyYpWHFpZitaUDeSfXZaUskgg
GEmLcp1IxMNbT++/nt9E9bz7Pw5sZ0k842ehtOKFOmF0WwpP4hZfrMMHwpLk4SWH
KgrvSymbuEiVTDw4iTn3p3FVetfDuVnK7gYvW9vVzoRKQcl/Me0crIJEjgSEg0ZJ
FIjzy8kHixMmyvyr5lo8cDynFZPGWHNkNrJRekNyAEHVrRjgSmbcY8m50HY9beoC
d+20DjfqLKW2VTeG42RW+235fBTH7qEgCgIc5Jvugydk+Mnt+3BMFlMevqNp/rAJ
GGRQA1rJIPeGI2W1Snkpda5O73PuISQ8ZmFXGL90MjAnSmnW3O1cPRYHnP3jEYhh
bocQFbDTXDPQbXa/pCsxfPzdWd0VOmeSgGZUY5pr7Wyb608mf3TqDYt3hffRUizg
HNpNGjyNQ1S48ATjDWaVr7YSfxPTe1msLp3hlPj1ABEC7mXrGhCqijUk5X5eCv06
OMSo0lfQX3Tuhwgo2ZTAXlWbYfWDY1hBBLwmMeHWSBUZtOcggnAeOMB6jlzOrK8T
WYm5OgKOnRk+hYuKP53bl0QNWXuTQAY+Mom5qse11qcAB71AUeD6dsA3S8dnAMYo
KUUNCTCQcGfnMA9/mUkExUoUF1rzmWN8FWGTTdTw9QhrlG0I3pqIVTjnrAScn+Vs
/IZP991zu0ic6aNGoLLRwqqu4/3oKzluYPQdKU2sG58rz7n1PL9CVbxBaKDM/prb
Y5Hh3tSYg9dCEGrPSfLtxchNGPEk9HUtoAbhhjy0hR98yRbQNvM1cGW7+KuT1Fvz
LLUYOg6GaFlcgzcsKSzMKHO5kYXOR57bncEchrFpOe05j+ghe9jStLFf/BNoHmeF
x3x0iARVhp2O9O0Q0jFca83Zo0vLmBltcXxG5EChhWVwXA3sMLny5HbSc6e+kVDS
F0/Zxmmnar7ZLRnsrQ1AXhJ6fKTj1FIj+AfHiQRh7FpN11P3vj/bZDFPenuKiYoh
zCUeU9WDYomQCUXuIWirk0ufG6iOGIxrYgDF/LP7tL0DTOlIAr40xiYof7woFZTr
EMD2c1R+Ec4WLoIrVfnu2myKg1Lf9+ZauVIONHL5lsb6aqvlFfejRj9+OQPgiygY
3xm6FIpbFteA8XM35Is4a7W01X0YFe5rwYrSWGDqKB4DaVAQP5U2UwFs0O6b6IfY
6FyF6yGrxtLdIRfVQPHgA3TPSm3V4DsG4xjCbNzAF4NzoWehm4yywWnqlAPKuf28
e4fFffLeZWgZiSUWb+sBOBoWdu47HiUBT74GcrWJu3PhsrLCJfTvSgVTbaCjf30G
vdEcvakT8ik5hr8/eVblseN18K/BfDKb8EBLmcfzUVJSoLscm0pVdP3XnkeqLvK+
uPQv0+Zh3oK89Afy/BqMxH6TEi0FOzEls0Ab53L3NEvAxCXxLP41u+5bFVjbAvUW
mkSJ0f/hbDyDdjhira7LF+lGcweL1MgjjxTYwBrnl8WZbJolgIG3ylFwwpBQLevJ
3FZJ1wbke6NVeNpIkICsM0nlhbsGjCRpf9PHAfHqJASMCieDUIKITWz/ljVwLFHj
827QHAoMDwV51mF9FaBneVzN2Q4veoRB91UBFh95jeiZ44vZSBmOWCPo1t8rxVPE
hMIDoMyvkvJpioKb4+D9R7QMB1+746tjZi+JDNCkjc+z/MSsqo332V5TAJRiim1I
98NKfIPUgFJ39YEuS3x4YLftTWup7TnGE/wBpiv8DeOb7qLSmwtbnH9mB51yq+1B
saxsHG37luemOejKgjT8FP7H3CzLnlAw81vGSZOIJw5Xx7iCLmLObQNSoKd7LjMm
JeOaX+0gVJTB/NviJQII7eHqSkX/3zkgOCC8/uRIVVqqTyxnsxEmq52iVgtBqTi0
TvK7Mho5YYJEQhwSEVNgxR14gyqgz8/j9Yhk41KUI5olDeA2RwTXWVijYE12fdtW
9NyYRwlI3Lb3+sS3aybbUbW2NUCfhazw/8Jhk5UymBXvmoaeOAA5v4E+zBbjY81U
hd2xgcqlk1RndPQekleiUSkiX9Tj86yKWrmBxeFbgHw6ikN67yTUWmJghjrHM/yK
y9J1vTP4C60U4mlkd4GRxW75pnzqgbn81YfxtzQZr0pYg4Nse/04Sei/C9qPIVkt
wH5z/GRS1imc/GeUlH7/RsOzNqjEGKUVsmAAmBvzawtoWOSBGUBraBsrZG81X8ER
ZO3oWD+RvcTbeOVzjjPQYNiaIlRqzrqwmriWyulSwqoN0CdmCxe2sUz3S8O2otaY
k417geXnQ4Awf0DXFGS2IjrtqiJIf+TZu3TK3akth1DKwaD4gf4kDlVhbcl1nsNL
Cnm+YYaHKFmrdawy4oLWsreuq4EI/qK4YJIdDa6DvpQg37KTuuvDbsYGTYQv1RKe
K8WLr51+QQnhrr+xuQ1Df4WWQMP901Q4P/vI11blSGPG5j44vLtMyXtL9caTO/OU
f+qWIuVTtapB0+baqhM0r47oyMhxp8+o3YBMjGbvgqrhADE7xs5vDCxmlTPeh3Tq
+GE62T4wqPLu6qzEAndvynFjbRFcHa3iA0FrE3C+JR/YmdRixxAtpi1NrdTMxp7i
XZAn7jFXIZSTvYYSn8wkUcKbdekRq7Stn7yeCbhRyEG1RI/l/A2gRdEOThH4H6kZ
1ugrcUAQp99xlGQFj5+XkgeniV+KrmWEdNQHjqksi+eH14zqX4rmWXhKLGM+pSYc
JjbDev/C2VMCJJwmaKqIUW6wHswb3FITzxhW7Sdt5VtOMs+Ep3/9eAxnWJWT9G8U
JMNB1YduivEr+j/0QDwkasQFdXfAFsXXchs3NO9ijty6HiyjSov/2mj4Ik1zgO9e
FS3BYstFYKX9J/QFJyxxLREhQc+6M2OvgyM9og2XzYvAKTVD/bgZj86s8gRsyb0B
dinHyTBDaW0Rs0/WG6/L9XV2XhVFsfUNdDAnIvXtI5FqvauEw++ht3klTOGU+OI3
Y6Y/vRhhHhdz4dL4M6gIj7zv8lkyyF/nGuinBxFVN8J9grAGlG3FCiroCn+xWVsW
aKFVtS3dqjrTVAZMsytIkDJlcDInO3dh4eMPGc9BeVF9zy3Wft8EtczossBR63Vj
WNd90uhvmmysQgDrWrYlRTu5q0gArWOz0w+h09QqUMd8cfV6FEb2JKYz/bbZcXWo
k4a7geZw6fuk5xiYrYe6EUYDEjihnrkkyONg4G58FgQWM4I5MgImdS0jrBWZwcG8
U2C17+PYcTJzMjQmeOp1s2pEJ7GVPYq+S18BCzY0vEXTTmVDejPkKhytSS73d22v
eoH045kU8Jvp/c3YTNAK8+CBfJWl6WtvSopHtZjA0ivMe3uSRIdIBbraQHVn6xfH
r75o/gOEKtcLJKSYm0SKZSwZ0cXQw2S0cbaUhUmfxiAIMv5Or3D81y+ER0bIXgM7
etQZO8P3lzCwOe6boNyl+42xq8C2C0qlSei647INi1iwKq2gWvmDMtSdDP7j/4XL
4KRzHR7z8yN1lJvgFiK1xmq+wuew7EfjXSOMqy4jet+Dk0q1GPFsgxpclQSJHTCb
nysZDDw1MlxuS36KwakiJXh9OECY2MeV9DpZtA8Myg/uuInzwAMTEX4l8GrrtFwy
FttsBFqI8GaWJuJrZ3hQx/c3THxMoh6PkSVoJt2F1erXvnlcEDHalLYW7zcAYnWF
H1/fCgXPar6ro7CObN21+r5qcdXNBc2eitVMksKAtSE3BgUwUbmgRqMnCeEWdATW
4fpTYBMEaFhKFdhgfgK6V0475sG5C6ZEmmi91mE2QbbXPKMSpA0BGVrtXa33by4F
hmPImsFCLrndMN16S9CFlZKQ/NWpc8mzv6AWxkXhPPuAMIVi3wPeqqolEH+wViKM
lAlCRtu+/z1mZpevdrGnBVHk1XYha+GqRiTkWjkIsNq54pHG4yQkdBZl+fAjnTHJ
pEUvZzy2Q2Sga6EVmijcsWHY8EJbYc+Yv7TpUr891VEMb0EHoCr62RCGDNJoy+e9
Eymb8EQmTfIRJ1PM06QezGmkNcwktpJ85la4FckB9Wbj078hwZ+0jjUXO7PifcB6
v1FdU0F/4tEbRQFXuCh+TCGIOFrWqiQDYsKrWIR+QI90bvm0kh1L/LENGdNhMkSZ
VVOa25toSl4eCIU6c5NMHMs6IdthnwHYBVsa9U8F1ilBNJ+452OcuIOgkGZ21+St
12kImXwBhpGjsB0Z7DIP2RAIqatDI2FaE/KQOyojePpmOq340x93Hiv2Q+p5Of24
MtGlY0jP3+N/OWU7Z6toXarwOKuFG+JqECRekBFelkCgUZbEdtPlteN85P54G5xJ
garDtVNHZYSAnBgr4NzxPC/wyZfy/FUFvmvALdCFdpsBxSJTyCHbjXz/+lxWBAue
Khdsftt3GBzSWXK1zEsu+6GSx2pTfeHpAK55QktDXxcSZSKmXYZlU0kMPuXoKlBh
laqV6ENTHudAVxSVSYEqkkEXjpURN3vYbXs1Zhz8KAlA2KMMGkqXPP09fg3vOh1Y
Abgv2UMDdmW0LWj4pffOG4NzU33YkyDF7A6BfEBtsrEXKlyzomG2eFpbe2LLub5d
qjJcfI0P2pnOQyIhgVN2H+2HtGEk2WhT5SsqvFP+p+5/UzwjIuqlbmpSauDwd4GC
2zo3dfGeja7QyUQedUcaWm0ITVzHOQMyNXcRUnDRCCcMqQZ71Dppexu7l/kFyRSL
SosPW1ShkTk4L2TYdtUaYA6JXN8Bf0yFLW0ZKnKIH3TUVSZwvglAqHAMm1/L2j7N
ZswMuWbuAnolGZDdbXZzkYaMPelxRYTOaIzn/23JmklUn72a0oP9B6uU+7ANdLc6
RKwPAI8nn9SiKfF7nsKLMDYlbjlJFbA/+rU6YZRMPJwn1R8VLJV5KGAgh7zJtECV
Sz6srjmD4pHGukBg3Zmyl9nqaYj3T4zDk70K5jQ6mWsThxtqQaJd9lNvnfMxgucG
uvUfYWtCvIZlUYwYHTqlZwYaweOp6EpKmuCHHlsBmASm5QenMEPSjI3GmH2qhzwK
dJHK+X5QHU69DWqdfp/Dwfdf47JWLYkStyhjS+shDVa20tVZw+7ieMH/nSUJkTLh
cmPB7PTpqyLOgxClabS/ccC8cyQgd8yR27wGPSW1PAi01VzTaSxieUGBFLR7CIay
bW+fsgt0MBJKBBHyxAoSy/iuwqQlnFxBHk0OShc3P7AEKMBiZsQFcQZld6pxVh0o
R3F/OtfEJ/jA1aZ5xvLImLr9dhH9BD0WcvrS/HyrTaa1FCfZfSjK+mESSxVTEoGi
SqO+NqCWwYUX+c6vXmLLwfKqcpn6jlh/etYEla3F90YqQFwTXoOohXBQO2HY95aX
QjH56Edq5Agqekft5rUAVbkY/xJnzIk9iKm1mDPBa3d2JOdVXA4XKcofk/M/rTdi
YJDvpUu3eYgttnC/Bd7JvZLIS4LpR5chnnFI3xbSVwcEstyOQMJb741GlzzUWFpN
C+j5JWBO5N4PUonJ9/98LeZoWRRl1dLG4KOaCFdcoQeVkGLf+xc0UwE+TLXSphLa
hgblAaOpucVq0t0RcjN9CBn67mL7NgZxctaiWQdhsR3CVIZpg1bNU+8+1G8Nyy+b
A1YChPaD1z5tHJt0vhhJM6MKtHDqCzECAvYm+y94TD1bFYdvVRMOT3nq6rtf1N11
Td5fmCrxCNN5fNqrL8xv1GlCyNzhBAaJeqdysSiADiyv9i5MIZop+lX96bGQCh1L
hv2nYEm7500/AiqgDVbAAdsHhi7b/d/ptZW9cOfFcxwtYJUCmEP/RGIZ4g5EvQXl
wO7tvsir5OHGmA7Wp4cqjTEsKytdEKeY5b01RB5F5dCk52/dBkR09tr6l80aSBkN
BdT1zuc5+SHnG2TU4Io8PZ9+uRhO/VxL5/fAEbVD/FlTsSx9xg4gmterPccq+/gr
iIuPUCglZTMh/gULjc07E6nsP61sAvma4EURw7NvS979IBlbAqVO1VEjr0NMgeBw
qrhsVz7VXl7VElxAcTjYpwUGJ2/lzol0F+6vtMyTxMtwZ/EvNoiw0GTvUlfTX7FN
/rhDAnynnQ5hxzqxTfGrQleHJysmn8RpDUKIlBXRnoKjlJAlc3xwNmDjuytb8KLp
cN8dCc0wq3W8zQ7kkDLZkXDOWmNMoyoMWG6REJXW3QmEWAg3kXfVk438MId+gpQC
V1sOfA5mA1UkQzQwakm2TpZmM6oRaAQgH0vt9LE6JXtXc+5sHm6LrTPMpk8bDY+h
UyfUaG47O0Oeq0oh02tha5ITseOYOYjpV8JSC416WB/7dZry3q4+59RvGE+h21rm
nXiPdiDk6WJd/FNzAp5NWLO9lEfDQBV3PgTs3zxf9LrF8biYYXPxq7Hpuw9G2qzz
ePJ7uJslq3ei4b2u0yYAHODYffVjcPiz6ZwMFDyYhvn/5LKZUDmqIwP49Xj62Bkz
N/Oqv7cX1MayOjxSbCeWZSN1cs8yfMn2ZDZuECDAudxEbe9COz2agFvkrzNXlple
9Rrecavc2lCOMCYmOrCaOn0X19xf/6JrLDRrwWqb4McCTaNPTsX/+lXqMpd7fG5t
HLABdFhHQIsBgDiasCyTvEDLp1myjE7f5YuiLSOdTProFMeNvbQ7qHURJ1sSVu72
jixm4C5kaZICEdLW8kctBB3JHJaGXa382aweR4sKd4XgAjNN4LIfgEhCfnzwh2+R
Id3vaxNJ2bp8xOjwxlYQkzIvzXp3Tr4203iWQZAVki6YZmfy9+5q0m0ggHcuv3NA
Ne1Is6SCU4QMF5PX+FPWjLLdiocWoLr4+O6zRfSL9DRi1lsWgImSFKdFxhkbwZ+4
/kkVHISyNtNn7K0v+2RLEIQuaQn2SpkFTqY93fswCBlXil8Is5THvXNOIHUhfsoR
p8f4moybgTXRrlRgtSV0Y/kcj3mtjtc1vpY33nRE7pfTClXVDrSMBS+QoHI76XKK
3B6sBAAFT5Ta0Dpy42JuZ5PkRKVj/ps+ag71hI1ZfrjXNVi4Ue0RbaHXB+FYGdD5
hwDk45yiyju1ZJWEqA7FSeSzS9lmzy2KlSuo4Z9EGimt4VP+SNPqKhDMvliceZNF
hDk/CGjs5FwnxeymcuJzgh9/II/pRdJsaOHJOqdTmDrHEmcK/j3vVv49+sxa5oxk
gcWZ+mZthQwQoSH80aaO5xzTubQH67h9eB6a314GSx7bJ2q8lqKIzHqaz/mEOv38
a3Rl4xhJtaHTmITLGlToKw3M53zcfG7yK1aB25zRAOoTO1Ud502R46MnEumEuwQm
MeDiabfGDNxGxV8XHl+USAdocqOilc8ALP2EwqPFj268RVrOjmSEez01fr7CopgF
lHO8GgK8busT0cT4kkYDYuXsp4zesw3doq7sNpCZOwXv6We13nW1amuBRFrCmklZ
FMAPYOkMd3xDnZ6iz09vMAsK2MYdmtSKiEQfF1gPLC1SlX3m/WDTSGny5Al/NMdX
+Ia9gEAnPV+DKTULIHDoTwAs1V2X79Xoq2wz0bLu3wKUSgr1RXF5nh/VbG61tb5D
hrpO/OWSPWlOiKC0AxwouJCpEojeCylbozlJhAVTjBSqY+45whLlEfGCRLAvsoHL
o4NXgF/IWOROuCtMQ6n1y2c1hj2INQqgyosJjq0pWR7bw6zRd/uJa1LsAB45Tsu8
7W5QM5tDg4T1eUET/mD6yrHxVuxe5QhCh2iqGb047RD1KVOpPO2C4Xg+G3NQMchC
VWz+Pm5P2LPTkv49nl6lPExRPN8LWx1MkCgRFhlrMxNYBz3LIzH6plbi9tOk0Gay
cV1Piaj4Gmkfyp7+2feJAKY5cfURUEryDIB9k3jx/JgqjiU5TQ7OUUn2+fJun3pH
ArDIjPMY6sjdq+q5u/hf0znvxH0Dbepp2ZMAjlpuPp7M/ZlLmHx4/7sNZzuS4xO3
1a+SZRHGI8L/mnyhRpLXpYCrctVCokzWGtSA/qA2++QoknESWHLmm3dOeMdeELGE
qmXksWFzlcO7dECJiRhSxqlqmDWH4ureSifw3CLN3FGHybFMUvsRbcfXebmFpMDc
X+2DJ2raYCIFSNQ3ikyh9O3+IAuzYWP234dvz2p6RA8eQSMHMfOGmb6+e6D4X6hU
fvkyl76jlSG/YIUqDwCbrOS2Ww6PKfRdA0Lb1jAy+837y7iDJwOCpiSS+hw7yPuW
aXQ3RsQD6oJDzBGxsiCtVED8qOxgQA0yHWe/XisqC9R82Wmwbhagcg/bcYYALWq0
N0V2IWIfLtGxCKxOqX6QHvklNoB2dV406+NsShVKrljCi/EIKpYO5rkBsmLNj6IH
hpn6ryoC75ZdnaNG5NsHfJg3GASe11uvSLkFdiCDCakl2h61JcBkIo+rHag4bMcb
MhNPEwrfkrBn+wN6kOh8betYXpBv4AOiecPEVMYWqwSGmhYxrP0jbLkB5oIvaMVP
HsYhZEBEZOwoGDElodZU2F+06ZKEBbpCi9dlfPx+Wk5Qx6oKPVBIAdPyXZUzr+OP
ZzfjHiaw1rlBrCxYJB+qOzzXdaYJshpCHM6/XYN4XhFrXwXvbO6X1q4g1KspbXzW
/PQaMpossi/tQug72i4UACW0AV0Mfa1yrTNLp6bF8HBaup2B5SAzKL5Pf5fOKYfv
JWNf3eBG1OpLbVFXjL7jPamrCr5VLImXVoIBLyQBvMBpFwKa3Mtp5NfJX0X5dNZo
5imTxLyFYVvXJDrA0aom24LHG9Ewb1ssVNLfIDpWUwbL2YRH7G1Di4/4ZGHtlpe6
YaYr99b9NlXOo4JSg2oeRpw0H135a8q7RC7QOJj82pMccgWC05Abr5t5cwAvJrDw
ZgqDMMOF7w2v3qQPzNVPq89uv5v4KmDqJoUyOfViA/zQcz6fhXzR/YNfTBRXuFdQ
vSq8gU/sqW2GenJ3JcgWPXcCa/mTx539xLOb/g6K/xikrKAqpRc5xZTjMRKbCUgC
p31KW3smgV42hy87JAQ+iEVVDnFJCaS62fxP5MFB1uZsAA7CGRyQihkjdKdywOUP
W9g2U5EdkygDK3p/6ephn+hrrxB9b6RM8R2OSKosjfIWuqR8Va9ueuOPlAqKIxN4
fqsdsXNLcFe2aAOBAAAwJh0zNiBgZz27oMOflGtsOoo2ghvuI/NF1PkAVFidOU+B
9bX2UfRE1XVvEaYfhkH0zKIWOGWTch8uDXrRxYnS7hj5nVBujRDvwvGgt0apOuH/
KFVXVaqnD2XuGVrUMWxXJPYlfb3rtTrtGOXNSDRJECOC/GR/C+qzOsX+qbsjXAKg
axU1tG9ld+T3Fz4y89QQBqVnGXglqTs3zYSegdHrt/bmnUbRvLPIkWwW+2yrr5jH
bmCxwFf9FAxmaB0u2A5eTLJlMctBTNsAenLxFCkQnaeFhntNH2Mc+BjYII1O4upE
HFYxNsEJyJmYh8EXwSqHIhL7b5wquKJorWtuekarlJEDi3kRJ99ZotG5yv6PV0dP
p5b9S21rJ1teJOFTOlKaZp2/seUrUTC9R9ztITV24RJewD7Pga1KJIHhkRAAT55g
RJeC44GGq18yu+ruUL/Mf3J7Nfm7tjTGUjxKhDmZSrXLmGB3w/itvfOoYucaS1ye
0+fMDDUGIMa9+iFrosu+2+gWteW7l1YV3A7B/XAv+PonbYcunnH2ZHKg/Ve076aQ
PTY5TelF73S3CTRuW+gbP3Qxtj46wbknp4+tlRSQ9oWC27zcVktjqMs849iP0QH8
noev78IC5yi0WC6k3PQBhkLezVMT4MSxVWOEFWf5FuTHnXomUDgIP9kbpmoL3hI+
RhYgp6teokAQ2nbq+jTyLfd7u7qusIVGgAOkbWx1Ru/WJNm1BZy8aNRUhUqgiWI+
Yl36538QV1EqDEy5kJTlvkX7iKowb2XxhkAajgJsTQgs6FbS/GER8+vN2bXcMp8N
G5XmOqXVsyDRvGsbaXM/Ff8BABlYM3WLt02N9RIVIrpUcZe05EWXJdyff6VgvgtP
7BuX/H2nrWKoKDxVzVirfuJUKTgZJK6K0LjXCyqFchqO2tktvZSPqHtD7nqhYLNU
lkHof6aJRhfH7oarEAZUY47UXwOSEXaHFOWzE5gTb1sPjAWuh1pKRIQWjOsrQsKU
3pMpSAuz92r7mO1kv0HWokA5utTMlltsOJ1tKdx2XAaIrYbxLgiS+bT2wYLDRVsh
fk5F+UK82+deYS9pkgSg8z9is0rdhbhiCfjTYft9DSvMRx+QbA+vx0NbXxDlAX2D
ZtjEaBzcZ7NXsudpkZHdm7ie7KCZpYK99VZjXPcp9FFxgKRHDh/F//RKkvfKeuGp
uKD9kuFCtRujIhtxf2814pMARSOyPgpENiNE1QLRXwXq0hagAS4Oficct5RCm1yU
D59fVqKg1JezC9XBmpYocPb4jG3BqWnPHp1RcVo6n1mFBEZdgGawKrUla6UPyiA/
pVOqC9WTzu2UMeiKiay4O1vTmn/6Qe39/78mUk2USD7niyA7DrAKcld74G5rrMDX
KLxU7SSYoHZkYt9NV7R8AvFwbo28sPsFBlC+RQVtGoeCf7Os+Yz16ArFc/ihc4UP
5vzTO1dQefwWKGjz94t8g2uO46tzrRT548Q75pi9vds3Md67KbO5s7k0E9ftxJ+n
do6yGQ+4MjyFAWppCk6E1ECfXZCnXUGFk5PPaYzgTjZznsMZ0+5+utEornliuf76
wOlkxXYSiGBau6ny6wmQZne97ZDfTanmxmzofBfSJ7nZiMLHEXZYeqfpRDhwUsLh
UYJkVC0F+4mOi3wfDL5qhyca8WbArCT44LGrEK+v4TbF9QzejtwUVdMDjVdo/sLU
dnx5UOilSDMa5Lu3slAGbGlNVOn9vNUmSV7thOI1PGheYFEcD/RQHaom2TAYkM4Q
NNuqeZC9wWoZJrD+rudPcFl7tMNr5LSssswLBUYwBLTvCHjqr4Phax8eyXS2qDvI
DkNtpZ7W2XYaKPv0Y6qkG/bAPAaBvB+m1gpxTBIHWs9kyBHNZzvk8ZaXa1dTvlOF
2ZnRCvw5Uhcl0bsvU6/Gk4S/dYzzXcQVJVrwprKqH5uWbn8jRSXScJWpBrL5GJ/X
eJbyf7OkNSaPFrNqth0fKE/BgeX9J/eJNwmFbrrFUnGMZw+JJ5K69n6QiQbeOj56
Eh86GDPjxF/qDKKp1jhgojIdOuc+nrnZNOEIWAygQiiFpkEHHKudqbQD285L2oLV
7Aouz+LH/ox5m6scHhV6GJvAN33ll/gB4NCuAfemPOxSSlYyE0INuVGaFb98e//8
rlOvvnMMFafwa4Q99pNoVCp4Hd+tBmJPUyEG4H/IHVqhgKt/+WU8GgdWP5amcptZ
ZPETp+xl2y9JOrlD7MNmiEBponX8jwqApN8lBMkIm091xwqEQNA2/cibTztICao9
V4IbSI0hoAHiyOxIPDoRKSXBaqnNj17EU0p9RrhdTaZFnMC5D6+DTvFgjubJjwyp
/1hq6tv8aFJeYjC0+nc7ryW1qBBkb2iC/DcLglCscru/9ci1GmBHE1F55A9i0hRR
x7wCOLTZvjbXIPohNROuUqhXy1KkSPJ2SpFXrH5e7ygIZ1dI8YopI2lgzujNG8Kc
Xh3tga3L73hWFUJdro2expeVan2tZ/ihQvIL86D45eHRFtn1IdLQ86dmrlBQ2eCl
1oDV8vrTf+ovpmy646y8UKncbZ5v7iTX6815KxX7mSIzktKLB26sPWnNwWGJVM6/
ztXIQ0jxpgwGfDAk7nRXiomyPTCX46vsDt/yKdwlDSv+QQwwXs5W9r0x/2s5stlT
nR++nhOP0xC8tpFRmjwBKdPQ59TPUDtT52VGFe+gzhhVdm9CItNekZcTefjj0Ucx
SS9C9ZAXKBhnaWjs+iYfBDLyDEjBv0edLAjxQxGY7n7wd8dzqtwYPZtl7cvpOpGK
pgAKv464cobNwX+KRgD7+exKqULf5vV02QWXNL6msoiqUWx6sMYY24R6ikukGIaJ
fDLF4I6bTcAf9VeEbQZzA11g7Y8wUonwITW/BTyzJqws9wmBEkrunXU8BKVrxJZ5
+j6IokLf+pw7wHP3mId4av39b+mTowsUPwucG3GESTK7pQzlbLc7960EvsY+uXlS
mV0vhqEySZI53hmpehdl8UvI7govc8hiRiDySfJIk+hhaJ3Z32ZUQw/EChUgQYk+
JU3uThHfRoJWdAfy50C+fSMgS1Cp4bGBWJZiuEX637hQfk3IsZ3lqqffplNUEmsH
pLvVhPMDUZl/fcodOc81gweYUN8wXuXj67D7ZQhx8H6yDOdVpzNhTo5ZyIPVL1dP
ywnyVAkggeVuQe5a9qmwVBBHQM+cPHZ1RZ23RBwHGKItIql46apA7KuPhNa4qErr
nXf+cTCgBAs+XRTEV7kKT5kqQQN2VD8mVzGDRz1cADutVg16dJ1ZUw6QjIC++i2n
fiqLh9R6WU6Q+9sZ705ZdlK8Xl+N+aJXpFfjoqwfydVwF5iJr1Ieb1+MBkxbrD9P
GkpJInCkEH+606ESPG2rRsNMxrPHXJLEQl9UpvRtGNqrTGxkxJt7Pp8wdSqIIXEt
YPpDahG93Eygsajkr7Fc0ofmnc+nUWcMpmNIvXijwaWYAETex+ytHOWLQE9uKqKo
T+ssqa33N+Xjx2g01FEP03KLT3SxwS0cnvPlxv2iUjDDvMdhw4kQhqltQFXkTX+J
hCou+V3QuoIUz7E+oQbItPOGns8ikTfHyImSsoSd0phN3CpG8fn6uRobk0AcjbhI
N6vu1rDVwWI+FPKxrLEcb1kgtG2DFf6AF3iG7muDcBKzsH+DxnNybwmQFTUvXViY
`protect END_PROTECTED
