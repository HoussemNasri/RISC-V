`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CL4+pkL9VkejZH9wxwjxx9kbtdPtzt31nNGJ/2D6XczTRvh+cBMxb/8H0ZtHaKUX
sb5Ohibz2Gbs4VPSFjVHJrwGvl6d0rdFrOZYFDK/cNo2GMCe68+T9cMqJ73IC/3O
KwOBf2fBGzH6GWqrFa3wgTIqGN5saWDE5g3nWU3YR9/pgQdQG1ksULrk2r669fup
U+2axo9Y+OIRIvIJPM3hJj7LlPlWgXSrU2IXJccR/dTUI3UPxcYx+UiEYEx6iCdb
XuCqGdjUaumhKyzHQsbiT8GSm6PGCvn0XYHgklbGtXt2TywWBB5d9IVo8SgTNOVN
h939r57qJasvQRbqLl+oUzC7Br8LJoUPmlc+hXphkEracspHFF/HptEu+CytLwjj
ethV1628sw9dUEbBlzd4XwyPrU27TK+aFW9s9zbmyAY0T1OrrcsP+hZV1QnGPIg+
e9JYl3RTqd+ngdtBVxEs8wMcKFk93gCSkHDsqWQ31rw86jKhuSMdBj4BjO6umWWt
0s5cYdW6ErAwppbs6yyZn/eK9xIq8ilM4Yy0LCnqaJC04mln6IrrBUMl0E7cOW9S
ObpB5IIacIhGc9PHa0gdDXEZYrj5+mKUCM4YL1oGdN9l58gR98Ph+nKOGFz2PMkY
EpBrQmI7TtU74smFp9QAZANfZSDwzLXrbJ1nMs9JMv8bznQo9qQpVvEaxDuPt9Cb
ohEbdfYMO6KaBCS+GfQxekpfw28PF145uGelXn1SvNQ=
`protect END_PROTECTED
