`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zmv8S8fMHPx43gUCJ24c7XXGexxlmxbqd/t6XejoBp8GxqEPWtwlm4qKYB5moC1J
gGjdv1kLNfv9e+EAlauqhcEniOf3z33I3wlkCea7v8jkiWCU9VLvNJonsX0FN6Zz
zelaZPooVr5BMxIBTiS83DGeDsNjrzPl+Cl7uJdunlPy5klRk6dKXgt4aD19vI0q
42k7VbTU6j3q9C/RvcCTi3XSIZfTt46/QtJozM4rYoHo/59TeXXA4KiNUHuT/b3i
QF2RCgs1iwUMX0o8e7qmnE8oN/HYAFz6pOJ9SQCGV8eDH54BLH7A7XvpvUdGLhOR
3SQ2T2Q9V6I55I2+pK1MnwEea1tu6hLyMphE6MK8qHjOIePYwMgjbpFU5dLRqJhU
MkWuFvV7S25gkuXBtGg1HemIndC4MazS8tijrqH/4qwRkLWc+McmEXIKgorPEpRJ
vSdFbthTXUxJEiMmXjJBsiebsNTdfqkZ+j1mAuFGlfQ4kwrJKeSObOMcn43o5of4
61SbbG0SNw0h019DDMTLt6Tej4i4rUFjovsluAe83ruQuc8F+/UhaylTySIxvSbx
13YKC4SfudSE62gNgvX5AItynVQsm1vd1o/wsI64nyPr3rBiqhBFMiTbErLgJ4Wg
5suAv+cRn8UJXjfLrOyGRDAOgV0lSU+twBcOHNJaeA2+3VNPCrfY4qnp92HWFOgf
4/4w94MrA9Swyu+dmSwj4JL5EsM6RMVXw70INIrobqTlyBfA2GBGeHqDDReWOetd
fWZY1Yz16EWP4q58Tqt3V086izfwnxtqf/W4dD8smQSVlF6hG9vhj9J/NKeSRH7g
HsPP3USGqvAXsK40m4b4LJyE69fNA2Dit6QU6ppy8M7VC9cbkleThtDG62F2S1Al
CMJnbJWEQ7unHdudZss7Mtq/1HbFaQsYfP5GPZzD8MJ75Qv+T0XtVNK4vAN+MS2W
vs2UxDrUg9pAGe9hymYT2FYXHFS5PpjAkDxTdE64ZdYWrGTmilAsXLHDF2TdzoDN
0mxXbQbSGIM+Lhj30tw/mZ2ubUanwh0sI77BJajiXpBKzcejhcOHxcXqFSw9G3oE
KN7GV596I7EXGouu4+lQdkn4HOnmI/dqXh9aYO/TP/k1hFhSATMsMcNv3y8ZLzd+
U0v83560fyilWT2L0wXuQ6LkbEUbNCsj2t4kgxjHDm8LRv7GH0/ikf5fsbrhpUgw
er70sGebumk14kyotx1R44DCQbfIOfQPqhfhijV27Y6AdvMGYKfTqNYghTqi84iN
fPr0Rus691rpMb9ipNC6++txFvPYTMUoBMRpi0SgEAAs+EodFixKwshXounzowsL
Z5lC6wwCTXjEk22dITCloqiI0/pEUos1W5IMAv7YsqnbfknovgvNUZVsV01FV54M
8sZCm07J5LeBCYWraiLtRGhG91d5Fr2KePoGODV4vLWP6h+96bKtRUSPznza4m87
UXIhME25KYfozS2rKE7+PF/v/r9KIHw+Gf5JSSytJUbf4nH7djwMlFnD8VwUlK7n
p8y0FCY5mJsSWylER45w+MzaTZLLeBtOVWW5vyEBXgMpsFuAVSymmMbXhPY/Gv8K
XjV1fp5TE9Tt4+gKn8KFbULa1UJPxDT5uhHjSaJaW7dtxH+JtJhvYHnz0Eon5hIZ
ShZXBa861sETF44jecmsPIUmHtXyPRkEnBVDVyP1bv1c41NLiyvUACKg29BTAplp
pm5S7b7LVyLHdCwZ39XUCXHSXE6uYLmBNFahUdpLeXOiyWBXMUJ8g3j1jcYDOSA4
0wogeHSaKia8bkm0L8OPxNFO3995DX4BLNP/m/fOod/7wkY44aLv8enQnG84VbZQ
bTOhby8YiLA9bN75kOOjUDTvNIMn2ulRY+dnYTU9Ob8Uol6o5N200C4Hc5HdZWHZ
ssfUa2AtrK2Nnf3M80HShTykNTSB2TaGA+TpWOc8KNTt1qYwLinOqfGWC+1B6+Tm
02EBnhZD0gCSSSM3BpCFvq8KEL59dk41MwzuG2mZqOAr6shTx8wXRxQvfPMfBxzu
m9thVcQP5JvinP27zawxyRG0/b01cJt2TqAlA62RdJep1M7/PgP+in9fHBdrkpkc
o4KU+yPGTXSi4jLyYvOA0h3jKlNkzeV7Qd4FBmKRztx8MibISQxOAh0eEGWCHiL/
uKOerwh+Hu1BKyv3sfbjVCA+/CHtTERVDMq7smVH23KrIbyR3yYDotzETqL4EzAC
Ubh5APiZOQVbpiDAtjgMO2ZtOIMRNjixO3QKFm342mivS3L5ZQcJqcZGkVzGnbdW
NP9MAWxEzhMV8MzA9I1iTHs4NCjxmoQppLnJ/cxlqK1SsaGjUcGLkMYY2wifRsI4
AekKUVphb5+F5mgc2R9H+YcObNjpUQfsNsdaKuHepKLsYqIcrcZAmbZvy7Rmkdql
El0NvRvQCGGoIf+ajR++H+ZbawYWtfXKIbZ+0yvNPFS4MScd9c4XhBGUpQseaaQx
J6kyrOHCRQolzqs0C7IV/ZQZ9yAQ3Am/PkW1E1OBDmV1RTXbG4xhVkmniSeMmCb0
rckU52tnT8z4hHhnagUAwdJAFr7GVvvabv37rzJdNXR9o6bMcwdI2ZSnIM9ws9FL
1ud2QIk2T2vPU7PM4vKG3KJHz36Bfx0VXztUQQbDBogK5+1hqcS89cWyjBTI9GYM
9mFC/hdJ5THwrBvC5c+0dyz9+0xQZROTJo1Aefvob/Rf1GOg/ZPBCJutIsW9Ws3f
4MsiZvQ07/1SQKCD6bRP5FGZXMhr5Op6YtKy1JFAYWfRWp/5HxhU2nZCA0xkwcfc
ncKZV+GnQxH24MSmsdRM1P86TdnhJlTWz9NxzTmaXVMdI0W0mZyBeUGumBxzvuiZ
5Tf3qEhYIb10QoGZTAr4DGIKJoxryRoCbCVnhXN+f3pXgfeBK6lxfrOdXnJVUcKp
VQOyItPpQ5F10KJ+tK9F2VQXStSiDcN+ZMccfqLJKD+cX7GSRtgeTYqj6PyRB12j
OD7cb4Oh+tO1Ob4ePWVOE1DXvDBcXoVzpeJu+JZmbZK1zbPBx/wrJbUSA/DtQcWQ
BuR4p4dGifZgIWIeMyqrte/wj8wPxfikUOZ/9VCPDzwKcdY4iOHiKKk5/o3kAKEg
/LaqidN7BiHaXkDW1kBU4FMPNefYORaWGQe9umG0eO8y5fQmk3zKeIOxf9LSw1Ux
xDId45ZjsH1zg1oN+p0OihFG7Mr0CRbI3SFcpZkgse048ABpdncENG1BWy68nTSd
lRseRowT+PVjuBpnFpbxh5n68xxisS89jt3SQoYu6D/ZxtqIbqecoGI0MQw4dS99
zuNqb+E44JgeEaXEl9KSW5VqY09JIqgkAdNpF3KCTnZIv4Hey5EjCm9333Ce6wNc
nQGlbICiZdIq/80TT6Y4tU3LZUqfdvfHO75DK3THcv2ikIWZn/HnQtLPLKPFUpNO
+Ysbj5wUm8Gm3HSJkb2wVOYA7a6O78iDp9G25c0uu1/IlsdZQIupyvXKopJwszAH
TY+loLNFwdWhUIeeqi2/azTJU+5o1GfMhxM5rYewO7+/PFQImsVHtMEr5VW1KOOP
CwZp646yBoHbYPFLkAT2lPW1SH5RunCmV83rsT/8wSA6SiyTGYl/Wgru4CmSjT3/
WLuRTjfa+i2GDIJkODGn5szfzEaCeBvo6gdwCdYMQm92QhGpWAT98zLMDT6alp0i
rqY2mh2TnFwkZKiE+jurqlZD3y+gcZzPhRDG/uFTzXn73k4NNVYWJ7NQAngkQfmC
cU1L0lrFURHhXXCiPbtaBZPRe1LhuthGL6DDsvLjg/9Cyb1Jerz4g7u5ypMO5NC8
XxpB4HN7hI+BzTPqmgQUCkZsvywp4juJQn3TzBhcqM5Cs5ArUO7a3DIeTmrvwX4u
A6SowB37m4/zMfBsKvNZvidHG8mmsrwL9FI9LPACSnihH05ViSH3+payuCbMb6zA
Mmed3JDtObrrkt6VsVraVBVt2O6zvvhr5o1LTynpoWQjzn7dGJ60TpX9yEQ/laL5
Z9IsjAbBQ67D7m7YpSC7W4DfP4g58ekHvVgafLCXc2/5oa7wtWu2qEB2Ex1d1wup
iaqwVXkksCYCfZVCjdszX2JSMPz4ZbsEGCBOGbXAuoXkTmaODlBazJHVxFZpby2m
J89iZb7Nde3QN5kiYUpT6FRCIi+mezbwZAJdHhbVmZXEzj1Mjyn83ycnlGmTH44u
aFyl7N5PUyN5En4kKpBmx4cRRwNkbBqGc0RgIpRrY1fEmrsGz6dYJQGKWjbKFZ9i
BpKoVv2M4nuysbI/KgVG8DH+F15JbXjLlk4+HhAThQJQ3cKOQ81k+VZMTXpg6Vu7
flZZx3D1Frc01JZvvGY9fbDflnqICd5WMoldoVRbX/1sfUzP1ykCmBvlZ5d6Og+N
HZPPrcoNF+eOtCTlH6a0/DBgs1d27zzdUCSVAuTuVn7jB5NqO4OCg0/uJmdupKn3
ku75Rh/UjF18QSHAKHYpZIgzpbfaQSXPl4nOzBRQag7TjCMKmlLRrH4EHO6XwoRe
XiQXTEpOuipPVEccOFV8x/zdSdtmjYW9PrDemF69KVsB9QR5xrJ3Ow+0aSaZvOiP
`protect END_PROTECTED
