`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HQ0hCod1lJoGJP86MPZ/CWS7iyakgK+PSbWVQA+H7u2oOumekhkzU+rIsYgg8Nmn
0YTRDKTlaPCL8hOT2ej7LMiyHudykGCLwBk53tMULN9w356uHjCfDEid4TsrbyE9
CCLzSSPszMXN/cBFofX5JEy7KMYIk9ohnuSfH+5N745ZqdSIdIH9pFKblo27DMLS
ZF69spO1v1QepV34eIHjijlNxDEr4VTgJi+7DaGLTa4ac9o7f/SLefqgtMERRZr/
jeOfrzWL3fzYAsVDY8Cco40F72MWMAve9UlXzBv6CDCMIX3AuHbCOOW20aAD0M4e
SFLCDbPXtl627ZD+0sZ205y4BXan4NrJgsG+XyrYPSNLJVIIAPOpJRECzfS5+j6P
bk1A3iFVc58hIHeP/LlXZIccGRyGGv/+869zyiLknuUenn3xG4MXXd9dOsrCtT2T
qoYAfMFGfElTqs7b5Woj45ngoI7FUV66tLkCllPkUDVIUxT6q3OnAL0pHoPTxr8Y
ruUNc7DiOlTQOq8ZhQPE4S2m91Xd/0RHtN0YrYYqhH7oWELg70UTP7Ja6bt2zzIc
pUMgeDPSLhrLOT1h83Zmp5kqYxv8nMUDJ40HDxndBSiuumCldyQPHwfY7dwGI+BR
HremXUySvrDskDRKs/7X1m/QldEd7vq2t+zJ7ly1n5lKUy+CzMFrtGP4ZXCQZi8u
rJdvGBQGF8ZA9V2hoP6XWlRkNtIbxctK5w2+ayoqbBSCAaHJnit0EO9iKYRA19Ur
nJ2M7+DrG5OHuj2ukGJvXVmc+5rDBatzCMILGqxjhx8ZQaqivSAaHOet5gDZpVe6
U5d6cPLeCXkGlUdSVGhLsiNYHmQCoLLeLu4f+YYjuA/hIyvnvERzGY03lmAJApAk
560xTrAhrnJGmvnxdNRRHRC84+e5qIvsN+EmCSMlublvL5nW43VfwseockUAotJj
TxlnfL+xpBpRdxqMhM/3s3abVsFaizvPCO8hYQDLBdu9HF0kwrNW6I5vhsrzVxcY
QyhiX92L8DfPT+7vzmnn0RJVFg9fUBT9mHvw6JgUwde/xbjHQgT60lZThibpaT4I
DWU+teYABZ0lGyr++FNFDB1Ld6QAz7K72rFeDmeRdUU9W4nIo40Bd+nIJM37kkJO
TNnIinjHIeR6B3a681j1nXWn4oQMXt9qpuzSfDfcpAmwL9BZGZTj4q+5pk+q62lP
60jbfpEC3Wf3WGsv+OLjoq1ZVmDNgs+vIIrr6Adf0ynHME6oR2jqZVxRdP0D1Hbe
KvkvuqJH1Q5iAfHnWFGZTUN13+zm61BIC9jdQSzydbI106ti0NGpSKPG9j12uC4v
LdSzSNJttTZ1LbWFPP0mDHj0Ct2ywD9GLoboq1q/rTHDHNea52DsULnbqnU+Td+T
AwtbRQPmGSSZhuByvwH4qbbmptg4Gb4wG6x69lFjryY2GEBc6zxsTKq/01PYPDJ2
DL924dCgVCVlvl4RtXG35qFH5gFlHPkLI+jH0tzAT6odus6QcMeH0P+5f399lTHY
L7yu3dJRa4TtvsHpVGDQOgSqohH++8T2XSB9V1JCmycF+6QKhIawXXAq27w0SEaH
9kmraRRErgB4+Xoo+sbg9l/scYg/Jb8mEyR3VY++GKse4lVrh/a173F8qeyw7W0o
4edlMCczPGloCeS82hnR+bQq3gnOYqtVgrHqhi0vC19yHxC55GDUfM74Vy5VHknM
DGgalsYCTXOuZNPQjB8WS04dSNM/cHcalKeBPIHf+slldTIxvQ0mLDjMcYyJCxZ4
3kQA+IkTv0f8s491sCo57ccD8LK4OdXE3Xel1iFQ8rIQKj3oDhG9Fh1PPS8s8wa/
BQlWr3VMtqsyyEfVcQh60d6U/WRFGWUUovDsYzI8PYlHzpsOIKyajr+nVtilRKl+
VhtGRG3PWm1uMrTHdhKB5jsvCzR7ecd1MqdTIzu60J8zB7OVXiA2F6Xf0zGkDYIK
/4x+VaXbLJT3GNNLGhUvi8D/tUs5wriorD61zxHnmIaTmoBCZ6B/YtSrI6U0rm2D
q2qjCikCmKFixIh/cNZmlQi8V0KD4yxmwaQOhUnB76KJqx2M/NDpEsDx6Y6z0G7z
reJQDevFX84RdEpne9BmGdviHEWCr/jKJOExB+q1ndJL1rQNsGSWGnZIhWRYi+DL
nugps4fYK7lDGXMtVVsErwF4UUFzL7m8L9jpnBxHI48jJwJ3x6B2Za+iKW34Zopd
xTdcDRy5ETZIRm7vRPLS4pPMvPDy77+er7dsbVMw6kzWcJ6si/o4hKgc7xxNVRBa
POa3dtw5pfEoFP7JoUTI62KgdyMMm1GoCJ5udrCqEAghaLwDCSR/+Psu6pnpnxKd
eeAefXFVhjbU3O+Q12DAviPNxumc7rQo/qdlaOjrQxLz/cfK09bvWhlJuYyLrZ4M
PRYhQi+HPPrtG88KrdxcNfxJXWf/qbKCqw+hG/XZHkYUqfoE+ezkXF04Nw7fEXHq
6ej/2LRFkD6sgBIlCCe5nxOx7KHdUwGPt0udJpohTX/jNxEwLlKyHQOFjPk4Y7Rv
iaRtDkv6jd3NJb52ClHeusCiHLEL11TCAfpfWFl9ciTCzsnQkMKsKUaO+Y+DjMOZ
a2KmqVR/t9da7Km0HefQerVbYCoIjZHxrfqKeN+bV91lO7bMGYbwad5xOvUDi1nR
GBu0dN9P6IBPt18htlxR78ZeNBpWgfyCUpGLNVpipx2L6nR7yssaZf1IbctOR/Bf
LACAU1jfJIcekUQEGoxY+kQOlTyXG9MFzdS1Ix6TAQ6zs8MJ8bOTxWn4AyHqX03H
Y4ZvTkDI2AzLdpqE8yr1AwzEJzNO/myKG8b1uJtd7JYcQHxtzjgP+7ElmyKnjc0L
0J2DEYA+iwaBOAcjyBJjoPRnxSHdKEcMngPQ75m7HRN6HF+n/NpMZ1b+eVTtRk61
uURTIxciBkiozY3+/HA7koQa+RjyQvSlthALkAeN1yehHQOC/QeB873VTCQcxI92
mmaFFnrUrUtNH6Uo7xqHCpjRRsKoK/CHLRVGjIJe5SKx2QblVtJ8o62lb72bf+7P
+L/Q+1/W5xVdLwakbzH6JBdOO0NwJsACbZWuGA3Ms6U6xveAWUu07PTSesA5HAYQ
NUHkYSXoPPas9Tu/hBwNszG4XFp4DlQfC40MWgincTQ8EPHIC2RL9uvSRcdAYdmK
nxTi09vmOaRn2C5i2m1M5+3b1ungoiP3ogg7kYJAdrV5XGWeD8xE9zOafDbXDuhk
mxy9S5RCmWKM58xwch8FFZVgE5VmNrZW2x4ieHl3pGBtBD8eFFLRMzIhIRjQbC69
Ds+b5BXnvB+G1ekFq0c1O8GrMD0C7BwNNTwehFkh5ZPXsIKHN1NqVl3GiMbUJghN
GyUlzspeoH6L+GdQl8y851ZXeuwfyjyQf8p3RacA78mi08iIQvCem17HnEKgYGB5
kSpQOqhom8zktdC2uauj78OTEHNZVL9V+4H/RGhzF23V7/ACLlRHt57NepJsEays
nXvLzhQ1lybcMCUPEFSztLUQLpNWjQJI6XN0cGEGlKj8EghuCtXKL907NOMMMDxO
XHskqAtjg962t+333VD+IJ52nnm01hLiUGHVKSavuCcLmD4roWcabUWhH18btXh/
kVvpv1pyHXGbtfVB4RDlKpI6w3laQ000bUGD+lDypI8uQHYGN7vojU3ze9UBeo2L
4ua89n58YeRcICDkkmOZtYxckoLoWykeR0Gi0GrZnOODKLOfQAdPhAtqDc+VT+os
RUmBtKUl4AlA7622BVxUJ2RzaSbV7a1Zj4ZMKQfxAIXzUkxQeWG1CBD+DPRG0odJ
YVxwaq/62XeaiDTDgt5Z56CWqKWFO7jGm1FTMtAJR1ZDdm6ZxiQ40/k63WrBaZ3w
k4GluzGo93THegqEtZ2iUerUR3Zc3PjDkSfEH2AelgtCJzewzvTDPhZkXBsaqWXx
LOImi/7rpeUnrqRUbDcfTPnQJnoZapmSO0Q41LEmhStWO5nAC4noRkyB47neBSpG
MBZ6N12GHXAP8WDaNlUKum1fJdDpSgj5Lr1vnKXDk/D0RQoWs8ZlVHMtSfKeM20n
BffwG5pChKQgHkZ5JrAQWBELOziwKafmPHaCBGKtf0PKX5PlrwlhVZA5UZFJG4rb
yjrxBf1MPOmul8CE68EsR3qppoiT9b278X7oBCo2ut9bE+R1RfVEsE99QEPiwexC
bL2Br/0/m4Ic5BljXeBUegSlMp8JC1oRgs+XS9x3VgrRW1R37aaK6dsxP/r+Fkzg
tVwdnem9gEKLFF7DAIxvtZ/H+7n1GZkhu+xKlKie8sdBug4TNf9YnJR87ku/XmeD
zCOkCmfB6eRYZcIB1t6RqfWTJfNOK4XXXlHpS87gDp2L7vJ+LIsThl/GJ4QKBqPB
HvPkO9HQlUYzoD42nQ5TAifCcArJaT4ZELnJi/Oofa3KK9QqINHru/fHhVIY4BuP
+5bjekSItXeeuYPSaDIFHRzNzNq/T3a2EUZLfxfrQwH99FAQBY8H+7yVmh1D/YpW
bBMrLpKb1XLVI0Bm5P7rga0ETnD8bsggSvhJ/bTN5n8/rGNN1u1bAk5TpNu3/Cm7
lSzO+JPUZa4apzFKLVQTQH6h2s4v0spF8i91473s+PG/GwLbImLWM+zPuJGbX9au
04f738Y97JublVXNx0+fMF2MALwGuDpV9avxsBf8hO+Yu+M0tf7YCWAArF6f5nsg
r3g2nBzGI3rp3rj98nmnbPXisCvfcVwkawzYBeIzZ1P1XLkTLaPysVFrLNOfI28P
rxTu1mrG59wlIaabQd4w+UYVBqpVFObonBfBX92XFoiA/QbnLJi8+snvXWJip5XY
Ww71JQdezbFy1CSzV77cyvbOtWldFktn2J/wvC4C5zt7oSsK2qqjLI7UZaLk4Agr
XJ0DOpdPgMflo7bgQiV4YXOYMkj6My6IoyzvzNqO2xn9F3MmDFKi2iV6z3/ooZZi
GRcvwkQox44I7+wXp8ZULctZX0FtoPKiJWpHJ5mb5c+27+O2uwvd968TnC3D5DBs
YCkDXTJ3hJ8GZO0a0Oqa9BvhjfIdeF3I/C3x4w7apGWIMwlty29sjlXHLTmnBgB3
Qf41Fh8ZEqRT/UpboHaWVlcusXyhBPtg76YQ81LsNmTKPs+lirEjKE2JKCuLTj32
5Tu9Qj3KHUoamDXZ2QODNeSCFpLgPFRizydlugltTzh5VeCaBQ2+fm53I1GQ2Ifd
EtGekq3EM7Ho3FBGeIaIbDquF7uspgLZJZBL1LKhwSgI3Z4DLLOVQ0GajUCptil1
gDJyv9P5P96XVur4CZsAnq1O0dKmNnMhepOnd7XGGFUIvs51OVc8ke9J9Ua2NMZm
zk+XYhIuOvbMDruzSyZSg+P16QSPsUR0LUp9R/mdaBz2cRgL2UWdRABbIwA/+ZX1
UMyUjlc08Ar8bbCLD9mN7LwztNqqJAX15/p5ILle2TMFC5rkBYJe8+tYOyZouGCf
ZIwgQ1O5UATR4AHokkP4L5dyQ/uKmUdPNZGZtcVfBWPuC6Bzq8G+/sso9AHCcDHD
GO7ZvAGTnde+lmMnr/5WN0XyW+EtEdHe3bTiQOQahja3YTVX+9CUnAmJZ6sHhVgB
nkBsVBZ79CPkf6s57ATbty1Ytep4aH3eUJnFL+HUfcJJtKUtRggyayHEp4pK4SB+
WPD98ImD7nF6tCHVO+a0Hr9jVvDfiU5+bsgOaS4XjyrX8ILBuTkxkLWSxe1DqsNP
NephAeMZTb/yoWopHMGEqa2p16XfsTdCS0vzPxLNgIRS12s9Ir6cpx6racs/xmq8
hBX9IsqfD5tn4A9YpdtJTOGxkAnWHDb0BU6XVtSQSaeRl6ysuF7E+6uKa3HYBRpi
FURhG+C1Ni7/t1FeG8JAGSccJc6Khw0olZwqp4hVx1kudHsHMA90v8yAgOhWpqYl
usZeOX6qzGpwJtxDPHrJblnqgPqFB1G5j6hVlsLD20Wo08Z2wvN0UB/HZ3oJdpLe
O4E1xg4/W+TR5OFVIu+Fdfe5JkZcBVqDBfuv2UnzXNNPyrTSxx4aRmEll6cGk+ml
4vL090+LafVoqwxaSKELNCuyvDT911dCIq0OZW2bjTGS2/Nw2XVBFJFA0ubEAWAk
MPAVL2vYpfcl2T4kkk0lPub4cOe0574LKcWSBHmHy8vJbuwlgG0VPTw8qwO0E2Xw
PlFnAvApkDgDwA5a/oDOC86VxTQX9lk8lUmor+BER05Gb0pio0LDaB2nbg0g3aQ2
pNfkYYgUmya8PyyYwGyZJJn39NsW4MlHjWo5ZCb1/gH3O60e10rwRWurtHFaiiGV
jqYV5pdD0Rva+0gM/yQI55/4r5L8AL3yX9WhMtlZsOK1ZOXGPFLjajMTFzsY9NOd
o8VKeSbKY1O6QV6NLN5C45jT90f4HX+1xBYC0xMb71QipZLOTABgbXJjxTDDRfaK
Xz3tyftDzoccRO6peovMN7V+/SNgRscwRbv15CiY7qMn7YYKK+0DdBgQgOwQALRn
X/rc43ryG8c09l0wn+PXDH7G5D7nliJVrpRk7p4W+0C2GLToykASRbz8rx/AbB3A
T0kRy4eEv0DFt/yMWmOb/g0uBaPPIl4zqAhsRMKhfyRXRsNN+Z9u2vXfwWRZqKa+
JYdlvXwhJttRpUtN125v7of5OCOkX0yL3OWkOS8FsYi+qPWkmTR7Htgl7WKURgrK
tBFeaZw4ggVZhiIJdM5N6buzkjJRqKhLNbhJBPIyO+dSCEJoX6RnKVvDGp67BHWG
mbQDR9OpIQvajRTFJ7k0aPbu9vKZH11mVIEtVdav5NFtiF9WoyG+r48115xkB0Ez
Uur0AjFDoGpJuh/RPLZXH/2+Vkfc2C+UVGrxqRFi7ZKCSpJ3wFMVko092wkeUp4Y
QqIMPvmeMFNMDT2DdgyrO6/25t0Szgt+dhCS7YHmLQO1icOnIzHEpulTfYKCchTn
qZUvmxaBhOj3qQKJC5UoHo501WAnpSeFXVtcXn0J5Ia+x0MlwDIZph1HtTXC9JX6
2OtAGI69In87t5aRiyN4AHUoHoaYUL3FDZXeIK5BISkM/cPApbFapdz6eRd5t5Y/
VC0JblQLXoqa2qURup7WqHbbrv8r8dnwnJa4d0tV7m18Nu3Y2QTcfwcSZkjtbjQC
G2LKnpnEQXRbu35bPqkTcaz1fa6C1m6ls/9CPA45N5ARGre9UUIAahq5ZRQ9Fv1Y
Y5AULaZ+mX1gqTGfoiskDFzMSRsa7NOoQ80LqLQUEuuQhtI0T2jWHESvWp7NX3AB
rRDt+fJheIi2wi9ieSiprb8rixEVcYRqtXlAoxyj1EGL96FPu+qaO/ziQynA6aUv
+zq0FSP2iS01Nd4i432Z0BjnCHw+c1GMt83H0IlnG1HR0ET+REqONwKsh1QGVPkU
LTihdSLn6EcesEQU3omNGYb1gOeONjrenC/uabEzu5PtmqMi5pgnh1/Xh4DmHUq8
Vsx3kRM5/Crha51oPyk1xqayx5V2p2ysL8h4S4MubrqDzj4+nMLEQwwOTiHP3DWk
ZT/2TSbZVbZ4if2wUBCN8RzUPf2HxCOLb3Q8Srd0TK4UeVPJImph0GHqQbMZE9DY
K1VDFgqYg4qP16th7t5ylI7zO0lL4l1irqGuitAYzN1/5sgfzKqlRkhtCFjXj3C3
1wfdpJR57cx3xbiYkNQqL3X/UAYG3KqUkDv/mRcXSdnoPY7thIpwWEsQpdoMibsp
T+cYWZN9y9t+/8QnFqGqfC1Cf26O0Z7rCLIsOwEY/niZkbR756LWZ0cZHy31FzKr
lmURMw6XRXpDrMOECAkT60EG8Bevw0Runtt/6svEDelELnkJAflo2+j37Zs3Dafl
FILOy2sCbkCGnHdhPJJsHJtcTawMoqxXyPl3cQSjZiAZy2wStC1H2wsnLhbtXqOz
GSt49m/ek1a0lzNx7aProqCdcaVTlzOWf+EX5cgpmgo+3G06wG/01F5Z3svo8sk9
SdcvX7jvGScCaLU9MOZ8F8xru8uuSg+ou38SdRTFixU7TNp7tM/WZOk25L4kkCWh
hJnI2/AVlGuPb6YGsz9s0td5lZcq3jpE44AIaUGW9JvKZXUTGmof0pXr0W8Ww+yq
j1fYn+ILWh7qbdn7SR/Xrs1vos4k1AUV4UX3unVDWB3vbX6Iy4HAqsLO9scega9F
plyd4oF5UsF8IQozOLzgyk3vS1urtoWmcitGH0N1kFdMlGV3YXYtRFcKQUlzzTMH
GxEky44SU2W1Di0mXYwwX41/zC0YZH/sNXgGWe9Da8IRARu9pky4NQ08agc2GsNV
Y3B6XsYHnuvyFfBGvnN8Dkebw+SABT9da6kJY5yMu3wO8gSXeNohmqiR4xKqxQI7
1vXB8seN73caY3DPj4uglc2FR7IHmerDnYtFNYZgoiQJ4lSbTKVBl0VFH5eWfTv7
/1MWl44z0YWLv1DnMsNsjjzvzBmyk/8/JXbNWU0zUvssCAeM7u0nnvkaHQH/rH+1
ZNDQxzRBc156sIr25+eP4ZUWObVXfJhZcd7T8t8VuOJwgE1vdPmXz7fz1BvrBGlF
3usjCmjGl03xS9owr8Lq4zLRXtvOXyYz5iHL0i1nJoNLXbAiObFwvaRxTkGq3UWt
TRiNIRaljO68MSRu9Yw5D4n9JRNIaNUXOREuQVXlYkb10btP/lHErwk+KqEfivj+
DB7Bot0gKRTHwiy/F+035WSEQPvNLlo/vO5i6TJl7kYDniKT4ZS+5Ys1k5GK1ysX
W5vazRDYW+ibLpZwi+g8WTes538BJ428KaYlassuxXurmglBzSeqa5Qe0UhhpiZO
EKqyKXJxngBUTPLEKy2At1RiwmMXJSaAM17/9sR5DlVAG2kzgRXkKhGHipxzp8j1
5nQlH6iFWNGOz1r2oQ2kJJ0iiImJtB4INAy1B4NoQ5veiqH1yW3V7FjqJPWsP5L5
QntGKCzftJ5DrqtOdZULBZH85fBU0QQ8cTEPAWgDGZ5TUBanys+IkCk88P4xqy3R
zWZnlhlWpLgcCAtVajmn+Xb1wK6wwMe2/NI7fg/jr8HvXJJDCatrWs8lCl600TYg
D9DNIlAmJwi+cvMkgxQcNuFtA7eJAbgkTCW3otqoWeZM+VVfpwIhv4ORjaJ1lIr2
QiwU4hnYupyeUGT6je/V9EaBbxxKASmBT2VsVT9p7bWyyQylorsz3MKzSS/TS+qh
6zPXxmpKZrZtxsvBvOBxmb6JU2BAvxpt3aJ38ksBpLSEVwpL3we4ngmXTnmJej3K
dGIE36iZz/1B8q1MW1HyNqdqvz/iY/qh7Hisvfam+Da89UhWBjhMfMmTCFB7BlFV
4Oj0odHOmLFplKczcOVxbTKzXKsWwYaJyXzWTBtWstj0wlPp7wMWx7p7DVSO9WWX
AT/LwXskyFFXQFw2iwYDtHAIatHm+3GVbCjunuuudBHs5GYys1X27tvHgePP/JJK
I4FvajTL+WtlqUbvGdAW+9G1mAm28TH+2J+xLIZcRovxwI44Ue6NOrKMSt5lB7+w
0HhlLGhlwHT0haR//ft6Vh9NkkqasxoXquABQ1r18RuxmQIRUvQoKp5pzGqIbc/5
2H3nWaWYY9AuSEHRDHVGvm/ZNcF4Vm4p4xctAgF6Bs1q0quhdSpD2VcgSImF0pXN
q9Lja8xXCV8J64X8/N/r/90/usV4bv7T3/oTVKIzMnIT/slGfYsaA7RTHYhZ1Mv7
b78fKgXWqqWAxAiMeUMyGVy3LcdA6FiWDKaTpavd3LAY8LAk25FQDF5yeDf/HYfC
L/U7CQDTi50xICyudHZMToGrDbuSKecdO2XKy59acyhMTPAjv0+tw49RdJWmMUdq
YHgNAFJxz9jTviKF/Imc13Ij2KHpUt8v+T9wpbboZYUHzYvKJ5UzMBLZ2e3p42Po
DIUA3I102lzg6rJGh8q/HTEs+C3hhZL462+Sh0qbkMo77Js9Lg9B9xSyhvSfypWM
JqZ3E8Wg8l+oc17ZVl+5fr4M6j2RGxg8E4q7xpnD5LAYv543Eel9uqxOReNyLumn
ZQ/u2L17SdZdnAfmH79BKe9VNjwbYW9+50f83tGZ2YQFTQ8sQlA1Gn0U5PRsvnL0
HH/GMOH8xDkqON0jNlUQqEgzjsjhdQ3vv1iUJIJGNTc0/oPseMoiVZGx4fLX97Kb
12PN4CRWglbmewuLbAz/+8Ln81leyWRrw6mJbGj2Exh4wi+5nxJQ2JhDAPowfTdX
2lxS0v5i7FwhT6iJI5ZMQQYbAS4mRpajZOWg7DU+eL9PtJX7y1vldeU0dXVBy2MP
lBrU2DwhzPvmUDCfYdPMFm4qkYPyeEfQnTPx67eX3KA7F+ILRxE26YPhYr+0JxDS
mUzlXL0B/6jClxygclx89gDZfMYkGLsGf7b4wDzhKZ8SimwtQIfBeMAV6CWvRDWk
n7Ufa5ypkPa+JWqOhiGWajjD9LM7iMnkbe0LIigW5sV8EyPU2RDpSfFHHVhh0xP6
EEZ3dFtAbSYDOU73UAjtX6ncUwzqRT0kE6oXHebHqPueqvV1sIN8KTZ75H+qxI4Y
ICUm7mZf7rdSOUb4McB2S+3/VHBUs+8o7IaSzRnaVuO+N+6Y8wAkxa1cU9YTdIo7
mtrooKJJBJDndJg5RgmUdwvJLjRjIXOaxFOmvEwgt+bmZDLUDOwJgw/J59mNttzn
ntCUHqTV3mgQn7nCpknzCq/xvva3uTCgAt3SnUho/YPh8CdrflbVcsrjvF7njCNg
q5KiJMddB0RN/QwJvMYSmEYHuzDzr9tynxPRe1vxhWd3sVmqOxzJxAdnqh7JMkpM
L0Vm6cx30HIQSgQUThHYupSOSclL0TDRss9cwRMWi3dlLGhhfpmXQCXdZxF7YKQJ
pwcv0EjU6C02K2x3XCaoqbp44ZH2nshGCqZqweu+kSX3ixzdG8Q00qcwyqRGAheX
ml7fBbvg9XGIOcED4f3CJS3eOjNsD6v4FmQbDco9f4zjBleAvIlHZBV1ELtnyfgq
UBv/S/GJjNXwbxGIFY605AAgDKmERWZGlOGPcXXDqXz43Yu8uJ2ysWpNWf0tuPH7
SCd8hmGzLnmMBuTqhAAhSadiEWIEb2cAA7pwCyixLxdEszgZcpw9rVap+AUz8yl2
tFcszqMua+hU7u4q6uIHMIeAWIttIsGVI1L3OcGZts9qIOtNsgyTIeQ0jy6LT5IK
m5c/NjqPlxQqlvAhKX8nVTKkM0sTFg0SVd/y3MXNBkHtaNTf/wOYfzk1G27Zx0Vb
73gexCGyV9zBmpDqGQdw0RbM9HP1VmVM/55j+qf7SDg7Z2b41CBEuRXb6SJXxkiA
68TX1V2bY6xfF8AGuu6sOntx8znWJrWILe4czr9cr8wt3wAV4uohrki/Of3sPlqY
NW3J7oVKwgiGRAseO3n+OZCnyQxBQaX+JmF3HRbjy/mPxE7CcOU+sBSrJNlIW/tV
6Ve7hJpP++8xZmDN8LdyBRbn90K0fe4HubW8LbpaTgkh3RZ6cLrO73r1g6CFUn2Q
FYObDfVut4PV0KaNQVmnw6pd1MarTpEtBaNt+/NszD5L7hGz/0SXn/meaB0XbACj
qnUC+WU1D2HMTfjoxh1Xt/C7rebgi2qfj3giuHTj9jVm0XzjNcNBFx3cSFzysYDZ
+zKiOkMhcYlb2O0g/yJ/ngUXdRconG5fy3CJmSutdgnyy0bPuOPP/pHpO2ukKPIX
oBVw3T1wrp70OFRidse1lKVNTfo4r8J6oElGlt9/cIXL2gv3WqR7B1vJJe4m/BbT
kfZHVVhEkJadms2yMZsUduUDkpLJi0DFELdKsa9k6WjYkM3GXmPt2HT5utXAAieD
DXKO2ezg1DPZAZTLv0bprsscvxLRBRsYMISG7PvWSPmX6O2QNMlfUAbHOmPhwxtQ
9EQLR7MnNUi3dIj64XXfD5UXFBX70+BzEafs5rXEX0PdSht3No+KwSQyDXc3jFZx
TYAH2zlDbsjzww6LJZqUCOvTHW5oYwX2u02Dj/VHGe3Kc/n6vvc+gZchjWn/PkLX
DECwwbp0zoIH+hbWG6g8V2/lQ6qR9gKSc4FIJQnRN8PCftMUL2hAfYnWCzlPAvYM
SDWPhTF2DwRg9xUqmlIel+w6E2D/HU/R+xTBbmInkgRTzvSGmAku6U3WNQgynkl/
e3nNJDHzOxYg9E7aiF8QBX2shsqp/If9w6E8SxD4ym8wUOZ5rK5dOpRjfPLytrFd
UCYGR3zbW3H5l3dwm3cuesDlJJhTSgQdoUm39biWw3saZVkdrhbFcWwSqmm44A2G
kyvNur2i8C1VedGfst+5A1J6yk+Ip/wJt1u1tcrvI9JWbKDaPeoSXiX1oxAQtNF7
YxwoWlbOQdmEO3bx9vmV0bGaBPJlkJtclx7zFdiAkjuzSCOxTl5oRfldnN9WaQT6
cHQMti5+T320XUFFsoBqPTSIfZYV9djX7abwFk6xvpJXC4NeMXkQ+5I92hVWDvWP
fxyzajXGITzPJKW2Db40YGKE4TztFttI5CxVlEwmPLqH3z77UCRrXRoFDhBYGxoy
LUCwPwvLkmeTWZJRhJ+9oHKeGLr0F+oxJM1mVFBWILtjYdYKmOQxfX/1Y7r6/QtC
SXCr7vNpo+KBSousc1RimZvmySqARmGtPO7YKwRioLNUzxow4+nGEOYW1nzZeyEo
+XlqTLIO6OU77H2MOxFASp00ZNRi81JSz6T5YxYYMEgYSnCznR3H0adclFDNhW9m
HYZFR3i8n8tLQUDWDwUhsBe1OOsznUDQWcaJHrY/aUFlaA/jAWuya8FyQIVLfL+F
QYJIF4zTT2Sa0lLzaWodWmyCCUVUQaunvfc8KLkGn6tfqsYjygVe6tlxiZXFAMsf
d+079B9jB9k0BnzIq6VDN4ogYwKuCBPrFCA4IVgRYy2T43UHggxuJkMoKcYt9NnA
SCO2UGUDAUAB81OB4sk3G1evVdAPAsmr7kuIF/U4rTu6dvf0vYqbCgLfdrwS/1kK
9ky9WIs+8EKxC6zRRh8DyNW13AZ9uqRhRGIOSFoIo0BvQeXJHfUxegCBbz/Gm2zL
CitES/A3GD3TzlfvkVf1MqRlCp2sqEZHASzweLKPnwID6xxHHBo7vB7YK08QK0ml
CDbCW/OuRpzgpYgYLqQlJIeI0I5Zjg1Ae6kGA+NE7/zVU1RHUCciNUvektsCr6EG
B6PiQa0qdIb9ebxivdevaZ1sO/iwbYlfnxE7UTXXZ/65X2nk0nVGP0YM8M508wo3
PBEJ7jg6FMN7OEUnUl3wTsgZ/cpzEC4K79SHUqqzcx0R/pi/xCXCAbHwrPLoMlZO
9ovfW9cdP3ExaxsqimHXNnK5hQqfs4iY9unXnlS7PL3ohYxftu3VZhN335wBlYn/
uXfA2RTcl7UuUvNkKc/r2nRPR+CJv4d009g7mXGHUR7tZy/OPO6Sz7rGkkoGWRGW
LmnXRMhOyNr4OX2Kl/4IDL3vOfiqlVFZ3YNTxY+OYVlKGVlpMeg2nIyST66H6srD
CmTVX/xbgIUs6UsJpwXhyr99RWp+jYto5Qf+fg4AkBp3Fur5IGUanHqaCpq2pVzJ
eJKejIvBIe+1LyASwr3vc0ZWE/ajg3Yn7Bc1GB4sQhciNmthp3MHIPerab20Z3OC
BmtuuXMRxT+cJUIRI9XMLJ2Z/dK7aQ20/9YRVGo+usa21lyVdqExP21VGyT7DexX
M9ufIgNegZrpHc0TNUedfPhKjr7VBhvfORmRKkpMOMB44PWo7b+1sFWvrznBo/mq
PlUVv6wySwnwy8N+ca3npx8xCEY9flzOG/yRUOxrYSISs0pBAYGa+CMtD6jUUwhF
pkTuan62eU8QQBoixcghmfLYVvw0K+oCWQCeNiorOiyGJfARNn0oT38mzmeLuYq3
TLdXyLjhLjm4/JqNP9+n5IoEj7i3FfdfFPqak4D3CF+hG21OBafZ4X+x6QbahHYH
d88J9Cl10vkscux03IRGchniaXKoTqGMQKCqLnq0tywIMTwcH6vH0FNb5HTm34PI
rD6xqekrB44ALK9Antye5d47rKIo0VHZP6mrZfFiarCy+TWCESRSlTohPI2ggPF+
EmPm+KDJcIXl9LfK68Zk0/DJYPh2LJS11OsZvPLommj/+Ak8pPlz8KOiDEAeWr8v
fZ1dTfOngnO9mMWh6MU52XmnFP9ZVQf30mch1jLFoBtgn6J5orBhAt7xxyET/TWN
7I/rSOwJpovt7q66TUgHKKvLxiyvJrGNoCEA1o5uWTEFCYvIbYVbxG7eqAZjE1cr
y6M7rkeOOlb71fzi3cTl9DomFvaSWO3p1MD+8uwZt2jLPNy55Ndm9G6m+w/egWes
fTJMl4KimvPLj9I+PutIjK7DQV/+BDfTw2H1dTuGtyGpTSsjY/bMn1w/KGdKcynO
Dr3eAwIR4MxxzgRtB+PjHC9esRG51epWE5wVPJOrVoNKXuM0NiuOkzuHkV7UbIrM
PratFEUX+1JKWEvHJ0HsWUm1nTiC0zR8WwcN0hPAdWnMK38TKQyKGP4opJoJ/Ot0
Xy1PDVbekeftOicAWu+XCvvsMcbCabECpwj/DqGFtL1k5xzu8z4eyR4FH+gUDDmH
1mxmRbFSjt+XzEU3oeztptRdS0rrcGfuBmKy1XLWU/tmdthfGoqHzsSOvO8xHBjS
UgOhBEXQnbaBNlHtrVf8ZeKAlR+LQ5aMvugLfOd9iz2HbH/ktX7Z8733hWo6W1VJ
zCBAWERTNm9yQGfit9TwTqkHrBlrvuc9N60gmXSwd0qakfDMbuUZ7gQfn0U0z9mM
X4m58FTbdOIHm/yRONFShjIMw1PKVPT9ZcpQ1xV808gwqWLxc2PdXsrNsKjKcarl
PtJ6Lx2cShN2eXt/pmyq0oiEDv6YO8qoUUXwPxYyKOy4gMeM2wrRTBfVLs9th5pJ
43kMrnHVEdqB3TXRnGc71Xl3ne+vvwpjCMWXkMJ/fDJqHy25Mu3SCqsBKnX2Sb/a
nQmgNaSZMHWVe0BwBfQLCzKSIvbdddYQEL8m/SaPDjqmwxkUa6GpsLCOcMjpFvlS
XCN7izpl4/Xyx4GumsGTNPPUXeB+86YtzF98nvQUe4fShtUS/JsLjQhufMDLuyct
A5yrhmCh7vXgOjJ6yWUkFX10BZhK05FkLydvb4v1cchRMpS6QzuH1jvdvj0CIIIa
hX6INZZxrtE5ZyFn7hYm7oMYBbSFr29GYjLAx36hcoVwv49OsUPPhmvpavIkh2/W
PXBcDwbsRyDJfvd7KHYwHnISimEq0zVERXS7V4QRvF8zC/sjlmjK0gxWzBJYeA6N
VRroRaZ4lyCAL9Ff9Q9KsmPfsJB8AMkon6EDI6GbV/5gALHv9mGiN51WqqsU6jHm
562hbgu/VHvY7rBtCPVx9YhANfraIr/LdoKZXB9DyJsSekLdDqD44+UtvVg4e+JM
BziOUJ3dyfJVDV5mNIxWzs8C9i6JWFjpnVI6C2VMd/UWJJH9GamgTUNPX1CYs+87
ZUh6e3KIutfiAZNCYI6zhwIb4MaS6w/Tkta/0ILd4G02oX0fV2zjwm/CWhbxPwDr
cSp4ozkIDIxBrTXilUPzBLleoxGTeYXIZl+3khSDIrpIKYCzdOa4jJlAHK8GEET2
Ypdxe/Z8pdyC4Ral/oG2hZmqNQ6SLwMbatKsJNrj35LVwWf5L6XrppxNI0L1yiQT
hswrzZgikTJpajx8eC/cAXWRm75wnyjssbTAVk7kF5Zvrg/N7BFV6MGF6HxbxeP6
7FshOWK5Anymwz+0yrxUh/lpGPes+m3WvyxaQ+GpbZ6hwlPclXmZpHoW27zSLyIW
mYB9TuRwpbdDSw/XhaJaD1eBVaBl3/VLrpBa1rkImaSm6vA7gpIuCgtU9bGy5UXt
hG1SgXehEH07sc337fagpICNsoUL1ub+RbcvkHNS8q0Bxl++FKAfzeO6NyNOded+
FhmxfeNxc+FNs2eI3ULLo+UZX9FYycDAekdohYsIzs2qDajjUj9fPDS7alqZYBcF
vDJmdjdaftC3BAgOv38UjFJmX5oYDgPOZu+DvOB+8QrPduiTX1rUco4HkKxvIk9v
0fCTpCvbkVeSUHEMwanlXmGG+Rs9grERlmZHs97wq9nU+f+VulQIhRz+4zWJqLyf
tdoy8PfPAmE6QSuMu54MKx8BDN8RqsRqZmPsd+9oC9Dpzijd7tLz2d+vv6ivrmdO
jLBcofzHU/FFS/CWiWBquzZTcKS417Yoeybq5IhxvPZ/Vu1YQZwZ2a1e6huk8TpE
PWhWfV7e4SittCSJQ2PG92lASO4eVXJxL6DE/bImQltqgCT6uSDuiVoBRELN8kuJ
taD0NzlrfF6nuK1WxaoPVHd9VX4okSwJFpWQjCynnKBPdhCCwakBg2Zb5S7ucRgX
xUcVBNbaApJLxGcUJ+K+3OCYCLW9sUQPkxEZn9lSWI7GzU4WdtGr7/+gjnNaKKHt
ZmFxQQDEYYeA1PDdeIS6dP+Wo59RxelohYYRzaJ8KHxq7qjZV6vE9Ywe1Xt/uAVO
nHaJ2eHFntOzKTGnWd5urIQsxTP5fQ2FXSFAoBuY4WKR0fK0Gi00Qjk//eOunkq/
RKeC2pB3Kq1uhD06MLER+B2yOhfq8g0K7bU2BPGVRe05t1I7sMgbciZgsHxtyInh
NQo5d06j5YgLs5TCWtY0VIwNXv2INVU/66WNd83dGe8qt38kTOn6z4clJ5SKX3c7
nHMuFnmUn0+eiPEATDikrbYyH2Crl1YSp3agr7XbTSD7Ibll7P1Gh81JFrn1EhO9
fES22MKHEN3qegCaRziV20xjEg9qSGApyLMd10CoCQl1C0GREYvREW/z/KsP+7gS
rFd1OuAWgEAuz/xCh8+E1qdb0QElWqD4WyTsVKkqR2kcvIEGFgOPXHU8eR4tK+K0
U7qIqWp8Q0r2zbXy1/7bQQHh3QhIbtCryHkXfRhJbom7rWcLp6+xbUL7D3aIgXAg
oustUGosiPacwf7/njZFWD797WNT8DgAoP1nGIpT7tN3B/0nKJsRw7KdmpzcIeqA
oBF9v5j9OQDRVQLSxKZPgxMhM07uFIcSs1nEx36GQAIPEBUMCv3o84adGqr4wNkp
nxVYVEmXcbC0MwmXZuMieFOc9DsxOX9xItaB5rhcjOJvQvpjp8Nw1CCU9wM74B+P
YkMEiKOjGxNiCPrFJr0NvEl2QeYHPaIxR3aoJxKKGyiL3kVHLQTPL3Jn7QPrjMoU
3bdRtEB/i9NnZmyN//pgPwLlw5S5GLDUUAOa4/b1Nvd56k9MqRg3kMo4e9tcmB5D
dPfe2B6fltqAqqsCdGwRUyQx5EC3KUgpKhGpEbs/8vzIsIp7BoJgVuUYPDkl+vCr
bPG3Z8pVgBunbcKj9HMXZWgXgwrWaBo3uQwASBokGYLN4gkJNBLrYXH4V/LAyGtZ
xrEN4LbFuB3S2st5SzNP5u5WDn7GhdbAedu7ULQeGm06VswX1IwIptesNW6VH4Lf
Wcfu85uBEFNltzgMlXDQ54XdYVwPwE7LQyppeZjs4InqPp12DH4hh8F29m81s4/U
doRwZ27vFtV2fgPAha3Bs7lKPwJy3iK6MctEvqxE/NM1vM1h9pvfyCElsYzUU9Jq
NOEz+nHx5FVjMSxsyD86SS4qBOZd3LwDV3iPCtWGwM6XAbZXmQM1IReFIshz6GYc
BZUakm8gpiSQyy/vyBt/dOXfbW+U9pKTSI+qOcz3hfFXVEpuMpr8O6DKb/FEcm0b
QhGd/SuciDjWFYZNWiU5XX4Fq2KngeA7Xnt5j6fNCzOvITMb8B+Xp7r4ui8XEmQO
Jt19K93EsXqQCyUVFI4Q4aghH1jA6ahaBfUxon1PNqyfl4Ye5DRGIW9gSE7aFMUv
pAweWV6rcixK74DTom29b7C1lZi/HM3zP/Q4xQxDVmuMhcMIN7jk/+xxHfg0435i
qt2tvno1DiwmVKmUBTro1ah9PRoPYt0EzDu/0nHQewbeqDCyOJHDL4I/Si2MJH6g
Tfh5dUvt+w7j7sSc3lDtvQWbhdeTwE1BrsrbHubxJQSrWe23kcQF7P1/ppMziS9j
BlAvwK01TkReAQx8i/d4x2oj5SB43Lk1u2WtjZm7umVc54p/Pzbx0iKsSKL7ZvG+
IAD91cR61VsSkN4PfKvL+Z5V8F8pkDVPMF+d5yKKBtThXjSJ76U33RLUzoj+/qwM
pr581B/ESpb701TEN1K74NbFHZ8KzE4UYOFIObjJGrYxG7s8G4ls8H996vioMyuZ
l1ylbS1GoMu3Blu0NXN4XdYo5RHxgV0q3NpIby3ZfEmtICtdFct9YFofvPzbSZ3C
EGnyL4QpDNtM8ny8mDWY7RTUTIfE8d7I2OlTPTivZHhNBw73QdOvjnMHNkbaZaNe
hXFckOxsXGWQg8DDfNzUHQ63RgzglN4KHxI2jOpd/mfcDLK/nRM7yv0aMtqJBGPc
2v/26n/0Qq1tpYbkN3vYyI7MrBgQuZtMhj3RFI1WALPxKadMPrhwY8woEwcRXiXG
r8j8IbEyh5zQrsTFB8xu2TqmWczBqXcz+u/+n/SGg647iU5GGx/LBmb7Id0acMU0
FLHvlq8rwC1dg1vmsyg7V9YmpRDqm2Gtgj7/8KPzdDND1fRyGWzNBrrqkdq+FphP
AqyMVVVqQP4ELrZoyr/48Ve+IZwkzpSOPpZy0Vu7zcUNwt9NiQB6w00t6gcUuUWZ
bmuSHG3ABDCjJY4ZorvU73/iEQjCqeLjdwzzBlsqCQBWcbLIGFiDaszRH4rJulj3
3VsA7z9Abesbbn2ndvkOv16LF8tJnEwC1mBs0swJpfxH6FHZcnacYuXxryTgMGyO
56N6HCKNIzlMl1a/7Xj2It4X8y3jnNruyaoZr4PbzNhTm10FZfjO2lgBxFbQ7hDi
GhrxRzMKS1EmGywZk6ENaNfqs1iGMiKowIim/T1/4GvGozFa9ZlLjrftahfHIdaw
tswE5eLPuAD4tm8y+uQVzOrn0hh3bsCSgRNa0lEwHPV5awCanuy1gKFwTgqkOSln
x1Yg+7/PhEe8JdhQDKasa1RB3T/WGWclNuM8aLyG1XTHhJACyMh41FdkoUPbrCbs
EdXpYC4qLGRGYtDjNGNACCoHQUaqRbpgdjM+Us389OPT/HnaJhM1HmpkNpuuZVUp
+DU5jLzsQOeRDVB2k+YuM9rZN5rdVo6fjSirIP2Taf2ozEV1iFg4DHho/HCwA5tc
9BoMecUBKiNCyMq55ZVYXUNtLX7TLJ1AsLo7bVU+0EwU18JtQCSlxVW1ptQEAM+B
2oXusaK5Q8KWrukBfWDSHZj2Md7WZw7ZtplkLh5jL4uv2PRJTaPQXmZewmD3pK4G
aH5khvhz883fNJ/tdj2bwnH05BiSJJN/3QxRJEPI+/gV0YalsHK2VlU4ygqarHHK
Mc2B3NR/tDDKmNOv760ELDHUKyu1QgPzBl7loOhuH2Ky0u0rlYu/t0H7SZyOL4ue
QxSy1GsuZ+iRNzsuYmic0oVC+JWmz0XxLku5V+YnE2RTMwzK+McpiDs1LQJNiZVo
FLGCgsUTCcPO9hEJLKDRa+ihuelTzjMOadJmM7ATBl/rcFFMheCE1dQA7hlYh8EK
SP3Nh1NytF2tfK+hg+zslF8ll82n8fwSMxipRjx6U7rxPRALbjpY4Kik9oVbfAr/
2il43p5hEjrwu8zvTUgtmzzABr79YB8r0X6vb5GYi5gio/gGhqKfZF475zkLABMy
TpWkXa06GWA3zs8vVg2YCjR5dvkT8r+GET/mMWjVp3b59YuxguLwQbhihOn/lY+b
5LA2KH21zWVVU7JNL2YFsksyt7xS78VvCd0gtonaMTpVQLCgK1Cv/tmR7XzgpXpd
P3lGdCVFnIpMSX8UM8adlEfnS3rEgHlxJ1rtYK9DVX5Cgm/OO62YVuDpZJxqe3jA
peBp3lSDhJSK5VSJTv9d2XRlh9XYNKv4nqBsU35l5ckvignUFTEruQGzN2UIQJ6r
4YAQCXS3/VSjyjIAtoap5dKbiH4suEtPA0EqdgKzBzH4pIGAOqfliFzlrYPj3Fio
Jt8c9i8pss8H5514ijT3PoiEuwKSysoE8mIAWzwgEwyYjg1HRMm+GFqVPmBe6aV6
Ky/hfHuc8Ca9brhbxd1XNTJmv4UKFT9LnvqUgk8IHOcvuBL0ETlOKODw2DsaU5Sg
x76/l7hoCiN+rQE9klUBtohFe5eLPlqoUIepRiE4kz5cDoDc9QtzVHO5cfUgQVQp
T86XNqVW0BfLvUrvl0xfO/YmAI4gdjXMpjxmlHYIIwkROVchnnQV4ZO9touiV1Cb
NUylMGGDucZPzcCUkTz9AJKLXFK/fBD8m8cdL+LAsOC0Otv4FyjB3jSMZojatIAZ
8ewiYmho04+MemQgy36qAoV0rs+uH3rFx7VH24wDIRzeRn0BZ5mX9Ps16eXvpbPz
PCBb4MceTw3xqpd7RKBm7N0+aojSnHI6qz4jdloURgioCazNBmS7lvcY625YXL1X
/mVDqWOTdZX6tIyPL+kqUE4lENKSnv/kVEhPe2k0rFg/2bve+CsH8mDGjoNIJSpv
neVa0YmpfkL1RZAEw6hU7cd+lCRkjAIGmYZxbtY8V6+suP7/tGQXZJ528CSWYU7p
+zB67i4rcBc4Je9t25ft8fU/WkZ698e3wd9em+cwICa+FOpXXOzdUQgE4T7mzukJ
bxsMkOFddVwhl54jwoecq+HRdKVScHEAtw0T8O8xS7YH8+3cZN4z7l9DMFBnTTNw
c/ND+GpfdGO9oTKldzkigaKBBgHs2XJSuAyCBPDKiYubMBOIqP3iFT3m6OjZteA3
R8s5hqaCKDw+yKFx02tJSHJxkygTCptzrMjzyORBSOWWzRR/6tFK2sXx0Mrj1tJf
iV4EccEbtBZpu+/HRAlnl2R88EctO+l5xybv48yUEAP+eXptUolLz5nyU1BTsuD9
XO9OYFUBavpT65FTpa6jF25xzsezbXMUR1l9aSbHXu1VJeuChFL4dBiA5t+qHajQ
C2enChNeAhVDSoLqT1eqkmUL0zU4WkrOmvD+XklujI9JRWwksHIWMsy9lG8Ct9Ou
xY/CK18RMMq8aiM2rTLkUKT0ZEVBNeleQCZ74DNkRi6+co49HJqDHcCGVi33NCT2
vNdnI0N2sw5WmUePvSGPxGv0lAH0A8mkuNYw5piUF56wOk+l60lieSg8N0BjJhOl
ims53z2Eqj0Lwau8nRDl5TVyZXm6Zc9rrOe/FIq25kTXn5f4LZYdLwtpgWN6P5Zv
/SF6NY95PJNxqhnMvocdrTZApS6Y0uRZv74NJkW7DrgaOYgLQW/gko7S/3miKH4w
d+R0s3xUqlL0PQQ8CuiqhTzuE/h/eHVfdmdq4L/PMjL10sok8EijWrX3QJ5siISo
U8N74T5oDP1YlzrtqnvIbKkeuXtGqKwdzkpiC9A0HxB6k0jSLFKvYPikbFRe+JuJ
YTmCYpSCc1mijKD0PHP5Y3XC6H/hhLde8ARTCZQDklizlPLmj3DHpBftiL3IMl3D
dvSriVpOM8/xKzLQvkNaAcIFVnHAXIVkvTr2Coo1Tczx3gOuDIOlwXneinwaXtjF
xv03VmXp7fu0bLHFUwdeT96u2RXdieNc7/MyNV/pKwAvF+ajcB0r5jJMYrYJsWjj
Apc+//aStO1PM5bUJD0lpPeQuYJfWe29hTBRX8a0xzkEu6h2DIBO7n0DTPtmRk2a
puL6klrpmRpzAcZk8xJmxGCWPTAeeQc1hDCmJjkxjTh1/46ubjH2UNJV4gp8kXHr
Wq3DVZsffT7E7Xdc9/LE9QUPCfEakYVnbBgE3FtH7qBzDsXba3Qi7kceNeAGg0zt
klO8HKhVJhzG7BEhLGNS2X332hnm0eHBch6pqG5/K2ePZ/JBXdIWUMKaFJEzw5/A
add+Ydxm4GkRxKS3aMlHZWhIA132mrSRIGZaVe0YC3/B4kWoWUHvKf0PVMtElhe8
O78KVx1VuEROlJtaBpXl5ifG2y/EIxUXer0ht/09LPXb3pj2S/d3ApQpTBRg7Kqc
k/h4CWLYgVBXvNX0dxbeb4t9W2kjrCMgc2ZsLgR4fshk0j6o3ThA8xFxZo6S4scc
WfpwkNTCaR5eQEscIgPsHGPMSwafJhIKU/Q+4WDmjLjxqx8uMR1AkYew1EjEem17
RZTC8sHzxQVoTbJWz4CP92DMqjyz4GTmL7z24p3VTVz0XrvpTs7YYxr4qMJmfWdr
M5GiGAVLXuRiLa5AG4Zyq4fvModfFnoCq/uIEFdDAsJ1oM+YL+VPvxPn11vD7PBB
QoHddqy4q1VWfUx50Q0tOtcDCB88I9D1r3BZqbnYcAbwjzbsbnpxUILSr72cDZns
+iSTfAE6MjQhmGxbNPHQn1mjibx4wk+zX1mHOUMMuLDR3C/Hi8ln4OvkbTG+mEXg
U0WGo4nBvYR7bR6vi3HMc9+Kh2F0Rz164ePrJLMPUREjxYWOQU+KuEokOupN9CMJ
67MtJyuBBPjTO3QDhd+zHUQiz+M+fMHR/ZxrI9CPFWE78LkbMQ21yqfBooJEtBPj
8aD1NrHtzsSq24uAYHt68HOFVlRs7NuKzpNA++u1v7/rFJ8oLn1bDBoYhdKAJUv1
paQBMTpzwDx1KUzu/n8yrS475V9B9Y6rBGeYeNYGtPUqjNxPyrat5Ah2VrSyITnA
bnPSr225ZDEbOxqYak82h06PtfaFmIqy+ckvkVRp73EdRGqgX57YqBxmcqQRtOYe
xqFBl9J+VbupP+LSLxsj9C7KjU2UOPxttjxnX1sVFaBngMQxQ8HTP6VYyZbwm4pE
9ImVIve/hp+YC8WhlCp4TCz81WnNgyCFKYEFELOBWhwyKxY+Pbx2CkODqCyeXv7s
RNaHpU04k6IzYhQIe1bhKxelJ5DQT4W+7oy5LHqQnrWihXIod59wi6EHfJpykpIF
25wkii2HAkzamxyq/B5AlELKgU0WcULFuOZL2iT92eR805Yxo/U0XloRlPKA8xEh
790D1tFjmlkT4R/D1IdWMojGjDz627fXF6IRGuUZq5w8ikoehW5kwOftp0x9kJhJ
bWk5mZSqd5xH1Ijs0IfWZ2lBPGkXfamJSmnf5b67Hm9TGl9aUuASCNNDmZSpuiRQ
TEfsYS6COBEUZA7kt7Ct8zUM9cZtpz8GvjoffmA2TgsA44DFJSRkI1zi5ByF96SL
IyWlaUi5rmhS0YvVqgrFYtnDfyHmSJS9pXozP1TnFRlZJEzumKLqZ6T/T1JZ7KGP
cP6XouVK0smHQ8jFt8v7hJGGnmUOguVmyytjniXrxrHY+DEQ3hjsA6ybshwnUgiv
tSpmlFB9tBtlvHMXGR7DsRsQ+L2iUet/4syRxv8I2GydOV4F1x1QKm83PNqAj9fU
hlVwWUzoWaBml+8nmC13Z7IubX9O7VxZdj7dBPvLRzG4Y8VGJPcdCJeodRM2IqbO
Pau9lDN8Wy2rWGCJ41iLKNHMLZxjqzFb9MI0pII9u45bzAubd3Zef+/7Ld+K8uF9
MGqIsBaVPMb2EjKJmzQ96fhqOX+72PUKLSofSW5MEmVhWA/onmeqmlkaxqNEERm9
gdbIqT39olW32KYicig7f5RTBfSgQk+nMyMcqcrWwUhQ2gO7ANlk2Avwo9lgKNo4
q114aI37JCLBSLwhK7rGsUBM1Wv6FefJ7b8rkRlZx5oxIFHcNZDNh7/iFOUs1Z2h
kzzu1BXk5rkDU7p3XVfgJuVC5av2cYLPgxLg5FD7QqBu6meyCA7WS5Ku8u9MErt9
mtJA8bVZN8RgYzKWhyygBeJvnbMR9UjMzRei5DBbgqK+91Fa+Ftg8B9/3mvj9Xex
9SQUxPj7Lyq5T2lU8MfhbR92SH3iTHEaeEtrFgel/eYdTB5wCTFD9XHyP8gR/oL6
XXXXbcDRX2uKmmeD++ULCSXhw18wjnIm0tekGjTmKF0tLuFE9LYmRzNLgFlIL9eZ
cK/oxzK2gYRRAqlyojZFXI6iKMab2uSXaE2WIaTvXd4JVgk1GrxrwPRgW7FSkV6U
qJu1FntO2gc68IPUQFepM/Ch16Bmpqq4j1pniBC+u8L7g+def5+gyWq55uHQEPrU
tFC9VxIMgsYvo3g33lNpZjQBDPWooQ9k/xwPifTKPxs/7gPRkBKasM0d2pnURBV3
4oJ4rsOpCQXDjZsLKgVrb6/B0h4r+tOMCfo+pNMvCwROoxraIgm5qTkUWpoFbN5P
cQe44XNW+fHVshulD9RgaAiLDSZ0iRb41LK2fggU0X+NDI/mEN1d8RvRB/pfBS26
t1mjx9OmC9FBjrloG5Z3Yj5zoPI01+JMVOdzAAXaNk4dI22Qtk85O5KLRSQS2Vpm
iNNfUEpj6dQ4YzJtlPcTs/UkuUcMGXDHFJlQ/h6Oj2mx2yXF6UTMHS0UXfasNkbC
4pjA+m6KhwtX66ipOwdND9xyUgfMHgcRaKlRd42jWBiR2GiFADziP+qhHU99zitn
7KcGFQSgVplHQRsxWI6vB9LwVuL3DrRpTqXL2r6Di5aDDRpG+HbPETvQEh1XhFYm
QNVvRfhIHRbErjfaaY/vK/SVqOx92Ehc1AiaRHbmHOuAyrRYd/W4V5DTbYnYHLOe
Jk5ZzFxsqAf0xuDC1XuSA0bSyTn66xJkrOstwZRKTuroScCSk/gm/MTjg/OWJKJJ
RKlSSOWPX5uJTUSWFL95Rx25fL6Q7YdxTB+6o3Ta5+fTSGPIJQAvIkoQSFHGk81r
y/1VL31anxYAkw9H0ry53640r+4xPfdMJupWktrsF/9oZWs2AIpAAlwWdS0/E38b
Lcd9tVHbSGJjZtJojqrqMnMklmJ7s1Z8awN3/4ENESp+Hum8LpvuVruEUvR33Snc
ibCd9H+NSfgD7CDOBFCQNLHSnKLDy8dg7n//mc03SzZS2B+QkYu3exyq37Axoljm
GwKKZNCjmfbbegfkb9JcyEtQvCb/3Q/NXrgLsJSkTnrcmYsmeuNoO293dhzgR23D
6ow0X6im7UzD9mYyDHgoFkRMmmpq5SRjsxdgThmB8mjLtHwO4NB/A4TRwcPt2cqq
EL1pS8M1AFLRi7ucoA6KJrwsn+u49yBkeAPashQkRhMkoSEdkPRiVj0AxkkLyKdb
fKJS+Xn8ZyhrCpAh3vu5Z2Szgos7f075MV/Z0RTTZ2t0Allc6sF5b0lb6gZJMKxu
CVcVIL+VbUN2aB7noc2eQ9ryk11Nw77X+flA6Rnwxp51NxhSgIUKS6cAEvnFt1pp
Kh2l1Ep8cpoWdQ1AblptbYHOtrg13CwhTf4bvaoLFjUVN4PhbLj13AxfynvqMLFF
O8KXfmBAwiLze8cX6hikxijetgUv3roEVE/iFbEO+zbBUYwVfqrlpbHcu0MCSb5/
BqBcKx/oYJFhXi8WLN6yAKxs4U8I+1ciIlGUmtr84xqwvSWBfASeyy5OEt9tdzbA
myl7CsER2RbFbD5LoyKv79TFRRe0jTmTUIvgPv0jw878E9iNsKgPHQCTFFXob5K9
xbXoRid6L/ojmXSmANQqAQUyOkyfmNQlZBYJsHpP07BsLkehfCh9D1fwPMvaLJSB
sFgruuTWqj+Le8FzkFC2Ry9QDRJYdxwgZRybKrWXdDbNr6VSJY8iFPtISD+4xZi4
l5YQXmCNpX0J9dsaMTBLjifV8V7rs8pCuZSOaEgn6shHu6ARkMkCLgNHJPDaYTNO
JDAFug6wQW0zFdb1y1tSdtEmkEKfz+qtJNloKuRRihiW33BjxnH4UFcF6pq/8cpv
Z8HzqBE9p8v5l4IZGArZCAT/yQlObJdV9ncg4TZvjycYurn6OOzLkEApmE73vm1G
A0K8heb1aQHRIajYQTHhG0XZcmd1LUDJ0ijnUeOi6xD2s9F1vNPTYb5iGH6l7lQk
vJOI5yfDwjXQngVNZ+ieydVyi34xECScyiquFu2InZLU5ndkPUq53nTr+cE7hoU7
1Rig16VoA/XFaNLhYod2mCXwJkLB0s7H7U2eReubBEkLB9tpL4Wj0IVd/PjiAKXb
Km19EcvJB9zJW4LmDhye9P9qW/Pk90tOF8Z0TROIiLAilBBPZ8eVLxTwO5kLb8qc
1E+4CxB0elgt+/Ub8jxbCjH5iA8O1TC2LbZdv6J7TUvoSwux+gmri4Pj1oKLCDaK
Q8C3VK8rkIJIzDovK1shhfUxA1O2NT9baTs0zs1ilDB5DNDiMrWo6PceMNkLV4Ze
tYULR+zeP1cKZAujjKJCMJufYH8VUgawNC4Iesa45UcgRrzEW3JqhQzHzMkgy8lF
W27ny3oB1oa+rFtxDEPSt3PeYbvbPryK+BecLQQZI4b13AZ3uCNKZirU2FITTNS5
SbICww5xRh5Ns0k4noSRY7It5KFfhkVYz55YGUJmXfa/ag9AYsi5hc8myUSyiWwo
WY5ZHyGaepPRnVKwXw21RcGnIvrJOYjX29EMMSlhuuW8+q5hBJn+bIxb21z8gUtI
bq9i4OrHkPxU7vN3fE3w05+Sx5wdNcIK84HNVYgAtYCg5myTFF1PIyMCCa5gGMSn
23gccjkw+u6GYTP1q4vVqN7HLG5NBAZE3ocliUXprbMBN4JBj3uH6WAGRSb4w/DJ
QkspfzL7XerUeeSfT+hNVRFmgzQGyeY2/g679Z/iPYH8G0Ld1OO26cFaVg3PPsnX
iO2TyByGWdthNPhFEd7KJGtiYHAZoHFKJ9SJyo+5iju56gwPkoJleMDZkSFCxcIe
0snzfmgQtvplxOyehUD1PJ1CjjPrA3R0OXGNArh1cMJmTCPQQsAwxuuTJFtuoWZf
iyailmB2VO0yll64YnurQAIX4reUAeCMpDDjKY0yrNl6Vk6VsBQJI4WwuUXc7cEN
IMGLZts45tCAGLoeUlotCUAIxBAMOgoCCIMLxXwf8vBP2Fc7QPGfXGwwDKbHcZCa
pVLzKPt1TUNh1DieO1dTpU6gxGwMRJio7yItqqH7nr/UiYXaQU5s8N/1dEYiYUVK
ucHGt1cdTzUYRJXZfHzZfXaogNKvZMpNdV+UQ0EXWqahgEUlVXOiSxbobWPDPPc4
kEnBioLsrqfMf1LVfHqCIYnM08aVX3AUyZkGxrffgYYlZ6hapCjNdGSnWm36kv/M
oMEYGrWupuriBwUfMubh/L4DpyUsao+qERWxFFx3gY2q5eBqBWceVLX6eCGU4S/J
sBN625OwNDw4pSCFB8FcAErACJF8qN6crlFze1Dgoeq9dP0rm6O4uRmKKZfiVeeq
FSwTucRCWPnjquLG7RjYPHekOICMgwaA0blIXtuTUsqHUavY42H+0dfwjPWZVdJ5
r6D2IMYQczMToSXxicJaxAaErqXQYE3ijQH0hm8DEiJg69CImgzx9BQduHOURs2n
zSIfPumTgbrt37qgYph7/eTqGdJrBHFkpEPm5YdNB0tUw+dk2KmGIQNIiVPNMpMo
YoE25DhLtm/BQ1E5IMza/3lUcx6JoA5y5mHeOVW10De0Cso+THioZ2do4iK6UEC2
7Uib/62yveL92bilU81apfaauN/r0WrXFmWSa33oTKGPFhnBbw7nr9ERpry+zRzr
KJd/ineDIxcv9kiZiOluSIuXnZTOikPeV+9bcnjUxV0SpMU4kY6xruMmG7pfz9qE
rwvyjBS3C0yTWkRsAffWVMloVLXITFP7ogqj4bZljPvFAY1ileKeeNuoLg1RI4N3
SNk8QjSaXqQbA3r5LpgCpvRiFXvGzSaPFEOFtrJINjg0HRs2QthRXFYqIu1+rilA
+vIDu9LZtgJ9g5inXAnwyM8r8z89QfJFXSUo0a7rh52B9GG8gKqTZ/k8scrDf9JV
0ROBQVUpSc71xauzjw1MpDSYEQfXcxJY4dxLpWEeT6uS5NZJe0ag5vLQUUXRO6yZ
d92e1jwOAV+uV9ML78ETLtSQVOeuBQI6TmZG+4izeJ77qikUXwEe4DNyPEey1xbd
IAcoXuRbZZKMXxOdGSWL1OQdoGk7Qh4TShS/xImq+qmSP4YBDiuHB38d6cKi/kLE
BZfYOY2EiB8MhR9aBVULbjG31s8rYglyCQiNm0DFU0fzaxsHaATSFvH9a2RNKSKd
/OiIDEEh/SEq+ucGJcj3ItPL5FSquCzaX/RZ1aYuXP0a/mznKnJ6S+fIYtbe5B1k
MgqjkBTKH47txOpmWJ84hYD9oL+DZHlCyXdAz1xRi+1UV/UO4dBLOo+kcQblU7y5
lWFFnDV29vPA2S1TZpZrpB8doI/Ct4vUtq3+TY2U755cVCuhjEkEtR294iIFKRzC
Uxh80QgfBptqh/rhhMxrGxI/P7DZLnZCxa7NeBWZzCxI71JGoX3RMLcb/RpW8DFb
v3Nvo22sMCdB3kVaBNOdtxNRZzHay3Wlqu9gZ584zz+tYBRKByFSdCATjU/3J2kc
Ak1pDK1OzST7WTxfarGP2xu+EhogOK2bZgP0JTE+hq46i6MQ/Zqr1KeDujaAKeeZ
Vryo0ESIrpsGOCaTDsJhTvjVxEiFaZdwuiK6rHNy7WYoc6Hr3vo02Y9unOhHOzvs
ItIBQ6yCI0JzGPfR4f06LH9U+cfmw/N09xB97vO/2mm1IRmPn7suvPUeWgE8LH6G
4yHSrszhRMdbY6vNbyDmqrM8zt/r8CNPaBSn705BH48OGSLNwYXnfaMavm35cFPJ
eHvZkdReO2r9RG/UtXd5BGvEO8tGfrUX7ImmAav623XAaySXb4maTLs90Ein+Te6
aHFc59eAYiEQ3E9CAG3zVc3k5FPP2556eSogR8omHn6ZOMOt+YpaAeH1hF2sEhEF
LXehbmzL4Xmp6F1adXa7iFHaoPFtpqQipg/yT2Z3XkgrZxWqtSHWcGzyECOVcmZr
zYeADw1myY4HhmF3gU7blby3H/4R7RJze5MvBdMj6RoQbaCwMskcVX/7WRDIjO21
6niJZsIKH7i/x00wFvEwHmih6nQafr6XIwCh1KWBW967bNAhv6iji38wg5d/ZNUk
cTGFX7+KghsTcvWHCYwV9balxtncLbUOnAd+27dwo0dWRsGNoBfUnV1Jl1Qq588v
Hm4+QSTP8t9ujjStmqd/wnzLybi2AVKfYYud1UKzKJr+ZyXHPZSv0LG6EfItlWDz
f5McVrw5oybBcXBn92c6wSdFZuIlH9kIuSWDZ1K+5guWzofBSXA5TIL0+joELS8e
CW+YPwwMlvoNT5rqDCYm1/dfhNr3T7uSORQe9jAUv7azWoo+ED9pI81xHUIQRMGg
5zisWOdLG8IlzVuaTXOjJ+lS6u9aM5BMMeYq5T/s3Iso7h8vHS3o6lI9sdrRvwTO
8YUKxr0JGeGpwZ5kuMWA+DX8bm7cZlETqt4aanULfjK21hV1gUdqLiTqAiEnuqIn
vdrRt4SrC8hljWe7r/ldWoqXxqUsqqoegiTvX3KTvitNSUjh/xW9INiwBNSEi2Uy
cobFgYLYt7hiYZJculEpQosQNZtGayKn47fUcxMItMGAojXIhh67hyAK7gtlnsVJ
mHy69hjBmMj0U61L2AG9ZB7rNIFW8KiN5MRIQCTFN5thzxyjU8gA8PJ/iySPCIJX
Y/G80vBrS5DEjOx1aJXr10PYBs/J7sGJJ7XtF7m7N1+ztwNPqvIaZBI7+xMPDS7V
3p8w5JR+GuT3FnfLkNswGct2fum3ym0wvxHWL0t2DVK+LH5UAYcMKPw5oKaTfM2c
qteqbs1XOpUpgQFE4+C60PnOO0GlU5WFantDC7HjYC+w4baAuwfYaTixBDgp/O6a
yy5cOHJFd/caeuilQ5uHNfVg9VmElACMLqTVuvGF6jscOXXjZZi0srnnDt8FFFBG
/byYLJmMlbCCXcpt+EWD9dCYq7XULZ4SVGDbRAoZngFkJw9VRDy6Fx81FcUuk8PC
7KES79S/e88MHMRuVqH2mpsGqmRdu1nWIaJKUUt8lkq0ZRzu+E5wvcHISpkdI17O
0OzV35n/O/IDJnkxRWYt2sDl725Sm6WuMM5cp9YPRIf5QUSV75z/Ensy7VBT2wfa
QF7mvHlkkAPf5aALb42ctElzP4huf4O+DWx4hSwXB47BzFtzrR2lv8uuXOieqbUS
BspQ7Afd8NgVD/kkOPa4OPaYfdr3qaowGIjsynIWl1kiEPfPsk0lbtpdnkZt358r
h76NY0kWYXViGFCxtQ6e7n3h0CXSz4xV9l9Q9SrQLvy4RC4jTAx5mz8Mj8/plHiC
vQ1PvYtAqVLh7jwB7Lh+SoZwxe1Z5AVvT1SAAvUO7k63GWf83zw+giJ+PsKyw4nK
WmfqyS31e8paE/upJZUDFaDLsTsBVPzREUu0wC+M0TImjdL5jslWn+8MUDE1rp2a
q7ZKWtB6GM92+PblTN7N3P68FS94VGU00IcpXEUWI1R3Ir5NY0+727do2kjTG2jo
Ia8jrTAHHCXAxTGA1r6bLSj45ERm8HAZCkHYVLSrDmrFp7OmshBiGycnCgvfnbLu
LBCfccn24/N+u6lnBfqY8SY9salW4vUuo3rssmeOgxpX3135W8mRaVHzoMVCYajn
6drTwBrVBrA5FZS/1q8K9EfA7Amr4F+DZ+2lO45UX3w31J4BeanOM1N3L36F6sZ8
Zqq1dwSvIAvAkwIKolfhWqGeQn0eD17JNHrW3Dprv9dCWvTSjUD9G5AZWWdgtHoR
v4OdcEZC6fosX/rKriqN0EwpZRN9YG7qLybvnYfNtUdES2BQUc7sqNxgSC8sp6wf
CEuCTp0Rn97YOty/0ZdvMHYofEqGMauJMxlnsq0efozrYSueEb5MiYHsW8O0Vkwp
7osJBibbMwFE2cffPwDL0WI0TA/IS22LBGBKHw92v2RF99RVCbXQ30kH1syzAYZ3
nJCa/4s+ixrREjF0r3mgqkUTlKyjfQl47RUgWyFwq/KicUNNhSs/J5RzpiITfhC9
5p/V9qh4lAdLzTmUpsAlNvO5IgBSiabWRuQiDzDV8ZkKgciQ/eNQranFLVGSzH58
9O3+fDct02RqDfMiDW/Xi+eVLyaS3wtffzCQXdrki05Gm6aSFXEdYD3NqvYHUqFI
tMuRvbKcNQr6f58/Nx9guKw2/I47Mti0keemPvAI5mj+kutziouT/jflHnIySPfn
e7d8xYJHcvfYgX+NRan8r+e25T3aA16+fJN0hSCknoORJdghMAT/dFqg+f4fxGAU
H/woe7+ufBYSTaeX5c4Oaw9XG2oHyTNAdOXOp/tID+u43/F7A7qW7JVsJj1YYJuE
gduVKUQWETDuMlScs+K0YS8/JIfRv1I1zxw5AznED7WU4/fhorKg9Ckskj4J+8IB
oX86vz3FkYoEZ8mtBT333aQBFVt7W3Rh20iXa7ACEbLBMfcee5gYdDFgW51DbByf
VtSUC4NSmiet+CXfObJmI3U/DpJK/W7pOTGOwkNtAD6wo19Znz95JArDL1CMrYBg
z6+2m7y5Z7DbrSQoSbnCdWmlgZNDNoefVzwOMugqnpb1cPTI/PJU1OQnmZnj5tU8
Zikp7eMmDiqc5DP3Pxn7DrnZyERd96p0K42mhGfR2NBMGcJOh8Lf3u/nvC7OOQcB
VaIXholE35N6WBz944w9+isDxGeG2bttfE8Od43jq9HjIcXpl7tn3GPR4k9EUTi4
9BKCQVVWtxYUFEwd0x9NB+3WP2Yhb4Z7aWB481r4mV7Eoq3UqPZnidI/YuUhiauG
R+PaZn/0G5raWaUGBJ5yrR0w4vEgnnJmMtqZDPWe33d8mJxw/dn8WiFMeFmxln3Z
eJ3CIWdPdmkms5CVoc/6P0O648MpLc1nSdOv1bPKJuc4yg5EIyJOP4S+31to9z3x
yFYAFrC4bTdQeha806Zik9GZ5muhdeWtuX4u+4q6iz9gsUjf3iqeXyS8KPlVXxuS
5fNGGIXS9VFmloaC8JMFEdd5mFhT5xO1nXdqHyLzAexoTP0d8H0jNCEnf+p5jEtD
bZ2AOlMuhMuEpRdcnbTb8TB/pMQLmHq7v+iApvXdjg+tV4mvD5O7uhu8Gf4t3hSV
whtG+PuoQHTo6dZKI1jzkqm4XKyge/UO0eCJzJcQcKqg6RFYcDvPzjrNazePXFcB
Dcozkvwr1lIrRNklit2VN7BHF1MK4jiwIiVHAmCXMOA3bkGd4OL0ONSRYSwQBotg
W4F9Wp8v/fTOWR574hVohU8ZiBH3Iw8+IDiA4LX0Mo3Vsx4Uf2hmcqWbx5ryVI77
zMih4/tgW+64ktHzhu/CVZ8OaA9khq5uQFfBYPw+l/gZsR2GgRt2r+owizbAJm0/
mBtdWW8+KnBQGYkqmEFOH9hfzHxnzP8LnF7yLBSplJSZz0VBbmz3FgStm4wppaov
Bgmn8239YNNDCDOBelzGMq6a7025CfjN+XjibeksVf4dsTBWhftx1w6n6tT3bWp0
/s6wPl/Y3VS2RB/X6a5AYpl0Gesg5742Ky9993TsCK9QTo1ZxcBhX6+smA74V25f
3e0GO5AIphQcVPABq8Q/CM/lQpXRJPP+PQO+gKdHycD1X6xx7713tKZP9ElGxbsU
RC/iHjWKi/WldfAbFP7+qRHwhIjL/dTghtKUriV4DpgZICk0vXTh2qd45o+s6RlV
5twq4PhyOo93eKXRQWO7CC6sGT4AVqZl/1ZZBm4rkY/+Mj3xm2aUrHYyhYSJEkja
iUJT80dNPuGduxaBXICpHxjfHHbGOlKCshfAM4CB8UTSCPoEvbKGt8Op05EX/FKY
HWMXikLiQv4XFdt2U5Laxe5Y1hHZj+28gbgETPDzuEizzjXTq+2/Z+5COFVwSjbu
OJRSRwX3u5NG7LO3oxTnQt10sSzCahs0PMJXLza3Ze1gO+mda73r+IuvRXJRu16e
QSzXwkEyUtGkaC4PQApp51T1ugaSJNebPEyIdTkI+YMP1lLWE9qhuoWdcwXLl71Z
bWbnyfwAFDzuB3hNoyV0lt90Ltr0xGy2Qh7be8x0b/ztCsOjaNzG7Vt7GdklM3Yd
kHWKAzQ1zc20o51GTdUVwqxBYd2i6xUOamquH1oFox4X0qi+Yh+G1f7BgMl4UVli
KBHh8GlM5dlfs1Z86+HTr35tGbX6V4E3y5wmuVgZ5RMZanaKUJOBzx7SBcgYDJS4
GsMDNPxaEI0xVVfTrvaGUn9VwMrHHuI26GfZ/rA1XMjIRxskRl9Ncqk9pG9IycYI
Pz8EMdKKciBlJQoYXMoOBQM97BzI9eAbDARmXvI8atRoRZMRV8rZtkZI7sc55ouo
HOrJXCS/Ughd3gcCSScIyz6n6yAmPYwLmFjAE4IAUyXFq+USn4GZzgdwKvHvXg5A
cdpCM15Fr6n2FY2uHc7ECR3ztLcZZrP9R9mGKoqQlEulOu5q86vbgrCTVJkdFtPb
1bX5a0AHj0JLxasLoUbIAOU40sE6bMaoyNYawyioGTVgy4NEeUI2C/WK/9BtgBTP
STZoy9KTNAoIhmlU+zfwY0RX6uUlmjb7X0+HQn+JQnxPCFLAf/MbfIHal2Z2dxu4
DFsPari9byhdNKrIDKkEeidOYMB3jwRwMQkxr2cJsNRbLAgDC8NF6xIErVoa+9qJ
D5GT95of7uzYHgbvFPKqGEPBkhAnVYxu/yt+gnbfOpRnHbdJmGIBLBtABIQDOdTf
v/vQvMqhW6s5aWRH9v70QiwPVtHIm5thk7a7eVk7eEop1coFrxHeJTdA6epidKVM
azfeCF5/+YUkbLzeB/wuOTm4ex07eBvQbS5KQcvl1j9fO3gkE1X4KmCFWUpB2ciF
xKcD/7v55btjSSbT/9WE9hYwKZkBymkc9cylDN3h5pu2w7MtygFvd9MoUlrjDHFO
0CeGOtrBR+85a6Jl+PdbCs88ED6H3Uikek/c1Jew09QXXr3oyOOr0zzolH+BPAC6
kTXQoUo/xr80GGbDoO7l/nwXT0/BNHfbPrIJzOegUkjZ2xrjitszC35L/hzOFc74
XzgSe1v9yrCxDBOmM8YLLYgomrTQ5BTACMM0TJc8rufpPaVAl8YF8Vspv2HbZOxm
EMMkvW1ndyved0UJEnWcCcS8YCtXLZ+morOzRuUrlorIli7/oNYqN/5RXSc0JEPf
iKMNmw+GLzAYF2BNaHbHy/eXOklpcx/EepDX13EKD1doQ49m0lm1ErSPJpcaV+XT
N5XPKrLVm7A9cevqoxYL9USHWz6rDHZdjWt+f0KAMbS3s47Q+TPVmsiNJpoJ7nI3
sZq2KRJ+OxdsbIJCJrTtZcmyQPOmp4TFxy5YTREwjMYXSEhmxZxxN3CV/d7ViQDR
6SKyjDwynAO+0eglKUWbdwTOY1mL0KNIBSOm2K8IZWqek1cyGGNP75UIRCj+CsAF
kksZhRm+gZM6lmscnTo0YaD709iZE9QMjHUWDijYRMgnk+qbBemwvKcebKDlNICN
s+52SQcl3xuPtHCIcrY9kbtg2H28RoRAE/aqi8hc51IqR/rbR8/7kBwq9VYWCOHr
fc56hpby3W7g7VyVWYt0dpNw63VswCQqteoX9SXzR95R47ZQpPnlVuL3os+n6WtG
Eh1t36l1BxIZPVtYKjhzOXi5wpC3XGr2G59Lk0lGzUu0v+pdrfN2jDpPxhC8WOF1
z788fd23aYFFMf33Ob/JXvWV8bn5XUO4L4nbnLGOOH7azt1liuHY92HKu6Tk6YAT
4UYMmh86rI62jaUo8txD8fxg/t4HW2iU8ye8eUXpRI3dBzqbLZzrvkUNPVAaHrzK
sjGuEJU3XGjCn8NWHwyqoBUiz1qLOXWU2XrTwxsiFU8/+RFEhDAkc5zc/ATgfd9F
iM93g9tYMM1jxGoor+q6vpPiTyp2qnwfEd72a1qkAS+A1VAdcB/DQJW+aPNRO11C
NCddAb3eq0+EE2n+28oWs0gnl0Qx7jRqOqDzv22CLxgga76fLQK3f2OF4LvtAGDV
VY2j0TEZA4JhcrpxpGQ4htZOBjv0awncjJbtkssK522LuRgfl47w/buW7w8+fwir
ZHWue4jEB0LVGgKYGxSkpN4GzmTyZT42AAX65YS+GNMfS4m/nlad5DwDe1NVHmn2
5IDrt6O/XfzhmzVCLrmXF79uthXkWOkh0yMCLXzNZsyJtuNDOjrIPemgZEc5KQNr
rnt4g5s2iX2nYQMgojeC0whAj6Mu9W0QxJaZ5ewQYEVjggZO1NtfR88qKsjQ5twA
T1YjtO56hul+wcvj2o2OwAkyeI0VI1oMBty2ajEuRR73TX467ZLA8KLEV2Jde3Y1
4Z05tn4OxMpvjmxjJL1haupLu2rFXawXyZzXeWC3J1cXhKhO+uSG5Uc5q+4VLXZA
ksnbi7x23uoaESBYlDG2Qhko88O9Swlq6SLL743NFE+uFvILVCSCWHsLcZrYsNeD
9c5EhRIvUgKMU5g9DSbVjNjLzu1o5tcNGuSyJ9JorZFGn7C9F7fm/z2VYeYHf6Ip
t3AQ1vCNqdjYUdKtykVigg6i+r03veMI6jphdw+vV84fPEW133KKkbAYFy6Dwi87
eReGr4aidWiRjC0bzz3yyDxuXHZ9S0qtY4XwRY4D/dprqtM86MHmIxNLx0nMNMbM
0VV7XL2Wruz+KLLrXn4Xa/mHAfYvzLnaPfWDRoKqp5vPuTkWfoI+C3IRsWO7qq2F
9/ELNMyeRqc5a1GURZK7tw6kAdBkfFwq46HjdG4LBi0Y9yoCKI45vu4UV9pj23WB
Xoh8ypmUtrFVtxVqAvR6THWe+qArRtbn36Cawq6H6VaKYhKfvD94qAFN1NFwuto3
K9IkR1K0Au1n1tz+98JOnYcIrixZ01m0IeziNV++jbLJMowVQ1VXPk+LqHqKJmIJ
lZ8PzgDYaEN6y3mI523f+/KFsMii0LenmgYlS4XIOTipGYgZDfVHdScswKoyk669
DpX20jliE+QCpzuXeX9fm21X4Dg9KgCDnBs6t26INtqaXcgxRnbZJH4w0LYeultX
7cb7HhxHbuEj0lTPjhpLzCk6BsJr3z/dQGLmjAFZBe6Bi3vCsKNCLZ/X2w441L5m
T4HvWT4Ea6T8ZE3wem+bFRpfcV6zmQl8tkj6THaxDXbbu7C7oKMzYLhvIHr0kOso
/NwDIYomLFXEijYdhTxFk/gEXK/1jPAJ5GV0WpPELK3UzhA/SjXFX35Lf/1EzatX
GpUseJgR2t7Kdf6mjnpUlK3OFoxNMkWmcP8FR1hoS8D1YidwRUme4g/i1UqNtxdr
NmZ1zUIuq2hyKuLdyEhAXhsY2saCuWE9YA33qWaQPPvJpa+1KBU9NMo7PCzWejw9
n6IJrlMjKD4OzOUrP5HHHPGmPmlom4ovexlR6fVOw0tcpONCEV5xH1a1gUS1TwxC
jrx0DbEQZVExOQYJsZzEnA0q+9CPzury6JpGuW+BVyzds3FWOy1ukzzhg8D8Bebl
8XICGYPsJr7hdcJGDm/qbMFkwSCKTKNamSrWid9Astg7h5SPWLlbwqj1VthDH+tY
h2IYTeHwxMVvh/wqJiNnIB3Qn5LR2Z/vO3ecIAY/wBDxGNM8FzxH6zPfLbB8EnzL
wccDvSaXVD0jUB3asMl9v4yyuInOkaug3Hv8lv30ksVJ6xowzYHw+7Iwty2k/vMU
F6BwodLyc2lFtfyaruXGIrODflStbQdJ9486yzcHkW2DrwmNf3oY8XP3fqMYraZJ
osGxXDfb6BKWXmEBXQU4dhVw3sDTyGOH4hWOuSHfrtdwdVhjnm4sCRxFOGuxWx+y
33+ipPYfRJnMabzOjUXELwl8B+P+jm+IkW8BNHiKJsEzwd3EwQXWCMhdEBQhAfiY
92Jflw83ppUwQYxtkTyYv1ttalZCF4Ewu5Auanfe40BesIO9o1A2Wud/+1hTJQcz
1XEGSgPSb9HLOH1LtWs09fZiw6WXITg8mwWm2rM6FqWTtglnF2CNrPRpxbChFyfm
v5FuEEW6wloLw7XMOU4ibvjNwQLPTOeosRYCXmXzsCbiDKYCA382j1oxoespo1dc
65ZJ2rIqR+mVAZcjkdChkOiEuAJF9XfACUK2BIgLZ1GGmLlNVSnoG3PFst8J9RsI
L+wk1OpfeDeC1hm7uRwb/BXmyTrSHy9H2Dyi1fkoau7u1MO1KA0hV+9Fk9xxFZIF
wZqJPWgafo8oovlgfpE1rwJh+FKpimPyxq9y+gYDBsm5uY5Jeavp4XBOiGVhFLj2
OdPkvJ3PCpnRM9zUmRIwilJi3Bj0InSo4Wi6WjeGuFVtENt4QwuQOtTQQ0/kYPOQ
5q0Pn2AehNdoR7+JROS315Fek8NpBUmh+wXi0MxgPQ86v2pTvVlw6rUnGd+cvTs6
v7KL6Yf/dFzR5+3R0uZiFmV1HV7kjVZk0NGICbrUmJsblz8hZQtBFTxp/59su6Cy
/a7mwnHIVI42oZZ20EcFeU4/4zRTVvNYfs9liL12NPQEgPxd4g+ZEPqVQDv+wxYg
eVRL/BhMKtO7W0Io21xW4pqkRZ6jKGgLulhNuU8kVUho6jRH9Ft7tocMMAeYqVYu
yH2PdnUEtvZZNiEHrmjw8OxcYiIQHmxQA0e/n1rDjMA4ikUkgHF4V7l3vpz4Blzn
o+HHr9zOiAPGRcgPUm0y/RMj4H9h/s5Zh8kyNq0xDWpc3ULa7Ajm2+HIobUzXYR1
YUX7l7UYbL3WeNimfJ65PVBSkD+LBOQHHI7WnyuIYTMrGycHxHROFuirtl0XuvCd
P6bBmAUCf+ZVg5hBJAWsQSEshpL7iPLuBbQTeG9E439vCbQFiHhPvrrb2wuw8TRv
LyKfjFm84BgH5eaMMvBmMr06YffycY/hSWJghlZPdNvj8eU3p+pwh+CBm8GySlRn
ipYngBPc5OqE5xHaK85W0uPmVKDoitZbzEeF2litesDMMDhViLELUz6Gs2cegf7p
NvBRSoO7/X9rPZVRV0LWZEkr80BrMgPas1ZIEuV70tQLgesStVMGYVQI7f05Lvo4
VyHBe98DOAIO14RNjWkQ7PYFmq+c7VoEQxqthPY66Kupc++R/ci/rrrY6YOWVlw+
zHsFUY7ybs1PK7vhiRSayop37EB5tUtNv/76NCFhh/ZvbEYVvtZfgjntbqUluPJ3
lUq7af1/H5Nc5r87lcBWMWwuuhtZMKC+IhiNG9w3HCDVq0EPc1vn1DBZIXeAehwm
eQjMh02w+Fvx7Z2vZwUqlWUtzB+F2mEOBNDal98it0TgfHp1qmuRF/yd3afXQpIC
w8NdGogZ/f05OJB0p3ZMrOT4cnLvIqwYyeuev6pLDFls9/zv5h548E/di9PZLKVZ
AfSPyIFna8wlPKjtjeoEwxa3gUbMkmwGGeUFONCZn7+Iz6nT3/XFFnuosJI3SilC
y/xq4sraRF9oC16mxj8g5NgOwmFlg7rR9okt7GuabkIV7zLBPADywdgoXVPuGWqy
PFWIbFIssQTIoNLI8doM57IhcHQJ+1esCjZ7cLmj5M5J51N0ZTJ7p+DwwKN2fcSo
vgSzXJ5E6Hl8zs9N/uzf/6ZC1kd5Qvgf0b9+cEU2BF1aVSO/mUW7rkWNdMWLXHcd
tz/HB8jLaisCIlsGRkL6Q1et1+yOA6WTRdPjysWAnFCqwZlAgHJfFIZOd0zqM8Ie
bRiFqKxJdZUbV9tl46CFjMgw5uIe1Eg6riZ9FMVkVwaNUkLFiaVZb7sf7IQ6S6UL
7vjyu2Xyi0xJth51QGziODyDGBHDJKLdxjMP2gnhtfuSVXgD6AzjtjzDpPTm6Oj2
BOGxltoTSzpjOLgXfFhh40Vd9mOuOrJYhovVmfBMW3cFasmywejKi1D3bUqPV1NA
87OL58K6QL4oJbtB1sn+32o5Y8IwU2qM5sIPnq0K0Kuyw/tSecMLz0jBWDanwnus
uZeIXIh1UmmH11eec+llOutunctBI44akRtcC+eco492Qilk2bBQuU7GSIjxDBYl
Z8TDBi/EiRT49Vqy+nMeDXq+J6w/yywN5IE9OeAQ+kSq/rwlbgXpSm3o/YOmRCZy
zhFkwoiVJeRQZPrMWTbCbeifQJsorlHAoimbXiBxQzEp+Uf+GAG9a0zTfrebhISp
zYXjRxK0oBBVqQjlZcQgNM/AIQi9iAafxd6oiNCVTwC8H0s0hJ42ZlbbAM9AjiDo
hO07Oj0V7fEsg5YHMNozaADMQQ26iQsJN1PqPpIO6wvXP1lU/GPGEVvAd+HNTkkK
t0GMiCBbq1c6llkGb0LEhujf3nZim0tEQYe/nLR9KXXbtGmwU9J9G1r3ssEDI5Dy
9hXhVr6Etdqb0Yl4FJr5lA1pZfnvaZOoqYGjUTPdSpiaDlW83Avz1K2+t1KMNU7V
VMiWVMznSJHAEhWwc4917s5GCz3Sp6Te4A0Bj6YnOvYxHkP1OmRyzU2kGlvaRZa4
VDosm1u1m4idQ0xe2QXRZtD1jsryszvQSxBpdVI6qUaJ0n8BWA4hkt4J3/GZcmWU
/SPVCNdOgTf0QMc7QYAIb+ieSX01FKsF2cYFrYayd8fXbQlspsA+r/0VSzCs5513
4i82l86+bo+LlTeMveUO8f7qPlwaZ3/ad9ea33xvhO0om/LRnWJPBqpZrlXqSTdB
J55XLD1sX1pmiVjo/uTmY+33PgcMT6D//8SwtVhtoTQJjkMcQo/s9x7u7Uh/DvIC
uGwtQkWrcow78kmZLseTLAIThE34Q8vjPrqEwbEsvZTLyGX+GKAEuOfJ+hgYf164
GqdUAqBhHnbse5moQdsK4/LO14F7q3fMOpLFEMqZi1HH+q+ZQqc5es11CDUKuos0
ra9k+d/o/HtMAdkJJiHmlTpR4Hr9PYVhbUJlY5hmO6kenjsUuUzlOkwR2Y+XSsye
7oo0h4kqPeCLXGFQaOo8FPecNwOl4u90x6H0hg0K8cEWGMaELYwhlGOSNamIc19C
Fq6Kkbh1Wy9PneSC+asUiMDVvMteoZLbCmVQcMdt8HLSOz80OJh4fiJU3RHVDQBw
z6E8Qa9XYnMe5TnX2PdWJxywceRdqGqveeICXWtQL2eczLxuhkpJr/ndmk4sL7xk
r8C6T2hXYJQWkXjahZk1Yy22wD7PCPDkIn6maxbSI1nQkjBqYVqt6fb9KygmUaOe
JLrLJJFv8IpU5c3fdLxuEydbyxyd+qCZLQPpuCJItm8fHmOgT1ESQQUx9vu74xl7
WrI18RKvEh6WpV+dkbl7jE1SeApQpz8On23Z7uQ1Meph6LOTCKPE/TFTo8Xyrsrj
b7+EJkOVWs2tExXjAG+6SzmfSZo8KpGsFe/qjXf6eKu/SJ7kGaVrTap4SLLMJu61
0KkiSRO91MGLwcJOqJhMDuzYwSEyMjvdFEgjMjyzA/BWRynpzlrgIBWy82LqoVcR
0fRJRSxvQ2iLjMEaPZ2q689dPiLdzml/azsT/QxGeICipoi7yM6dx4OgvSCCg1Bz
g9l16gatKoH2KqtOUNRWLzx84jg1ajqFFiajWzSq4mcraJFhg7KUks7uSNcADYZa
6R4XA5KUmUD9D2ntIoLQ8GvBeojNUoYlgcAQCDLs2YNOEztw8qpmkAxjC5hCMyYm
3XezoZ8xwZS/5qOImt/M/vrew6ChChGmzH9MDXSB7qpVpUAggsWFMrUpXXonSNht
XxZJlTyXJpITKfFYiczQNnEAM4qnl3h/a4UhJa1KdaVIwCr3IfUPK6HmjmSMQYD7
ucc/Qtmo7ItiXx94n4WGTymex+RagrpYjEWxoV9tJ9zfktxFHEZgxIIRUy0JgFop
k57EgSM24IZRyH0j3R/ddh0+js4lMC/ekUsgxALIetqAAGvcNySPa/AvYrsaQo/4
Vh4bjqdNpM4FNYENOWlsfE0CSkXyx9XPVpoaMdBBEgJ12JsllEwS2yWdAQvSjThc
BtgatiS53NlAGw1yMkZxB/jKLsS2gOWZx6Z38N8xq96MCKDyvM2HL6pNvJYt0Rte
nmh6u6bEMnTvG/ulW39TPksbzL3R6kqpSTQXevVpIrt0bTMMi3mdPU8zoWddcVNr
bVx1vo8TKn59S15d0qBMMPZ9WipylxDhrSUQJ2cxzpBdkIU0NG0/DQwARl3TG+w2
+QSzoaId88vgbqP9P1/K4JtMIU+1wM6PlEypO73rlboxaMKrsaqNjvWTbLfMBgvg
Ym1f1Uk36HKzIHxfHlQxLXIDADJiwwB5TTaEY+BvVt4/5FvHQzy+syBBt4H3P1Qs
sDVJY6QpG4yLFZ9YmKb7b+14YOH0er7Z4pTNKnnIbVG+hIMBW037m3r6gwvHI4hn
m4GCAaL44YmCx+s5xioej+o/j3vMUn54dkG16zNwO71HUKy0pPhLs8rNC+XMxS1P
YOMVM3m1mhMVnwIstJIBnYLAZLv0R+12XwqylZ9+o1sYy+9/YhZpGtLyXSzj11xF
gZXoP8fAUdi8gfYbTIzEcJm12+NdZwG+PQzVpZZcP7rB85r0eZGXBhcMl4kI+C8Q
27PrXZblYL5/w8sv8qv3nwct2ZpL3bkFfZcQL5/L3+Czlo0Jk/waaJoRg9nl8Xxk
81yiUuOp7oNPa5KXRm8nWEN3RAcT7ehNTe2lBxZ3X750BJK4MOdnjI2wXwWBdMNH
751JyYdt2oA/laFOeVyD4ePaQTdtYygQHJtmG1n50MH2xrbea6/96egK0xqR9MLh
psiAzgDCiL81ab9D28QSxwnZrO14/8llJhGPmZhapRHCeOLVn9mHd3gGtuyOaVlC
lqgRLa3lOkQ9Rm3koyrrrD92F5DkMzCeaYxrtPc55+wDjxEIy6VZfDmLp/fuL/Eh
+rKHHmUBiSB7MbyCr7Dt/pGsZhGv/hPoNqfvG9f01dgkBthu6TEh4MuC1Mrh+Tk0
UOT7FjOBE60CTxiB5hSqcbvIinlWaheGIBVNtlSYGbPG8fQs8qG7ZzbXrknhqwgy
8WjnAr6mKWrUP3SYfsxUm6ClhmSCWsPUDuxRFWlaOx453yIiLT0/CaUXvR87pNAl
d3aXnbZJvmNUE1E6/v28k9RkO4Qduy3hEVaxa9VvHCFpzxlWRVr2QqRWwP6iyuIz
fxTfRvGOsWWFKehK/iEUR4mBKskYV7oLsBbVRqILpNNrMVdIPnykiR13skq6GGGZ
TSGuPG8hXMMgyu/KkalXvlYLNuTNFjC9+zQgNBidz5U6tRLjRGYH07j9YdzWX9eK
Ja34vToK954z/14/tRKOo2wN5lxRSLJfT0Dgz4EvqhL0Ayd1/7FMGlT1z3yQb7nn
SPP7/DORgGSPd8No0rbPlPs9suZxkjEMGwTjANQ8RdlCSDuJS2TdCbgQQURVqfJY
z2H7ltcbkBSf8pvEJlXSW76L7QHtEcDBOYzJakJasZ6+PGRSCs03l43Fo7IHykvN
zGDuDXhYNQ1Ecw4On9FqrerN9Sa05YnaQN/nviE27JyiKfZUfebiEG1499YuX11b
bD701gzte0HBJ+xtSXdOZ9X8LkrkIhvCB9AivD2Xl/QudW1qFqjSqgYA9k60jy6a
wk30HzD9W/eT03gTvPTPlA9kMulU0QzSYBIMlTCHHW0GUYWmXoL40mzM9Gp9LiTn
gZQBcLJRNYx/o5RrBlV/faQ/C2E9PUw3Mcd0ZYZ6bGJABv76+R5Z7MQ1cDXSDZpu
8MBRGEBHTfs6oMYmX+TghzowyLGIPmW1keZpp3esmbmDlgdWIqrrIoC94aAyydBN
N3bjgkOBTlPR9qanMs0mXJvSh2RC1OBsVJP4q3lUEQ4LXidpRluOSdUE/vGPvLth
q2xl7dTUmhRdya+145uYNMLcd9R8Nlyrkdh/pkpjVej+OvtrTT1LjZhtwhQPyhJy
vrkfhGWw8yr54sQEljC2+iWdBZgZ/oU6+h3ZyfVsGkx9QHYlDhnL1LFr8bmVrPPz
OJJ8HONLu4lmFqoFPW7uEyhGNeoS0h2A5Uq2NW/+NyhqgFPMHqgofHy5ftalR/+g
UrGttv/y0Z5u3uaIA91ipjuP4hlXWhjFeUWlb+aVbGCXF1ve7VgxuwlsaocVH+Oj
OqQw6ELxmig5tiGNACoXM2pPvYE1rNVj2DnpU9o3VXRH1SLCwWCm8vAzC7xXi8ag
t4ugiU/C6p4TGiHksWRdHbWtUUvMZ7LOWiw/sn4r5KysKfncQeeNQ9Totq2dJ4hT
QOzCHX9u12JzJAcqfKvKcTnJRD31q9S33MAflKOIfEVNsLgc3/7LGaFNil+bDzCP
2MQ2/x52ofDzRU/2d1rFiOXt1mx7B9yf/IZ3xmZrJA6utL7poag83RY76wePxjnA
8QqLz3lA9iYIdkJi1w7TWBsiBw2/7cXxf0UuLFtQ7Caknt0pGPIV48Y+U6kC6qzs
9lpQDopK83VMyWbjnCkFdHpqZen47dRlk8qWSlXPO+f1Tz05HkmWXz9yMH5K5h/+
uMfQR69CPAGMipAlMlypFfFDM+SpjZokZJH+VucaKmAEdq+W7JPByieOJZeC+psS
emHlJBsghECiCgZeYQxQhiK2gZS6tteNpsUrPP4RVTIKqHwTRpJOIF+adpqCfiG6
06xTD/d62EzUGrCYyZZSRbaxrbHJRW7RTXCX8r9sqw21MeKmSDZNpOitu4U1VkiE
02cHaNRNFHFWsVO4OSrafJPtgW+DbQSdFsSate4tI0kJQdD4QZUnF3mH/V9fI2o6
A9xA38pwlMXOjD3ckOabV0x4Wy9u1ZeHtwVnF7YogzJmx/g9eFCmQWC9jIdfw9P0
db1ETucolBzLR4qRstEul5Af5VBhUacRK8aS7lRLZ+qyHK/hkANwe/LTdgpWblgO
D5SEXiC6N1xQjb2CgTyegcACpPpKiOJqGmMtanMDWPfBoIdyhIckgHmTC+Bp/V33
e/NfIUPkx8hXyHLIU9/84TmO/gT0N84suEwBwVB6jjVd4KYO4QGtA7S3I3YvSIf1
ygMPv3eLGoN+uqNrKOrlwlxLJq95gD/v3cOsPlcxynGFYq6EzvXyqc1IO3hz27uU
vfmtpHK4CjxHY74i5+vcTyH0ED/jTNpCw393lMfPvi7fkKcj0D3RbIZP72MNdMJf
RQAq5hE6N4jfkELAosYn/vUdj368NFy7oR4kPexBamMpBJJkU5z5Q4FcMtMRWwso
4t1b3Qn3Uf5ISCqrP30fhBxxUyCcxgdfzQpr+ge1KVBhMD6lBt0oqZsaJRfLkqN5
wyvAVO4kWTSn9pbbBfPCfdeQpmPqIcBtPotBdwcB8HSo6oMlGf3evC0SypIYIOj3
bzcgKKO7SNFC8d89pKhVORXezNI35OO+Wh1gQMyjaADnkBbuczzQwnwRxxJTJ+Dv
saHJbAodJ7FRofW2ySn74nH/psvAaGMzfRczbmXCLpfHa03YqGldojENV3CLdxq3
ISOvDviiGPtrGyPp9gLcwA==
`protect END_PROTECTED
