`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/f7yc15CmDkBNnv+maudutYtUznkyCtUtQwi9GTetUr8N5AfpOqku8dUroBOWpWu
CgZo/J3mxzMOuJozf4ETivD2CIJm08y2CPtz16/+L9dbolkT9jodDTDSqrh5Vs9C
ymBXVxFZxIvHBBmfNsGkBpNTPQxQhJVdJm2HtmX0sENz3E4fT4jif9wxO4VF6Mks
I9Z5Izi9tZsq1S3YP6a30EjYGfF2mwGGo5JGqhyMX8BfDkDxTNwR2qzKX/p5sIAf
3WqGAuyOW/eJX/v37ouBiSCHV+rG8Ej/gf0JmnYLt5BybQnmuM96GB/Kod0qzFVc
pGMGVC/yc5khXrz+oQ7QqBAFWpxqwsATRj6JGjk42jczUQ1rGryGrXtpy/hL7rnr
+B5yCIscBJgQcvxTOGkdB7m2MorI2e1OUna0+r1k8Nr/VNILhVM2f7uSbRlCKXN3
BZnTNNOZTMvsj+9Gway5yqT/v2WP5gctdt8u/9gudVlNTgycTI0N3ua13bUkcrt2
/1APQ4jWhkgSX1CLmxXM/28UIVb1KAaNdkbocDuXzT2TEM/zZeEtMHX7GyJy2KZv
/LXXmB7xxlSmCjvQLR5mcPKZeJseKATRIfOZgMrtlzsOwFA7hn5EjZ3S1v0JbVBi
0f1PpFPAUqn72JSeCt3IZr2UL5iBHXGNsFGA2gMhn9Mg2I/PepoFIfTGJ3bi4T2O
`protect END_PROTECTED
