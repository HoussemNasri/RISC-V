`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GtoNuJJrShm8NtEWIfnpoliZaq0iFMV5UonpW/FCTIWxySo8il5krV1uLp2utJfu
EtOO+2O1WoR5XZMm8BeSryft53LICorOhfG1t/VT8nwY1ixab91748yL/VBHzZLG
u5Wv/NVwpjsFS6o8xjacFJUyHgwoCrZeeMJuTo2KajospqT8FKghPhMd/J7mCle7
ba0VGAjhxCDHNJYGOG/f9sbjpR2NnaJZ2dCZBpq1ksmvNIAob+06+9N72VhrWUL7
BdZSLFmOmvvKloIdXi7Q1HDsSvPl3+AwlRU9oWrd1Cxy1lr8KQut0/CxnomCIOf9
0nUWDbwkhDkw2Yh3sPqrsJPA7lGrsnJUMZMumlGPzxmlRDy4uA9Jyn8hFsP7Sp55
7KP1BwMMtCJcafdCQjk0wzTUDveKcx58bNR+VN5ulGN48rjOoHDILfNV5DPU6Uh/
1k7Rah8dLBMbvoNT1seQZA==
`protect END_PROTECTED
