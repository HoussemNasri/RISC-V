`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IwHPnfAF2Zw16DbTgeTJ1U6VZJgwccZxT82YqhwZAHcYgZs/iAfdB5x8jFI9esDy
7iLxdPWqA+e0RJQCOoKl8GDxSNSzIj+9N5Z49xczHDetemhNDfUqu4UczdNdyaqN
6abpRYeq51IjUvOxUM9VZRqe6zyuUVbZqLHvid8/mdw4O3uP0SIWpgpVwRFyb352
Ar8MYqaZE6ZDmY0HBJJsNVQjtPNgILwbbvz34QSu8YU3fN3d7M1tvmXbF0YAR8sH
5iGVAqz9rFPGofEMq0GSINSbPbOqO3GQGWa/BH/OGaMEA2GXNhkfftgD88COnxAf
epLRrSg/kmsf65SvExJQXgjWukhRsY2W5hQT/rvTf5LCVxYd4QHfdop2Pzh6IYe/
PmoQtnS6+9KSFmGkCSA9oFJyXxqAhA7D9bHG+dsWKQO/N9uEVqF3GEKh73k4Ij/0
FxPWxOPIDvwmIU/C/3uVVJWE2b3V9vpNkaac/vwd7QwQVYIA0vMEZxxgQH3qdWz3
KVmPPDIE9HsIvuEuAUkBadhEX6WBz++IAnfBXiNy/Jc/NNZ2EyIQdkGatPXOwg2i
h+mrXL8gFTHMgdJOnSbwRN9tt0dwLsiW8gI4/VpYuHS+GW0k4jFyVGV6EK9v9uG1
SxM2Nd44MQr0Se6vLGsewZe1Qu++LZowxjMjFXH8mKjWlgTqBf//hhlr8ccGp15x
Q+W6ybwgThaBbutbzW78/qhMZtHFrepD/GoGmo6rPHGf5Gio+wwjfmp5iz5ZmzdB
rdU5OGwcp3GyLsoTaWqyD4q7TVi6h0fpNLtTMD71d44ilY0cT6nLXlA63JOKnTY+
OpGpgQsj/DO/6tgWHGaq/3udiadtcU255C5O2lbGysBPhpCykAAE1wl8PVk5tjOP
WgXo1JgadN5BEiSpVxTRXz9LqmDE44THzp81rVC/y8bksXulI57CD2pwR2TI1sj+
USaPAYDbCs0gYIveeEicULH4qcwQFoOrtWRiFxIuPNwC7nP4fNx66w1I1xnGFpTo
If85sCWPpG03vGTls0jtwiXHCgfrPxv0R11X9Sxyz+GF6jq1cNYHvdvNawF/eHuY
G+dO+wTHNnGpxYZO/B9uQfk8dREYDnz2wVX/1877MpjFb3toZPyEAQFFPGD5g2ZT
tgnavk3D0c3pg+xOCJ2hS/YQVEfJBy0ZXRJ/ZVDXxeEYjzQY/FMldGTaCsFIb2vp
1noWxELRXODqSkD9bgJjMwMYzezDqo/3zyRT6mnNWcG4zbgRiLgLjdW5IRFeBTNd
t2/CP1JaxG6UgIaIORSJFsCTcs0JSymnfQx1WoDQi74oSL6EZcesT8kt5bpnDQBw
8Mpvug52JNvzoBtZLvW964jeruJVqVt6XuunhO3qtleP3Vqf1mOzjyYJPytlmobv
o54V9izYjHGp3EpAnSeSzilBHYSYqk9shma2qm8Pzxet4mnDW5XK0tf7SVFA7A1f
L1nbuifUnyjLUGlANdJB4oMGz+Ca9ngv0pnWwietWOejNghWRZKWVUp/kNccreeS
92CeSNDqvZ3Dg8us1OKpowGz+MBhffNzbmZ+B8H7E3l64yAr+REACJEMoXjB8MeR
u1NvcgwyCw9ci9jv0wFN4hT3mZYExS5pFavF24Ue6OubaDdephUI2Uo/pksR9UWF
nyLCaX647eQfaiu1cKzxfX7nqA8EHzJvpy6naFkFekSXIXGOlpozWZ+LrGmHeG1U
KERfyRW+/r1UDBBaHjIv1R5pnyWk/s0/x2fuF2G2xg1073ly9vXZ9aNdf9/tM1Vk
09lolRTP/kVZqNrOHCr04k5DJZPV04YQyLDtB473IKI1O2vk2S7SXvMFVWLmhdl6
tRFQZCHeJPxfcATqS3puBdabmV/FzmztHebIhZxO4mJqrbl0qecZa9HXOoxaL89E
sPpj3irP+QQE2QuwKVfzysPSVB/ko9Sezu3WeNW1peAqBI8GKSCaeV6WwK2bHk9L
6HE7IlxNzVwN8QFis4/5uM8Yt5s0B3RRVoc6/W/+4BjvzW7r7MvGYLyWzS3768Z8
8Lf9pOis9l5k4Q2w6ZZ0+DWTn7Mo5eZ26oXy0MJZ2dzgDxEXiWI4HLibJpQ1RaPl
2ADo68byaepjf7YxOLqFMo0okCXAMvHrCjkumLpEnk9i9mhkm/XW8X5Fx7pqzBrE
KXheu9mLQTGxU4LrAegW8LgkLoQbO53rAFmjbOXWkUwmguwGXtGjvsGXimN5U7bJ
DS3u9OI6lJBlZD2i3XRnS2Jbu7zYpx5LDAi7WTCUIBRnJrQGN35d0RfLSTOEyqmv
wRSIIGX26whRdb4SjDOYyWHAhL/KOlsYKArHRyqt/w3L+2mPYaV6eQRz8RkD+SsP
1yb3sJxyXz2PrGrQOD7dYLQJ30eP2Vsl2ogdWMQrA9DGJbfGWNYtutIWe9zxnjPp
Wwpx1SHedjw4jfj25aO0WarmZ5fqDgwsoKg2+AX3db87p+Qmie9i7noy4bCTPHHq
xjl5EoOhONC4UjvzYgiY8ovT4fMgfX0zrXqDnbhc9XIBKKhbj/69pmFpYUJY9nYT
ZoOakMS6wJrHerfqHhssMrJH5d95xbZFgHCF7Wj2hNyxt9xQFiCbc/I0OncY1Vx+
bg6PrsqMEulL0mq9kA1S6Rhh8CNsTU+a0Kqo2t/LoRJOZ0JktBEmCrDOakpP5vCw
ROlt2W7juboocnyQMTptK4VniwFeI0ZkMN/1DI0tdLMVZeHVlZV/kUbKYP8QVN6K
04UBLpIHGSQROprl2e+iEMMrxLj3ELqaD4Wr2E3RH7f6ntwX+qOdX83tR3ymA2lI
uyZntM7e3hVCxF+g8OZOHpyls82Tqu/eCjt8EPJsfhD/DOhtUxQSOYCcoFpFxfzz
IE68mipYqs5UahSb2wQ/cucleKL5jSB9A+j2mS9/4GEuSRIvOt4+WGpYQdWv1vNx
2KBguFefLNrEacoBnTa1rJlCwWBYvAT2buSEuZRX9EojlPpllcV4TmneoJAt+f80
3rCvsCnvifbbhpNX/SfJiUHVamIknHnTNnAjyYAd0BR2ztLC8gw6IQDI3DB66PTN
czN+MnP3YLkbPPvxgsbqXfJY0igtI3IND6eVEP9+KC1ZnCP4TOcK4QWIMqDNe79n
dIXdSevmEVFLNo2rNOeW2veLZHGRSn9v2lhKrVak0lV7ofi0eb+D1Uy6V1ggDhK8
KRpBKjl3L0QTpvy9bmL3aW5pHB2a+4f+9IOTQ2bp0A8ljYYilE+uWqafZ5C8Y5nM
mvgQIvro/3w8k/IKmjzcxD/16c3Jbe4+OiA93D3z+2UCQ2iEhTJi7whJ5zXpqgCR
e1ocj/6zpESb1sAB7xaERFO5u67KwgsmOU0FZ42xxAdWosA0JAJrw5OGUtR1CHSy
3z0S0Kpk8XTxoVuJK/kFGJZGH+6thVEwLFGIS1EHrBOVwE+lJJtdCynfUMYW05cC
p/8OXlxgbomB2NPX87yYc88IicoAfYsPUcn9NXEnEiPCN3Ms9KSgtMuRZcS/XmD9
+pzZ/YlL/0JgtDaCWQvzPUSJwrwGHcrCB0Mc33zZjvAgC5ulG27jCeeJfUm+N9fa
mo9XMjh9plnVDIT7gq1BaspYCPfOXWrTq1X1/YCPvztCznjPOk5G04+8+W1od7ln
uJQvJ0Si/Yrkb9Gyux3TV2M2puaVAJqp6n17BrETjT/PUsU+jJF/1bgHxsl+Qi8H
bkSgZxQzkwtut8qaOkMhjL9vgku0dmdkrfHnu4AAk5ZU6d7BRhn9mMGPzkoZr6uO
KO8Vz3lnOJw66iyNeCg29jlNHoWs/HHvhfUCWjJjXOffrLNVbzzPY4JMWhPk7sJQ
R5TPCuSlDtbJrnixa/1eKBb+oIdoeAMuWBrVNNzQt1AjEU5G4g/44UCglRwkNAAj
0eJerxwdWFVkI92TAVvDPBwP+w2O6SJIk9lCNNy6+nS7wTolByNGeTBuVC/32uv6
G5EQBw0zDKLY4so3//Kq/PxspojwmWgB6QLuehQjrsG8C9noRu1MD/P+S483pJb3
YLA9Q0dGjxVZ9jl7cLnMdrxU+m5EZ2OIoO/aC6d7zQfkSe5Xz2e+KySgYMziMPXv
FlAQ4l1zcfXRK2+Ru3vF6wsRQZmxfgBNP8nk4mf571Qf/hyLLeLxIpFSph7xasXy
VhQNMly6dPQebrFUZh3JNQQd/n3+Zhe9XUSPbZmwrk4VQ/20XS/CbSLLaAl0Xx2l
2LSXTqqPzesjrr0DSPfboIwqlzhCqWfXQtpq2+l2EkQTHLPfQlrSkXqc+Fw1r2+X
x2b13478B8VD0AAi6w1jDVtue/C9/h6lOWil944C8JqsKONf1Avt9/OwgzJX7W8s
lUTxRvDBoHoPovUxXi7XbybQFB0V1r+ahxx4gFUYePhw6e5WKPjwc5iCuNiwCPTw
Ax8dkr1R5DX+6uNdWDcuZv+HKQLRdLImD2ducgsFEN34fgoFbbZ/0dggQPTs81ph
U/LNVauLJVgYxj8LP7Ep4KT7lF66sTNsjfToTnWA+0DbBNLhwztFL+toaQXsblEC
Dt5j8/WfxopraBwqPA9EqWUMfZ+eqwoSB7RQNrJ4pq1N6izE9lpbCbnVEBBTSH9+
ToqY4SPzq1l0uV64V/c0K/+VIDOADWzeiG+s67Y5eUGopYwMZ/rakTMky7N8hjxU
/2IzVszuzMZDGT0PyNxOeXpPa3nVjYYTbMMuSuDb982Y0dhDWSht+i066rTWK+KL
+5TqQ3ob6NuGm8CSmJp+wd80dtHgpA64dPQCWJHaIM09LpREJ/G27DcDcvqTzS+x
8me14JI+hmqOsRoGavm5rhqv+/5H0nxkOxxwuwMWuIm5US4u73XlkfSLNpRbhOYr
tkum1qfRhKmJn8BhXdGYpDdfAQZ8N2vNBwObXb0YZmtV9QRP/rQ0eeJUAlMzcl7g
o2B/qJ9CQaAclDVIrc+2Af01HwkmPiWAi3GMM9j5VaGF+XS3UUWivoV5FX/ZU9SA
iZzTxjdr7DDzSF1kBV+8GlbnOomLNusbqOlfQJziMOROZOKpSr95EQ6yEN+aIgwJ
tzaNUnHNixufDdiB9k0mlcx2qcwJdLk76mLX+Z2LKhJXIuqUKXdwtllVjRZR3Lgs
d0YxMItz9GcShuBmb8HTfAYPaNApkHN+aMZxD2Hnuzqavo0sUGUKcKq+TVFRSQhk
/imX5+O0c0TOl1ceAHK36dWEhJYGLXHIcDZMThswr7rmTXsfNXluMsbMoD9oEtI6
pMoJfNlX9CKDDd3sCsZRO3/jxqZvL7GxJMqxU0uHb7l886VSRX4866higBYSrSzy
zEHOLlgnKo5Std4nR/zDZWE/8RLAEgdLfHdFdzB4/TvjcaPwHoM8fQvTnFkWZGGj
qUHfo5Kdx8WOk4i48THG2Hi8dS4eAGlzuc9OmHPcNnwE3RLxTWnFWSE3k+lYDW2m
NuxABzdX/JD9aX3IJh9cwL/6pYXLut6sK9WgbdTohgnWNhLK+kfP0y3Z9LG+Dea8
giTtNRTK/sAWSB0PF1LjgvHzUFZAcUI14n9dOy8sTw8V3yscWUzzITObCvHArADL
BAG/h5gahbq8c6MtXHhkp8PWI7WeDHOayA5dseTuW39eZsmPerR5ohGLkUI+PvPP
PZQc/MyayjwSgSchtt9PWMqJzNDCD+MY5ok3w3a+lUuhMOdtHqQeLKPmBRBNKROw
UvmmJELODLo08zUaWnAQh6wXh368iQbzoM7ezWkcpA0CoH9HhL1e58YcAB2hNp6w
QwsH1GkKqzWVp8SiShdgCw0ws1XRhbcwGKuO4wuJ3NpPK70HFQBndzRLiIDcmuQT
COEMtjzmXhEUk5Y8ZLM3O1/GaguG+ClK28XHcBlUO37KZj+bYk+1V0OCBAnc73dP
U1lpWy17+EchAzfrkWhu/rSyEkzovODsTmNVUq45lMy2OIY91Xn7N4KUKwqYKoo5
afGMReqUA/y/VrfdSdKnae3hnQtVS/2LMB84RDfbOpToDgYAFA7e0U6o6916wmKb
VGgIvRnzFU5F9tqlik3XfLCJmrUqZ33wraNOe0XNrZ6Rtk7TOebDtMmGF+sXa78e
cFzMGLPx2UU88T6n3+Be3qN+kudDyt6pP9r/UnHuxWmB793fCHjJJB5J1S4oAndZ
goWVShxPtdWWZ1O7AeLh+yNSJfRcDyEHajwjyZ+PN+hUOf7SnSH7sl++9+cgcFti
PsOe55dh2SWPdpY6+x32IrjsqOLw3i4HP2fIJr1vcZvL7fJda4F5PRYpMRorkLl0
Sl0iNh5OizsvEypdCxTh9JbrqycxAHV9tWfu7AU0iocPcUfKroASU+lFApqq6YH3
LKjrqO1lhMIO9GIF5VdZhy1lA3t6r/1uv6pkTvk/leeb8wvgTHlBYUx2cdljZkio
Y157cJdDh6hrb2x7ub0docIlLO9HMWixE1Gb+wzJUcQNi83qgQIiNM5rbMA4zRvS
72KAd+JWwDwgqNceJcTjpp/hpBeWLx5/TZcGAG8kVO+Jd6Zdjw4RWrtqFJlVp8Jj
Wm66l1he7SqWAciTbTfSrXpdVV3S0qjK2SCcZ4JyQEJ95qTH1g54oHpm9Axqzi/N
+GJngulvXK/VGMXFUmQpuzO2udtalrNx01nrE5PfQFwUbzlyrYyYKQCKnr/eFLu4
LLIzFnHYYSl1/fY7ctrmq26W7aco8pQRuda5PV8SBpVdICC7d03YqHLMVufO83K7
DsSwC4yiQ7jV/GuAtBLlAxIMg77Mq+yV+7hKF/MnynNZsyYSPDw5gR8U7g+pB16h
Tt/JUL3wNfjbBedseEmTmaUft4vKJYrZbJAfqZzUU0/oQ4HlhlCojfVB0x+eMwC+
5dcQkY0iwIWoTzD5LBkdRwPIr0T8Bf3LAzTQE/8urMp1m40YTs8IncF8L0DsS1PH
gVRvnOScZElfJH+U/BjgTP5y0SDU6xNIvycvqKHTsP4MPQB1i6MdNXbFGG0nzqe3
Wvdfxd/V492wuetAz3PL5rpzECrKs7gWDE2RoB5cB7qIsVMPJVU1lRDLnzB+i3id
Vw1UJNiIDFoFYl7DZoR17bFtfjreVoVRWDt78NrfL7PX/U0rSsn1T/pMyVYn9xwh
sMAQ4e84ZLEBep9hmthOhfKGPm25M/DS6oVNWKDCedVeWFVQWoyJK+iVDh5POBdm
eFLIFY+vSQtmXxZyaYxbD2uAobNf82IYBKcODsUoeKD002vJtOHPA6/up1NEdlie
e9Mp8gIz0SHMZzGUyfboHonJoXkCoWlV6one6BL5pXPwpEMsIJixmnF9zVle/S5P
nk1VCwokeduCcaMiTgsa5izu4SeIB4YQQwaBqQKSUIRcaP+kLzQu0Ea6Volz69Sn
LBwxbn0DNo5kPlS95gpZgCGI/2oIMwHCD75H39olNV7ht/9tepYGHrYq31MaCqbC
j+WxypYqbIGZbVoBCr77rPyCFEMchIKo+ILv4NgzhCwtmnIksbvRpbsZJa+6QkSn
DcZMEKGoNyakO1vNIUxPy3JCi+VkFIMf22EUNdPQndIZcLPiYHyJSwqAdGXVqIoj
5dzfxjxx37DVGl7gSiaOxw7X29O2KFhyiCuSFhvnqqzpFXQe2noYkM881tKGwHtd
TpiK8EG2ii9N7aofFiaB9G8m7S+pT6cnPLL5/bXz0M05DOillnXFsNeLYlc58NIC
hk7u4r/W4Ydp9RDLIM8L+1mQHd3DJppbVjwD9v/EKtTU+v102USio40z5VyWnWkI
Afs634aGhQCv64j8hahvVNpDlmHX0UD7CqFzeVLd65g/37QWu13jV5lpyg5Ur/U4
FGSi1uws5phKa8/wt2cGVnUmM3IUSR7UgZZSwzvj+nLr9+3LIDparv9s8lSc8Uzz
JMAnzlEgGVuBEl/Bhrt8Axdew/rhH91j/thzEOeo3DJR8yBpfrLp1zmXv4KRKj23
8uDKPW+DefvqIPxmWGgm6/N+I7bw0ufOjwYJxwR2/dQ8N/LeYvTSWOVA/fFKYzwT
yp3xlBh6I5GXXmqaAPr9ryoWfcVVVrYvqt0h3LRtfbFmNOcapZIMjXgPQSmladxD
QGl+qGgJCYR4M7wsZFtIlM4D2j8o8XKemxHDus8D6tp9LJYhEuf3HHBl7PxKJzQo
4xIzupHQ+lpGE0u/oND8fvgY6yu1NwGsuCSQxSYNoH4V/rxBhWWQm8b7Z1wlCGGk
WJUYjWfCUAidJclf2rG1mVEL0jRpFK1p/rvaj+I/ciZNtVLz5hMX+4ce7kuT86Vg
0mKpyaScNMl/etaKZtWZCoKqASSGXq8+zj4le9AUHzzNBIBTcaVfaNHlvFyFeP/o
VpxxKs0HLbVtGY8NoJsSfCvp8zaUTPgQIxCnqsdMXCMwSnL2qQ9VktE62OCW0tEU
lvEmOMPUhKMtdx4fqYYy8mFq9Tx60OS2MF20R0rIY0zEEaKbN6OPb0xwKBw8KTvp
XFzZb6P1s0D2Km0XNPGn6ftFsSoKQEXII1zYzaQIXD21PvAieMK6NYSAvWkOeYWt
u9M7hNg/TCS6Kg8D5oQTl8eZNcNOTMeQ3/kSQ1B3a1zXfbQOQcjt6qtX+UvBAx1w
zeWcHJNlWj0Eogjy4TKIgjD8kbcBkM9tLa1bet1IL2vk94if6MGZGkWkypzY98VO
9tmzfjen+vtCToYv6oyk3scmkgny7tdHOpJ4/FO+nW5ZcEWeSskPgQBoLjLCwEbY
GGkGkFNowAviJbHIaYqM80IictSUru+4SAYaZabFp8ZxCEA7FnmS0lQ1WChfvnhP
e9q83tJdiTd3znQNF7JHZ3H1UBrvNRsqDpxlAoK4JfK9Vkz3DmxiE3Qg/mXleTwD
3aRd58LU1x71plPA/ANPIRYeQ8yy11ELuFSCC5rm+5xe6Cdw5CPlQQV7nT5UgwsP
ZKbP5DxS6wtBG8rkJnMrcQikOI34P7mKjIbg8b6WUL1i1mdUlGQLEQPjzIN0R9XU
NcS/ZykdhK9ndnBW1C+5KC+nWKryrnx4Hx07MbUl7lgELHxK97n0IJhC4vwtiH3t
LauWxYkFcsTUqVsF/51LWtgkOhyJAYQT0g585VyrKmyxjzxTs+DzC1B9rcbtz2bC
Us0G2NnpBoFFhHaBWwe72b9I/64B/MNtcLxP+DwvbKmJwKHkjwk9wnK9p4wEMJi8
GCpxPsCVLAVHFZ657UDbyDyuv8Qik9nH0tHHfyB6KxORaxRJxf4EPKQyksC2j3m0
RXwpPwrKqE9FhRiJTRPk1oyRSdRCPYW/0wGuPcZCLo6YMdLKD3WRP3QGsytL9PPI
EGAsBoTsmQg0wsbIGnL+zrro1k1zAaI61MMDFrdv1QVsKVlwZuh5j8WzkDuwQz/x
n8dZ6W9D1AWxNt4Hrx5oj7PL1DJH3sYf0tD9kfXwY+DHz9eOO88cS29ToGRS+HYM
r5JDG7xY0THKLjOdnX4kQ+/nFH4mGy+/J/nA/gwj4+i3Jnt3MTo26R7M4bbPCXFE
MzbgjsUckOC5b2wSTov5ymI0n8j5LPMkcg8B+9I1xHYkd6f+flC3vkytdZUs1yWf
Z4y56Y90ZEkniYc/v41uBix7lGgBp5glbTmz3vFez1tOVizwR/6k11mOiDcyB7Fn
mAhEixbs952lJATIxX6ubp0aGwgdbRJwtwXJPL0q/QdsT+icvI2cejg/GB7LdKBK
x6BgyT2nRsHSRC7km2MzqD+ET0sEXfOiWHYE4KGFbMqk2K4JCuCtGutTf8pIDI/o
0jsHKo5trRXhpo4C3LTaZdBSSc1OBphp0bmrBXrVfpMhXJojw3HT5kD9REHS55kQ
SzU00EzO321To2MeWcNE6DNmrIdV4mlWnpblBBPQ5eGh3fNzC6LaEyWu9gnPhwvv
x3OFluxi2oRsLrjkGeX8MMK/wSZ0i18qj/shKDo0ePUh1QIAiPetP2cWREHuO2RQ
4H0ecXw6W2JUP42doaOjuWSKxwJ7WRQ8uVOkSVoAIdMOJpcbFN9pBcX8LZDJQ7L1
t2Cu392UyOto1COvqMzYmS25t21BefzyYzKPtib/2PdQaCULgO4ARuxX04RAxUlu
cAgDEo/1qh+HPaR/6bTj66K1NmKPIZXpG/JpjcaQKPgwTXcM+wkEooDYbxa5drtA
zomjkdfSn2RhsjztLFD4YKGW13J7TeAuwYqezFCj+VAd/MKavFGrDnEi4aGOoGO3
WWETeAW+ptxgUIEljnnz9Xxyg0K3KoezkR5SNEUPBGn9DPXboantda/zUjQqdMv4
Lu3UhsxYcUVTSiq0jzaQCo1w2T6z/09I5vYJOMfTJFRqKJTsP6xrxGqPzk42pccg
L+I29mCUNlqeAM/XCFDvw0L91lXMZP10XNe5VjPji6QjR688Fx1whozB/j4DWPge
j+58qNuen7D7OVvPZttJpLX96Bma2BFwHOaGNS3k8RPM64hvgPy5SriaUgzfqNSq
k8KbcuN/udc4rePhF7newQs0OZJ91OTvJgkfEVAvEJJp2vvGWWEoSiJq75bJk1Ev
gYl73ArC3RoEN/NOYIFdXDf0FQDXTY16C89R2HEVoFRniLeN2RiouAVBeqQXxnzz
qnQy5M6PW3Plf5SZqARFgRo7KatovLWViZp47n06odFa8/gVn/kCSpwTUujxXmMF
rypZWTD8N1KW2ncXZ7qJY7SA7ysTXu0h3lQXEhDuWYRPIIWHupy2yLAIbW9MHVnl
qa2aqokMJjjPig8nSqam6UsKWpnDIqUvq8I71ZgrL9gBiM5lo3MHNSGHN6aRGt+y
0CGPn+4KpvNaQxCMefPD5SqRgShxLaOMVi3LE5iG7fBfQLG2UceIXftCVMAPmcEn
HabnYHPJqBAmUiTrEpso/zZIhQ3iyDzIhEoXOQ5Rt5IOrKKkGbpt26I4bL4Tdkgj
l3OAmu85e+g8IXaS40BbbmpYTKbfM3eap+ws7q4ydh1fGoE69QRhqqGOcuKxnQwj
EoRXPFR/cypXs5XR4S5XT/vftZ+XbgyAAo8s8q7jic8VfDxj276UrxcJqgiIxWvg
5o+d2slwfd5Rr+VIPR1VXbfvaWai7/IxvMM/i8EnDkgB7MwdKm59t4czsy5KQuUX
hKXtP4vHUuxsA2NZ2JbGGpjcACcpaKGCAz5sbQ//UT2iQfrTdLs2wD6PL3wSh87R
5IiDbwyxfpUvuKIxxsG5qMtHxT/zXLEj7okNgZLLyWd2SZvbvUIQNe6dVFOC0ozF
j1ZPC02zAbPSiGT+nPYzvK1loMTrnyDvExAD0Fqljqnh9JBQsc6FDShbZb9KXjsZ
ktIa9CzPSpSV5QX+OiNmjXPvnJ6EIv3S0oTTr/5EJXO+Hz0Bl7h73Iitd96cIlWb
MhAkFxSCS/Y5Y9r2TZBOkiIBBuxQ2uv5DLEStxj3uq9xQMx6c6r5jNqOnPbjoMGn
TZeTLCvIITsp0Rp0HO40gax2ULIv5nyc3Ot6Pe75khcQFGWhgw5erlhWveG+wXf9
qf5mREP3e7Ize03nnS9tMFZnq6ektFM1vPpHL/En5cKMQwRKnH1UFyk9YDgRYISs
8szQz8/R9MrclL8YQnOgqpP4fK3itelFiMlFVfvwBlVn2q+sfv3d6femSvdAsLlb
uWkzhggOZ7lyUyeXRWaOoN9rO/1O0NClYrrnSef4UBUS5i44gOvlKTPW7qUpDCsD
z7kORHL4QymoeH+moXy3lT5oYnOHP26JZLBO7V2kotbKzrwbLnUdpD6wgaZGiUx3
MhPPHr43Yd2CB/CFbhknlN1gkYGveb7A6COc4VwpGPHk0R9Y/4VJrn5PLKrbxkE7
i+q3aZu09DHdHMatb03DxAXy16fSGVpAehZ0rVR8rHCgC1D/ZEratER1foAoEl9q
KLWJMPOWT/WysK31fN7Q+RNtpvPACLAS6xKj2TXSZ7rTovADi+U9Usi3TgjlCN3+
C7yUdwFpOoTM7gUmsxxBmbPRjaowi0pUC1rJS5CjGkWj+6Qn6wEbNjrxdn/jljT4
T6qZEXdpe3v+eT1OfRDLh4DSMqYZV3eWNH9CyeRpVL89JtZ6VxZU5/f9Wo7Z+4mH
cj8tmj8O/oPDWYUpLNm8EpfU49b2dfxDURnmEEoV5q5SRBDfJVXIPF9q1xDaLw0W
4RMiadqis07nqTUMSCH9qrY1GSoZ3E2784Dz9lGcw/kYRNaj1kzhY4B/OxfW8g8T
vBmI0JDOs3O71mF9gdy3pqPhGbrxahdE22wKB+6OonZrUrLrhEna63k4Mz6wbeDP
B8pLRNepnEg1Hfwi7aIKyQ6O48L6feZVHPiSSOwYFGBH4589GKBA5NZG3XmuFLxh
6OBjVQM4JLcprA0/JKjpwD+3EjBONw2nUsTm4I+3ZGHFqAdoIaon+M5nVqSGoqWu
/zVXyAadu4wSaRlR5NNTlYTgFtYSSxDnQu5v903ICioJROf5RdP+Q8m37MCe2i1i
iUgOVFZt4yPDAShmdY5bpRWtSQCuFy8IvO4qg837TtPpmV2KJkV+/pmdojOxEr8T
UiG7yUpFG0y8SVTWGh7k/WzeSOCGAcaVjYMFIeWLAimXJAL/n0chPR8TBE/ySp5g
qLGsKmAIhsVuNJqO1z1gALBV97edHm3Wqhw15rs1IWovhKq35gf3QDd2kpIg84Cu
RuVNXujCSLrnX95BMMM1Iqvfg7SUdgKyCMzJlbUhjwvYRfsAUfg+ssF6vZi9xS11
PIYBqHfhmaE6cgVUYMToUo+Ol7Lhtzc2k8ZXdDF9izAI8bJrKdTeqES38oI3cY9V
i+DCQ+vOvmRsS5K78WdrjFSNZr6OB97UiV7UHcx3K8bcP3nw5IYpVD55vsPDyzpP
nXKNef6zuVHSialAZIJCmH5Vf80hf7/pJHt1KVh9Y0Iix/AMOZRwC7RzbxPn28+i
w/MhCnUSXaaSl5HnXM/sheQQqFqDCstJnM591Ae21zrtAG9EL8oGLqq6VwDeF5As
juAw8qOgc4SOvabg+UCdxMhsTRJgsTieSv/nhTxABYDg1KqT690DuOyb8stCRGfe
Owkx7V9uPprMjPhpgTuZRIcGoZK6ECzv/aZ2fkXHEfwup/92OC05ggI8knokD6WE
p2VQZXszt974Swthdpq7P1C2iu0GunslLEVwGGvG9tQeQ4EFqtfzWLBbH/dhGVsr
cXNX/YezsZ0hv3Bz5VTq2tuexxoHTFCWlOT+LPDAmCmkIyvqohRWChckVqzIeFED
+YjxSWRE/8j0W6ZXuCFMzM/NL6nRHLtOiFidJXD23cSk/+fhrplI6wACDLmjvb93
dQ9Grx56YG3yc42hyF/BUs8UTE6Ttdz6lTyfjLNXg+28hid09k823RfVUM2CMFjL
F/v+0Bdtmlahj4kKtdY/+9oqhtxfYTpCeG+C2RezEEVHUudmG8r2/qoz7q9LzRJG
rNyF8mCI8DeWWpGCKgNe4G5TPzNg0caJmEYlsm434wKj4TCodU9aScLONrOtMfjj
9vocydTzXZL9OkZPZ00VRE4bLqtutnt3L8hb+PJ6y0LsmF5Rz0YI6NwuvQZmX3w+
zR/axTUl2r6IUIE6YL5gEBOSYeEC4TIKgvsWdfu3Ypuk9MESLdDu6m1LwcBQIimv
tVkMQzSQ9M17c/udKT3do+ZtIWwjAND1eYiXm/t6xILr6SoeQl+UcAJahsAkO2xS
mUmp+NcvWajww1If2G+tzWhsJ2vYwknY1cRHUt5s79+vxb6cWJzEyGhOZ7ore2/C
B6F4aPSgFLMBso5ie3ktXo1GV2sq7xCg59JA/TKVyrGCNHbupj5vKQb7SEXrjkxo
RuckgYjX6HfEg4JhcFZCFG+rwtczVH/U0GCdZRoZ/eUWSlWbnoP6p44POVbOJSO2
xVG+2ks/ZVpV4hlaT20Lfak5ep4iIj4pSIDvk0tiUGRKTKEwb+C2m7V30ZtJkI66
INnQzNoY4ieDdhUssyrVpi3h/8PqNV41h0P5+viNcay5HGUfISUaaNseFJgYVgr5
/B1BrrsGSYMwb9NcGRKAdtC7TxcAghiLjMrGQWLttlJIkVa0N5w6ZclpLknYmTv2
HIEU5V0mRbSLYW4U+R7FUcSG+CmIcrDL995BNCFplVD6jWt4Po5wIsoNYqKYVigU
KF9bkcu1dYGfMNKs+YioN3yxPx1Moew4cydR6yEkltVUU5ds6QIDJhQGyFcjISsl
00RczjjPPxSxyFrjExhk0qiDrA422tTn+19/lksEWyW7jlUkzQmCUK6zHfFUnr4O
yJYVcnKXw8L5yMji2KtqlpwvIH4tOzswyUAKd4y2SrpWl7gvAH/24newA/kksNNH
qekbn24CPDpERcowmRkH/aNZ3rIXvAs6PrtwdaLpE6sKbwVUjp5uVmR5RivIUUgn
+bRp5jTPUxEZo7jrdMh++2NlnqMUNxj0mEhtjLMy6zj0fBdz8DaDW/c1YFdUW/3o
ohpGwq0+OXoJermBEzRk6xYIm808wPiACpW46ekwRflE0VxOT8mhtQAIProfwgMh
upTjBDIpElaE9b6h/1nYAhKTVIGe1c9Q1y8oJLS/OP0T/oeaWecJ1O8rFh3Jcxqy
DEvYK/Gr0tPvbXtGoKuoRZJa99dl6ygOCFp6xw3wQGdg6Z/47IA0GmiE/gIq9/gq
87m4lFJ1dLdyxxZhxpRk2RnmIJ30QFOCfBJJOMn9WjGCtiiE9mbNqVvA/lP/9ENF
ipcVoyTTUG/CoBQ38ArEcj64V5GFtSR1ypNrO63JoDLcepKj221kiWhw5/zBwOXq
qrGoXhsJfudw6HqOfPi1Cn1wS+hP5zKwE1L1xT7fAi+PuhHI9tEikQnUXTggvb6P
bNX4UeDUOIxUr/Cd1srBQmnlSUNzG2PfnSgwW+2+4HUD/VLjnlEHZfocQavjro5/
h6NIf+NRRPilxCQQsh2TgStAwZIw2jIx7xal3cvieVbHBodqKuimY/BkaKZZNvU/
w0vuaF/wp8K5mqkjSxTPNMDABkOn5Qq2/GOSd2bHR2nLGksfBVYnTlphjBtGsVAd
1I72qIHeFdjU1iwP5PaKYblt9m6oPFy0wWvncAkafveHsBrsqZ+g2ENVgH/FJLfl
19UeT1VecfAHhwRdzwi0yDlLu/Hxjsli7oEI5lvJfz/E9bYG7VaIcKvtT9SzSH6v
0ASv3bmYyeveTc5CaCF+51zFpnzMMiSpGVnBe+De8SLI+ziz+obSmwxyd//bH6Vo
hZtHL8Y1kyz0ad1ZI692U4FzyKWmHH7WuNb9nXenMKOdrp689CfAv+4KlPnYXxrU
vAnAhYRT3cXOyPYJh89YtvpC+EvqeXuI2lZT8YbpHgN6P4gpiE2d6DU2gbZu4Sui
7GnEvBj7vA1VKhWQbJFnEtF10O8l8zIIAVpdhvPGGU3BKAI8g+/GJbIHovj6ZgiP
Fq22KkdxcqKlRBjQKVhGwgroxuoZIYeZQuexQQxUmiJouRtLoyE3ZWauoKSXBpOF
Ev5dGgi0iXv8rfYpXMHRJFXkwi/cYTHnxtTm/7oAR+J0Pm7Vc/VNLmrsdv3LZ++o
bJlbruW4Xwd50RaihtBjmhuvNCR8F858H1tuUT+IyF0AgiqgayRNnIABZOGtymjH
Um82EQbMZ/fEvMmluRNyu+x05bPNlwdKD3V5M6IdAYQnMNNUdnltRGG5dUPayMsJ
NbqWYEfbrfmA5Sb8pRZ51hhhjiR/0V2ddzryHiWBajp4iWkup39rq6TsJVTxgWpZ
IKZ4mtOSVf/oURj+mwJp1J73areChT+/60mj2BuBnPu9/skQZ3KlsD97mRT3+lWc
f2osY2lvhadP7qRNjt9qt0X8RcBY0bOCkzPkS3YOygSdMDR2su44f5+kN9/SocV2
tRqtubQWUrFT1+Ov5y5DujTDXdqxS7B0Vv+M68IBGwhmdR6uPPM0QVKEybG26CZW
+3fYBKUN/89U5HfP5+LQI02NTDBuqCuuZhieI24DC37tgLmcTD/IR+J9us/eLZlz
8oZvcFd/U5gOvY+loqzUqB9XrhwkOcydtdq0RP3KgMMNp7MWtTToo6s3yZKNzBvr
kA4Y/hlK38VTfNO4owSVlSjApM+WVefayGf/ILXUsmy598G+x/eCCuCTaDeObFm8
6jwv7mskAaicJZ9s5G/WtNuQ3WIsge7WXyQlwPEmsT8V0NJW9OyeGwV0VNJQ3r8f
3tj2gunhX9IQivnNHiae4R+r/L3kirSTRmmcRT6MSOncaHsdgzYisE/qSmDu44TM
1kCLcMAnx6nCIU9kfMimXEe82x0UtZnFTkoaP/XgG67+8f2Y3WhVIdc8t1gIO8Ei
J5IG04oC1dObvbu/YZMstZPMNMp1JH6mgw3U/bE+srwtRZQX5Ryz5i3fNId/sCyy
19pPYfiiu1685ampKJDBr2dsLnwqAHOp205r7ZRUZct9nvjETycW2rSOYK/sEmTB
FnkAyGTjMtWPAqhhTG/YUkeaWIQUPLZZHkuepxCQdLphTROVuqumememFsGVZm25
aCDGckAvP7Mq4qbhs8cG13FIENWzikO7YFbSZ75T5uG53WU+uCldO2T9qCa63gNK
RZ30Lsn0LmHplpzUTtbQPTdbXLg2aSTP84VN6/TLeD5bHOLbSEeTxeugDPfDWQtk
hlMeePjHjNcfhtapv5Nices1oBFrAkg61jP4dSxbvu6AKUVQYxrNZUlZ3ggP+AlB
X7VlsnojQI8+viVhbViv0HvRcnSeSLwSk8J3ZfnDxt1xqIii6CiRhpJnRPmh7xzB
gxZSXvqRFBWgvVQmL5Vsws4aYpNYzzMRejCSp19yQOB1rueb6O0a4dUdH8hynmMi
eTr/ewK+DIjMqIJGZFoItOeEFK48MKhSQoUrOCm9OX/H5IyzxIyxaLsKCGFkH+/C
IomftAXftPZPh5U2kcIsCDwCksH+fKKT47qXD4mVB6hjvElHHAOHZhAwM9iqTW/u
Ol3wAad83Cdz4y4fUdfImLRXbZJ4DCxkAUHFdiL+DgWnFi5qrkdBrQZRZKJNlzx1
6fwKlJ5zFCrLqJuBhxQ+1Xf7+VXHx3K7ruqlcvLg3bXXawJNv/Uy7RyAxNms1UwC
frXw7tHlmwTqsL3FY1e/rnAhDG4PMtSmz60KXwF9peDE1kavSUsBtnZHWr8Pamby
Rl6E6RZ030bHZSTto2XC33usys4OBK0/lW8u/hTRIbhnRcyLQ9MnHmraQXGiXCS/
lUXIkf1/pAppfS5FBLDeQBvS9nVCi3YpCq8N0CfqG2JyFvXLD81GhWY1AfaY838m
KhVuMnN9LHTQdXjRZLwaTlMrDLNOun1ycmpKacYiReLBgHnQPZrWX+aDdCm9am94
1GfwNUbNljbPYPA/PM6ff+yxKaUN5jRcYWeXgs5WzEe7TF3Lr7ak5zV9Ew5VJU8I
Kkdt5OweQtq0iyYQfB9P50hLxoMdQCy1zPnYDFS5I08+qdepG4sFbbw4VmQuHtQ0
UR3VMuEIaJxK1ac7g5oDTZ/Vpa/7EnN8CnoL6xvUhtr6rowZ3a6wg90qKwvADKJY
pFB0nj1vgYXah2Qcn14wSoSMYY5Ry8PU6hV9+r+QC3+yBRlLenxt5VAfZtiFKO4s
m52Xsg9wuHR/hA9oy3UBKAj7On+x/PWmcpBfXXNUEigt6JgBtRBhrmx+Ue3OV+hr
GY4zZREL/ASTUEReTKpbt7sNOezHGiZnslo6P2rgJMgTxHE5nr8nqZ5L33M6Intb
3JBVHlVe1S8OyRtGa7p9Db3uCdRb2Q8w1d445ztHYjhkTlLTtSvRDae6VMulAVlj
S3vJUU3FAGuiZu9pNvTDQMKvZ6+91H7l5bvjDxPu/PjpOkgHVZ2kdvdMRSen0CvK
be3SunyENiP5VVFYty73LuXztCf0r/3MZ9ttkc6YK4ZKfeyTlP2wV0qTgd9s7Y1T
Yw/j1px3+JeaKeuq0haOHvP00jEAILk1Ji/sjJvrDxC1e7XPINKARejilqbEVFOE
ePOAPl4bHcOOUc9+i5YnOQBzjAvLIqmUaFiB4bmtQnahG/M/h+5RjUIfRGZF7JLz
58X4VkzwyHp/s4mG++BI4iJHZq46FWnmoOjT4uhNIdOUOPF7orJUUVlITNibb8aS
LHGb7BSEuB+C2m329gMXbmF4/KNwyI3hWP8huOYLuW88pIfphGJlGUFLxe2lfMAN
et9tPXKFvXIQ7a4wzJEthP+FW5rSG9VZ/NKBPzFA8aeGIfIXETxM3X9ZZXAWtNm7
azyOifHLxaK0Z1CwWPgmz4shackBvbxpfoEugpUSORrQni7I48ovhGyjMGVXGaWm
bfOs5/y4zg5VSiMvSKCrV0TLAksSYj3vniinA2OqQhFdzGA0H6ss8BjjTUiPNHpT
p4fDTsOEzuswNDbiAOBO33075dqu86SqnLiod9XwWym8oVvRTST71IiDZf552vMS
Z3+t81LlLhLMi9X5Cp5AE6zGQd+gm+bnhj9DjMHwbhu7KnGcrgw1f5nHzerANXWC
b4A6uX1ihj73pHso/7nrV9hoNfGNzJrVIOWyYfwu4k75eq9ub7CXwkx5y2PaXTQ5
Z6VtwuRICSdEafJptIrU1aoaMvNW2C7kM/YhBIa3E82xr1PTlwQI46AjmZ5C0/Vf
gDbvRBVoWqCX2SvuMofUr6biAUlt/7e7U/OqFlCY1L1ImgPzU6A5Wf/46M5q7x/i
6VNMtiJ/gZG/tUSZub9NB+B/OpF1i9LsVxn0Rk4Ar9DNahHXzpHVNx6iYwE4hK7p
ZiaapfBR3EL8nwsmvphaUwSBZdpnD7AAGr9N+zm3+gGskJKmTg/BRhLzAYoBRnXM
iCOn7Js1QbpSBVNci/PAO5dOANCjB23aFl/YTzTofHqsFR1rGWT920xTzjAv15UE
37T0dmFw+4afvjXLVTtlWUtydfIbdoTqAKLvkHFwyYImygKZ9U84Hb3DXKMsjJq4
pYKPHX/mnWkebGTKmv1qPUdbRjmsawrJp9liDNMDu4+yHskVacX9OjCU3Edj8iqf
hKPdyIhICi3WtvnYALimRDthfYlO/v+b34vt0uBlXRqTfsY9ibjI9Fk78ZMz5ADP
Sem6rk9nNMCqCyuFzChvzgLEAESrkBBsItbkz6+XpOyCtxJf6luWiitnE2TRpYXa
JE07oeQb+0gZPjRWNoqZxMRzPtufkDg5Q0qTi+CLFb4h8RdPas00j/B0kp7Ngubh
MuYSsA4b7xkgwxCIkDo0MYaN6Su1H/4U6Yz67EPCnNEBBfV9yhoqQX3xVBNEVQEN
d4zs//RCVrE7DCUL6lCk4C58eizNQTv3K+itrROOdMfRKOUclbwSmWvJO6Wa9MUz
wzBci8x2qoXf14+prx7e9UEdrce7jVIg6BBSZXsJA+dT8BVThybWW3bKCl/lR9tA
BDrZA92jWL+cmMuTPDTC/ZjVuYJaqXZxJpB/4U1UHEAA55art7Pc3F9MeoflPN38
bV5AHixy+BEn6lnaNIRCVz9GA5OYjlzom5DApScHbx7KFfs3mrAY27Wxa2HIbkQP
rLTX4D1k4H87zhDaMMZtYJZk9489Cc6Y2beMOPCxXEDbWsyIZJ5rkSAp3k1zi2Wm
l4/hIwH7b9WqM+TmBS367jUIXVDXjRhh2RjxuRQVSRi5yL2g4rGaaNMMZPYlNsW0
RsEz/aA7ZbS7DCOeeg9m6glKf7BCTkABrlSsX93rHMg97f1suqKYc33Pv/EPDg4Y
P+Mcqgxj6RwUzX1m5E34hPGV4RsmiTl64TBbtf7sKpme10xsFOe6t2I8O5mNu1dX
+GcfKO2SrcqIPfQMymMK1/xQ8xhWb2ZAJqy0LE/JN8w6AcORuNDmuzxEUqU80BIY
RgxGdoEHXuZ8AeQ7FsM8AwdCiNDa2kdk/A/B3LzXpk8h8o4bprxaa59ecHLxKn0w
HGnKEWB9eszdfjnLJCPiVbJuzytKRRNIxyzFTWDFVwY905aaz6XwbTdvPbwI6z+y
Oi+gQ0AXuSWemrgAoZl5XnFQwrDT403Bl5Viy76QX3twyd3VESLoNecTIM1ZHNFO
75ND5Zj9l8jvxTUs9JIR5/LX+uXyxydrp/xXpEp3lmJLKf/S3XoZZu+pFaXCiZKe
2bYZQTBqnmeQS7fP86apC5w5DkcswR4QLKCDfGnxoNvpIyCEzY5dQjiqEeK3mjY4
re36mMs1+GgY0gUgyANoU/dbsXcCyBU/zP2DOxsaExOy0D4wYWz8X+sR4ZGBWOvQ
irhHWctYRvZPIVIQBpOJFcHH/Vl3DJa+JdM5lAyvsfc4ijHtTpN/zKSFgZFirCzQ
iezyXBKLeaWSOmj7jrqToNO9AvAp/4Nxr90/g8aJuoBQz+JSAzUgu7JMo0aoTdwF
npkvHzzy0DPWnGmhphIjiAStDvqkUDR3mDTsHf2v2rxuXuzYo2vYsfpvPeJt2kr8
/srixoL3ZDlPFR5LfQPzo90/rWYQaBT5tMgPr3yEEsFd9Co3Jdodm2cqglsFYGt3
0z25Gma22QimbeDrdnwJdVtLCjx6iIzPvR5JUyCEddtHdtFodRb9q0WUlKX7ubN8
FQZIqF3xkCnZKXaCroYGBFGSgGI3prI8sa6e2hIn42bKmJgfoJrJlbk3J4cjN9dx
TFtRn4h0cxglVk2x08plXzqPoJFsGo7+g82s6OMcZbqvVT6Cz53qNmcEGdSsuCHT
egb6af6enZ7LK4pRvR+U+1hCLPnY7Iz4BrMqai+eUMD1Xi/4QEU9Edeima28lpRP
5B3RSir4q3u/HgPXS8NBYDH4dYWnzw/45jF/1iW0rFCpkQYe1+PCaOx0IYRXW6w4
HplbzdB3yMUt1T3f7ad4QWul1fBqEElvW4+jDVwoJG2BvQB+izFmRBgn/HzUbkVq
ka5Ej4Lyv7Pp3X6krlrRDwgKV0sZpclnFIzOyQ4xwTx462P/IMSLYdv43tuCxC5W
4C9d/XOQRMUgCpb89D/gTI2tBeTJ28dzKYfENWdmI4ywhKe2MtDkqYu8YjWaTnF3
mAu4YVYcUU/iime9azCKxFLTb/QAaTX4/45xYwkgJvj2n67e1qc0BrBrIbtESZfV
ss3jc0jZtAIrn+YfarFuVd4vCV07/wIbEFqvNuYzrWp499moDZA07PfYfdYsWikO
VZVFR7RU7Y9pptSN+lG7+BVY7UmsKfSfKE+dkcROjlXyBLxU4mp12asTcSqg5UvS
G0ERFJjZBYg7AckRETQUWa0Z5gausU/HpxdYi78263h5IimHq7hODGLB1LKCSHF5
diPMIr7MLQvMbxDk4nrrII+qAElDeIf8/phIe3/9wYy+gkZBUZ3jW4SfCuAgHn7L
X6juGPYgWdRU3t+NKsSnJuwKvRCsZuIX22ee/Y95/c20U0xLR4NDCgB1HhkCuZwM
I457CCgntYTYgA2j2mjs3xa8Zq/AA6vMlKXTyuizZcpzG2UD4paJKi5xatgpU4W7
wTO6OJs3lzzTHng8e6RZomn44IFV9PoJNCPYJv9T7l3VXgoHapc3EuhFtM0PKKfd
iECkHXaGm01yYHRRf78fOYPY8w4b4iCVUG/dUCzXBQd8ra8fRaqMbFFE+a9AkBfx
6PDBrVz7kgyYcSX/Ws65eTqwXKcPAIx9cfh1mod91QFtJoZhNOF90H4dqi664dMl
EulpF4k0oRU1TELDoisH3jf9G3iE9ssAvdhCESbKZZG4itVuHVUVXfIpAc9QCuSh
5Y35yF5rFnCowpQVFT945y45DUhDJXDVUaf7uMOVuEogzdRx9EL03TxMaJr3+3c6
+DEqhocfbkQ3VpC6WgC7PoFFJj6deIGy2DHs9DJPLZdbcvf8jbdiALQTjftVzZ/7
xUIsBMu9P5yGPhuQgsglsag2KwJw+bmB1+jTZ6Ktq3ZoyAq1phtQoyMziZA0V/ty
fIyigqQIvFHh6n8V2aaVCnswT8co4Ra3PN7COI5s1kazAdt+Au5BQHMqYr4SsQ77
OfYJWhFoNIaW8ha3mz7r849IrRbUQUOv7AdK9bZOqnGJzwfrgZMEe3W0C4D2Y6LS
Kg1VPxxMdJ1xyIp6ukSmz0LV+WXeKwAyDWZWPK5UiVjD0f7T6qoxlHA576iu8Uh+
eer3TyD+vyLHnnAaCyQzCnbUiCBD5OF/XMuvBDu3lgmnYG9feSCMux5Uz3MjX5z5
mCtEd7LMCrZFE+Qyg8BNUGQoagYjcfeDyK8XeitiGxWUI2Jiagitd25StK3tdIRf
iqPF7bYHJ97thwpE2DlfqD8WYaZoS1ZpfyANvwnton6ISmfHRgbeVI1M36TNIjvb
2tP6P6V3Yn24Zc6uhLbmmDWhNa9vXg6RYK7yNecAtobH2KzOk0hbd/M7DGuqjPDX
nExOomspqHN0GJ6bev+v90sI6lOoItJjBwYg9MDSeJxjpgXYmtLCWogVKZimkw+l
GO7XOQKZV/ZVp+TeHMWY+wWgkuqJfjqp3hFwx2Ea09BcCYNZCzDBIKViSzsbv53H
5PlwkXiNdnPjr56c3km0QxGQJzp9TsHoJwXyHHEzhzj0PvLumU/Gm8ciD99oFJEa
xXIqGQkEtqlf/PcgHPDnZIMfiUEkF/RVyeEGHt1ve2ameiRYUMCVZoBtcLxq8eI3
/nOVD2O1K7xUoJvWPN1708W+eCA+2W1vVOgnO9de5nmTA/V7pJiB/W7Hrh2ReQ4F
K6it7G1sljuKG1pkI9HYXceCYdVCQW3CbAGIApzYFxYeOL6lyPCeeco/3W4Ixjjl
Mfbw7Aff8Wbl8LWfNIYcOT+OwvZp2qrBiTjjAOePhyPXK2DCrOD8eRtavOMF6rcD
ZFW7H6tZdtXPtu3jHY1lBBaZFo4QvNeAkX4I/9NJLUMD4nJ0RxSJu67oXv7IVl95
2QDtPDoiciXeoy9h8kEjDPhvVjX+Osx6NWGH08bMgmwRO/1RNaxPGzphOkUNISjV
EYGEw98gXl7uePOJ78spv/0Sx7/3Lmo8U8Y5VREahzSKC4pZJsV84skm8X2MKfPe
M1/WblZq85fy9EKfuckKg2xSkOS8w9i3gvRtkkITlr41BC3Zbo6IjC3wqXIzvx7c
2pLlaneoEqyro25mbO7EK6pGo7X1i86YOenMmdLkUP0DbiNLEDB68k/k9CdxOiec
yNzpZUlSRv+XjQs8XIdBKkpJ3xvHdG9K/XVoKtDHiTUYOitop5nNZUG9edFCQIkg
Rjbu9X6sU9yzHa6PZiKCyqFDWxLuLVLH2jaUmH17Y5B7/gEasmCY+zCV8qXndyZp
Grrpt0WBCO2R4KiJbxdpNM1eUw6alj6jXN+WJ21aU7GQqCgi7Dalk8F8ixO5W2Nb
TVbJxGsGwEgEaXGGSXEngHdWWzg6htwh4CE1F/UHtdSGv7x7s9yFxGkG0ZBRuC0K
ExRHG86yRGLlNowBh2C89K+ayPbSYfZODK90V5Ll3JnD2s51EDf1yz88wVuSk3zz
lwQbBuDi162d0eHWxsO6q+nD1I7d5lwSax7lYO9nkwe/vt4yI1m6933yg3KmY+lR
pbRAN8KbEH+BpFCpRaV2B3Rm8UIHS+Axg+G/2izSAG6oyOaV99ACugMdFNdRM1d1
fgNlsMmarCd2ZWvWndEOo1UMWoRxb4V16zcK4bNC4jkchLQ7QVWrdO1bg/0vJIjm
wkQx8sG2KTmfxNV0c7lxYRWwDFZgK4NSjH3+del6vUyPUDT63OiaCh1HVLtwqZj6
e00yQCEa/Bn1xrqwO7ODJrpmmwx4RWRMNy4vNzzlOoAHnBBaGHONo8DkBGYfZshU
QIy4p4k6obtXb9K8XWMmY9TgPgzGrVnsH5yBF2dEFmHP+WLFRXD8cZkO8YuuGBkZ
/K53WxjM5q2oir7UYB4uVbDfjQSSG8jPm/tVnRDvx1K5aqtthm7vBNZe0rAwcou5
utj8v9ByUtC+n+9+99NxQYYjrhYxWbGeiBDG5wrYwjb3mBg/RD3qm2pJbaZVxD1d
YP643JvMwZchS8jqy8PVWAuWDwJNftg9WjLryC6TdkyX1KQIfBBCKGJL44nwkUoz
UNp/d1vRchUuEGFFtwvvtM2lFqXI6zVbn3aqWnFqFh8/eb5mNVWWaDAj4bXjccLd
5EYNGNIz4u+YGo1zlLchPr7pAVv0BlgeRMEQYmh6BQIv1rTDRxqBgedP56Hq8t49
pOnfTtrmVi27mJySttEmiOcsVzkjPYueUWhT8uXYlFIS0fGn1mErLoDlZVEqgt6A
V1UcYa84rXQxs6f7Fhf3ULFN4gxUITGXHYq/U98d56uxxs3bWwlGfTdJkN9VBy3O
IoXxs8QwgnZNmKAAqWF0wnzSO+a0Tvu2N8I7GmzU+cBqkJf7iinuLyi64CKN5/yu
/Yi9LRHgPePNYEoNgbmCSxnYoGReOO1FVtXfu/pjaXbGFumKmuLVckWDFFiZKIts
D/ZRJOAe+DXOGSupZwx+ZGhrC2/I5IUeTJ0ijZWl3ef0HyLqTR6taCKXuZ+BUENY
BmGiP/znQcglvahVRob+8qRywgwrqrVoPEIR+KMpEw+Fx7+HNHi/aZxplIai3qYq
xPqd0gC4mne71IDT/P2lPDu6+YLU6MDjat07vlYZnmDDm1A5jwqDANjyGAuKZCOk
JiXJLnNth3qAGLjeMYeeGFcmSWLIyJVjo/eCD/3wGJ4jHrJiQ61GZckF4WF/8oXw
dnrRNXA0YEj0gmIE+VypjqhSTioLBRBu34L0nfkrvCKhemCgreF5ntvuWz788QW+
Qri26R8589S8JmTHfkVbhLAvI6Kyx6YPeuu6l5FxtfFVY/HQ/xiJG0KarcKBMy7k
m6Fp1wQGbyjUgHelaB3hCSdzlK+17YFi7SqAOeQEZ9cJv03T127S4Hmd8Zjm3OGR
lc+pcUQ/SlnEQVa3gNeCXJqqEMGEl46G4CPV/9qOGfDNjGlnVmnLeWWMTcdxnT+h
RCLycMsRMaFUm9+zPxYpipolUx8IGTsUj5wjWNxLEiYyHjxANsqDx8VcNRFKqpIG
YxaWxtiFr6aSPZOmRjRMhuCRCP5UbE4nC/NQ83ABSREtQ362S17qxVP40SE/a98K
OvZl9RVi1wSH22skFVGdlC5fGaC9ytT8KFwSQ2YfSaHSH1+1AX3vkYYldnvxfaVf
rUyp4lEy2yPlbh93Xvos2DXH2o7LHS/xyEnDzBqOUZNfLi7MbmOxXFpCzYwojyEH
N1KoyMWStt0LYPTT1Syt18yICdm+PaeHJvh7ztAZG3cXlMd4exsK+IGMVnx+q8Z6
HA1ntNcaAVusyd07RMHb7MH5KKsHqht1Bj5sO1IvhpWy3+10ohsS88JShnfQfzFS
uyR+3iiROh3K15IQkpgkbpQG8ErOANpnoCOWMcuGv+E3Gurhbp/82pCSWbtKAAXX
gZv4mECY5gCPOdJnA2mGnLEcvxidaHWi0NSOVGl/t34cTHq0E2ZvwXcYHUCd+nkJ
e9Zagvhf7mLB0t6hK0Ao+fezFAXbcZ2mZhVJq4riBc0M2MlZwWMUtH+no7O8AmGH
+nAsEKdZ2yg1EIKQb6Q2YaaNZWC/8R4MhpkEA7SgPPcumbswsc60QmNsixgDlYPR
/H0EnZE8yuvqAMLabppSfLV9VaPzCWmIHYZXERFg0Jo9bwlUAZXclXxa+LYOBOKd
+hY2BGFKghYRZ0UjWSoswiVY8RyCs8guM/TVhsXXRP+rJ/n2/J+o4xCM1EhabDUr
33lfZS8tVdiYrHJdqnn5HT06MaKIYJvJic5fT/0DjorqmG3HiYEoOmARJD2Eubwt
hQ7yj7QK/K4iZG65Cvr2RYXuU9oDn3d9FqHkT8suF1eGLJmXkNrLDUCPKmcd0Riv
r+yi7mxrbgK0zs+QZWMqpv94OCFRFFxZeeKGC4VSd7a2Dt+deNfaVny9ELyRgSGU
g9VTleyJdGVLmHMlHG2wNp2Y7ajBQOFJEyatCaJj1fNPNCQpzFSUK2suPhVzP5NE
Yr9PLHSPIYQPMWa9oYCWt7hRepGCeo2MZQ5gud0SkzQJKFKkN1bIEU9xaRvUgBg/
21j0l/a8YyRvegh9ZL6nnfzJj5ScADVbUU2HHi2rPXpL3BByfwL4b0GoSfAZcfk/
4o7Xvp4b7FBc4ZrxmUMWMQJq3fBoZYlABb+Bg7kZER+Z8JiI/+hYQ3IofYo+SdMc
6CxWqcqp3OOutf4eb70cB0ehCswVk/Pux+DJNFK9nyNRQxLzF82618ez+juSXB9w
Wa75NulKbCicAHOFZt+5oW3uboVE+qNMFpugMhNEMl7Zp2h1kRm0ClYQuUspOVWm
mNeIUCNQNBTb8pzpL8ffcFlTWWcYJ1KnNj1T4Q5QuZvEk1wPINyE7iKxqNiPoamy
VuseI4YCxXiGdg7xJJtDjDVkAsKcUUD6/+Nk4d3lfvQ6xibo2YY9vyS/4JPDi1Ye
rbg3njOxCYiycF+241Q1Cv+aQKggEZyfqzpXre72N/Ucw0omXAEcPOroHFzrMOjW
wkJrYcZsxwyO5RzDfIa1SIsrdDNnNdU2jnxZQ8LTpY+by1+vAbQm2+HNFZcF6r1O
Y8a+PiVPjAAyyJ86Tp5JNLMKsQFkxgzX1CWQKY9OGdBwvC44n1dX42rW31Vxbzbb
yVLKJxY2KFfw1lOXefLdy2nEe7jnJe3+Wv6z7BXwV8IFtFbjtviKimGzN21D4hVq
oh/S2IUk1Y0WAlRE5cZlpZOHgsLDBiSZx8+kp4gkQul6A2g8ERhwQX4k4+GtkiUF
3hgBH90/msfVPCGjFUEIlSKHcCGot0zOnGID+Z9D6GWcwUuRexb93glq7uresXx6
X/dG1d+j9ntVWQxeeM6Ea+YeNmQNHAkfn4sicO5x10soSBrc3biNwW/ZiWzV/w76
1i6l49WNhpQmvlMz1K1MYWaszyX/IggLCoL2K21gijuohuB6Tlh/Zxqj8fsO1cOc
FUan2eysVHpRj8zXVfeboWOW4jAlfLRcECv8DapH7fOlEEnQMznywnswsRQwYBIv
e9p/aY4Ym/UTLYShJ5sHKMuCLszJKrIsVV/AUkKMY5kM/OxN5DAqWQ+ptQInDvOg
nAm0rCZe4tSMr4i8NL4MRkoJdnXkmjV5yTuYV0GKysJQM0bW1qeQLyavXz7yRccb
kswLd4rCUSKA02Uib9Ez6sy63qg3W8CmLDJv2cS4R/CxmQLq7rK3veVP4jzcIzJJ
qxfsF8bnhIYf8M1k624zb3tx4xqUFUHzfgZsFrCpZ9z0eo6mDg2AWG4bQZBINwo8
SNLGX0wjabHW7JAvS6YpBGMVogcxTA88/nnP8/XzmmMHf2wTWtwCrICNWdsH5a3q
nuHND3LacMPxkwWf+lL4ucFTmLlyeuPW8SPvou992Sw5m2EWixkFhTFhCpn6Uufb
0B6JYSc1ibKyloZcVQ2WBdExPrMFZ4bTbi/YgD9CbzXJY+hYllZeHgGSnDkNfuDN
B9jOw55jLyGBuMNqxZL/hVeyaE9d3t0HtY1xuead80dt5qOrXS3voJWiu5Kzgpy1
G+3mjxsRblDHG/PKl4SZ9Gi94YuK3f8sjonTSiRaSdA+E2lEmm25ZG3cW7x9iYSp
2Mgi2ChxUihQ4+7Gm4Fn6jkBy9V9ynzU/H/iQREH6m/mhSlktRpHN8+693X7pNTh
oao0E3U7TMULiCybTw5IqqeYhJw8nLHhmkzGHK/q0azzpbL4aR2zX1YvOivzA9wH
SWBrsKQDlpeWG+FJjAN2vlA1pc9GY/KGD6usihQIUqFCzd288p+9t+df4GP04mwq
c/1ev/7KIEu+iELla8x/z/aHByud0VzymPKAcFiqvvoTVFz00k2XJgYt9dR1fbWU
fR0gLkzdPtU9DHOCuTeRtHKt7AOMbnCFCKrbOlMN9g1W+SWE90NEVHuwE/R6KzYr
jGE5KfUg5F5B76xjqBI++OLjr7H6rxsDwsFauWPVJEIF8+Gorn0RPuX9MVthiUnw
Vcjx7omImpRfX9tUNiywcwf6cwnj/DU00gtbRuZwDcCZiBWDbkYpegutFp/KTeAz
JNG90PwPOUX0RTz9SyMGL2KUMMOckQX3NuMyRuXI9UMK98Y2tWWh5ey345K3YW37
yjrkjzDQ+IzTExz2k9JtstyMyBWhmRrlsioszBPtKPjqVPyVD5fGuHDkCtDFEvbS
6rfzVzLGjhc0jim9qqNBJlHaIo1elOqHi6+jAE8kX8/pJOF3Xtlw4mK8P+K6R0BM
rKu+D0azTmALfeK2VpCzTF+lKReOW5Ed7ISao7dHvjTAeobBRZXUPwLlMQaQEiYP
WaG6H0CvL8cJALhnpY+KfNOsKXE9r/CYl/iXKZrNmK0rSddpCYUb+fOsjlO11OCd
r3r1xo9wN7BsUWKHTrV6PU2K4OkHw3Wq6pFenJJo5eQy/be/hTVKWZgvz9HsS3sJ
ru2DiDwHKBEOXGBFUGRIjcTBIDIKkA6ybvdbCuakD8+X5pohR/eVkRh2xQWbZt10
7J86PCO/C0l3DOB2TUWSMhB2aq/UcGFknVAcIgW1P7SpBSeWMLnZr+zPNGFhGnYu
o/ZWuxyQhB3zJMbHxx+wtjpFKWE/UJAoh9JLmUWgPsLP5egRzYqbu/PbCEuT+z34
mu4SIoNlCSOBvAYPYRrPvKveCGb42v+LBpuoG/3AdYK9EfGLXPJdFwVFohUGy6Fw
9YELUe7eG/sJQxQJN2ooPzG/4rDUnrergyJ9JC6LJa2jFlhX/LvOlL+IOkUoGpFo
GOgJ6BHFu5vyLB+yhgETUKhg2yD1dQE7ZdegaXwH21HRVwQ/+A/jBlfeJ7gzJGO/
igUSNJ724SXlDMVQgv7jHaDgCMs37d2K078pC+6NtRUkgv2AQyF+5V5B2ctmhTpe
1m8QHKNrEJtEvdKLkqkVhOMWKZ1KRDpCDqMhC4iZ987Mcw4ph0Ln8zsnEbUkMFqS
Op8B1swHf9rt/c7oRXnHfa07VrHi0XZCGXvPhAz1DRY2onCmVDJMdohuIFNH4d/3
fQxtjb17knHs0mVsyRo10I7UomYFX3qaXacqwsHW/6Q6/qfm/Bc61RgkLpIERJM6
ZRs6b0BHXVbfqC93HJkwHpyIuzOcgRhsuri07nfzD5MzsHC+QofNknQaiSVQfZVU
glw8zguvcni63G0XnTQNfr10MzqSiSsiyCTSc10h1QbiXQDWcXIsyRYKqs1x9qe0
0tor6wNAW5qVki3L+50euWJ64wAoiTmu3Wo0TZ0/RsHkk0fbAQGCnNogRMG0fUn+
JBYLw+3ZoTOWWUMt3wxD8Mj4gVomf7eaLqUu2cw6EXAWurVMr2DEKTnmvyjE1Ujl
ZdKeroqCrM/uo67WbuupTjVsFbXa+8WfVI4clc+LCeRzdBT0CRAlFfOs1yZN8E+7
lfY90kNJXc8oI3mkokBOWvFpKoKXjEtLyp33GAdDpdHwNIL+cbPAqwPER/126IZj
4atXG8HIqaGZbVkpbrWCgLmqLjq6nniE0ng+OA2tPbHQn2mipJDBMLK8kTFoUrqY
tbU8VbVHFEr0Fxbg72I6i5e9L5S7TP0/wwiJTAlF5JTxn9z0iipnkxB8gYAF5eQ4
pyb7EdUk10essbHZLsAXOtrdoYA22fLd13rEIG2SAH6j3fBymByu5D6+e35IoSB1
gMOCykEgjxbh3stBVVCMp4KP2ytNKFjBo/I0VzjHY9BQy2dG4LlAqyAnqkBcpdyP
Pu+P39+lPWQW/kFRvEYPBNVTMjWttbWj8pxQ6dMuYsmVy8yZX49gqaTh3m0U8ds0
qI4W+bON8tLIXx49oeeQA4AlwonSOq8UrJVnaJhxCQZfJwnSuBor0NX2AS8m6Gkr
Q7kxr+7lL/0FDDRaBf5TYd+oPt4fWHwM/zA7Sb3RZfslwA/wvOn8gbn3BZzhNG/2
J0cgWBNpSapHwLZCLHrfz/5+qwaIBWw0S2a57fsnxUR/Q8cJ52aVAwzQsasAGAom
D21HFE9tv0vaa8fOEYNriVxCiMmn/+ysDNbwZ8SsbK5yBjJhNq8IjU0RmssFx80V
fOFR4cxe+80PwX3XN9pjrXmtAWRM8CU9tZas81wLayr2R7BKPNXNsUoMQ49njGDw
elW4srXd48vCZ31KL6ZmrFH+MpgX4wrA64JIychy96qN05GwxnJmWJ/v2pC4LeDb
Zq7OMFS73DXmIpuvpg4IlAc+FKMYjWcfxjtWCzV85sEYSF1QKQDPyiUNANkGmFze
AhXp6Tg7AgFbKH0wQSGvJXgx/GhRDzWoYWx6fW49OelXV59EnqtB440Cl+jVaRuq
X2GE+7Mu041KDVeQgdqIXy4iWZA9s1dmjotDgCRzE4NZ/FqDz4zMaaDQOEvIIJdu
VpofE1LxOedQjDm/dKiHOvps5UgFT1UoMVp0TwntH0KzDhZNCn0SnANeNG3xej4E
XHncNn1T4kJS5zuyExPrtStTTIyxn/ThYhCPO85zWWX4YZtP8EtdOhkGPH5t3MXK
r7QfLq9uqzc9bvxnnKoOJRB4gQwGRJ+tAGICemvoUB+yzyll0p2MQN1DdJcd69Zz
3AbnY2QmOlDfxljwmk4z8uiQvoJHpuXnoAwuj8yrS0CEKv1fsjBww6HjHjGpkBiq
TmV4yJA2sRrsve6/vrmD9lCqicibzC/zb6SW/qbvYpq7jGDB7u/y/bxoyNFS7uv+
eJWMHc224hJFt9iUPYFMuEfqLQs6lQj6j1WQQS8XLO+N2s6B2j6PU4g8Jg08Ee84
RecqjOaKyXP6v62W38pEU7BDyLpLZlZxa0ZDM3s3h3e+vMfO9Ks3pihUIcOEClHa
iVuPlWXRB/WD8GeIKjD7JblvfMlUmeyK4bzJewf84wF+CCaESecvqkTzmkUivrMC
ETZ6miNeCQmqZh+nEYKXmstpXhOkomcMCoJ9PBbfYas37n+hSxmrMRqRAE6tuZFx
0RQdDb1+XVn8LVbRegIHDlBptDSkf6SMYc/mBdOaIoAUYgIgaO58dDAuA8POyDeF
XKeM0aA2+RQzBovC/Sam1q2fperXJcyGAi8iMSZZkjcevvkP6IFCE0gL7mq47SV7
scheC2r7FhMPwgwZgjoIP9fo96lDCJGEF7BaaibV2YjDF/plPGsSyUo9lzpobhTb
d12G3lYICjezIzEywYeNNg0Z/NP56ydNN7VHI6up8XpIzxxAFlfLcjrrTXh6w/Qk
NBr9t4GtDOCitXyRNbGNAExw1W2a8dw9ElSRoK8hMkE8knXMlJgwoOUxVb/4L2L8
D3FkREKSlIj72M0MRZooJ9M5TioWL8o7i3qgCNc0g74mdWLiQVYsJD5GhaEq3BwB
w8+sHND2vSCwfMe22st/d75iM2n7ZxecRmrerSyLzoRohZfB6lLFNKrT58nfgH9L
7t7mWFs5eYZAfRr90cBHdErKbePx0iLarGcHOk0AcFkYHimTOu8+adqfeRhfQfbp
SvfLwD0U947hB7cuYqVPqp2b8KuJ6KTlJV6Kg+2aJrPry6cSFVRKfmkNmtec0UJA
2gTUHhHwfUUf9qXgVIxa3MRzuWIt6PiSnZCQENK+lhNQiQrdw3r7Fe1TR3UKxNqv
jsbMoHB125jgZ325ad0YNjP5Bay8aNrTd2y5b7R51XPX0Y+lPS8tWUc9+lrenFY4
WrZWMiOnZ1h4yTDnUyrd6aVKm7P9fCVjfQIwgu/mf0YWNAg3nEuzUlrDMfTefIjo
IGEcTt2xZru1KjHeVKD1IG4AQ4HwpoytuvbKojbR4bkja+d3f1tvaX/g9aZO76rF
PO7Xg1WHYUSlkrLVpi34VkGE1LpQjjVfzfznD10wdAS1pPEQso5orFALQPoVF+/k
N3EYCjjfGX4OZEpnYi3Xy/iXBWfU6TqTnZZfEg/19eHtvljr/D40xCDZWhZ5qY09
SevyyHH+h7599SmNK2HwxeDQYq6b0LrLv9T18KXfMG+FTeleFXPYf3SR0uNUHW8l
ysRuAO8OEfN7NXEGWzrb4ovHzXjsy/jtFI6sV4jDHH5/IiKsdfyyHFCVyswPAvIK
AFkGv2eevvFLkpUCYCpnVHPVLMJJXdomc78nKAQCsXUBMZ628zyrbualuWfjqCJx
hamyjkipF3T0CmQ1GGmnOVhKsFXWpMVPG8YuhYLitfEf3tHAYTfeIIaECYpyh6Q3
219icjrWdkWuQCfp/P781Vu/JpKyUG2QXBHzeW25Qmma/x6LP+TPqw5JkgucFDEL
l4PnoOqQxtZaOuLQWFyz8FLMSS7RfbHSN18ssoyhK9AnC1arrx6zECmmPqJmTU2f
LHIoZoM/8ug859BCVw7m6Z2aPXU2+fsCvbHsj4+AWLj+r5kiK3pxjNv5s02pZIsN
7UsR7VrtgR7DdKoQqjivXZ1okFRhmerhjZMJcgTzPROIG878t8eUlHkSWGMvLmgK
iwUwWqtT84/i/L2JOeeM3EBS5G+sLjBDPdh/e6XoCtqDpfbFw8pL8DpdMf3yOCfl
PwKB965jA6xNG1wB9MqGI8vK6eVdud7I/gSugDtYflwtR/JLgGktcRfr0umMJJ0S
Ky94xNPqnxm+VZzjGD4uzRS7WZ6a43e7WTFgEKKqXLQktVp+Fj8h7fcQfYgXEMnI
B1cqcJHc08SYVjaDWsSo6iBqiZ3BQDeznEFlWdilfgNYADorwyb9NC61DqYxzvEK
tRMUoJ/H1tPCEyFnsJOvJd049W+1qPPo33LDupouZrvmKfXuafSRkzCzPGVQyNjn
m8J8XeFiH2+YxIplHO/N7evs6/S1W1E2bbsu1DJcJF2N+3LoCohRate+drW0qftw
XnW5PTW1NFCfN5ZZB6CoTCmcm5sMViziqFsujQ+1+gstfXvINraXD/HrVN2GPIF4
4SqcrdYpCAQNxDESLJSmU8SyQQH4g1xDBWANb4Y1jY2xsFKRVC04MNqHmvgNglcL
SktowWWfVA4bOZ5otGm2RI9iHORTIppqwe//+QkkJCizN51AI5ICz8ttTOqKTVBh
NYKfGOU/O7YDOVn7HL259JSzLbXizRidKnUHQ8F45F8YPcLEhroj5TrRshQMOi97
7cRgswBMWju0BJV/ZJpr5YpBkRsYzbeUByKnkDKcU5YHpaM4PmdS/S8nYq5wQS4c
Z1p6EGUWrqz84quX5VnjLUgcd0LvQn3ABGpHxXQZ+aPPioKu3j5/lmfJwAfHwkTL
nMO6zhBKqoDgUZC92alF6NUYif7+NAbD3MFbCLlzffbWQgBHqw/4NE6++l7lnf68
PNKgUrayj7GLApJY1sjf214yMaCmAjUw/atkM2nWojdiGzCp7jYt16eV66S3NmUv
+XO4UpTrNbooo/vqnbu6fTNCLNdn1rjpaNX7pmMm24l70UGKHIWAXhf3qLurGPHU
fE+FsOg4YT9dbFnwuLxeO1e/sctpNIF0k20BcXouffc18mPD9aP9FOwd5VYyx5z1
sq5Gq9JYmz3GctvVo5sZ0+/ekU23RSr8uB5M0zitCh9Bclc8oko0cFPjIEktWpYz
lAsaTRV7fn02Vgb7V3UKut7cJWmT2pZDitfWUltrmvoWghZlr61GeVmAx0m+CDpI
V1o0WZIlQ5tpWwGBF13S7DmeYPDzrZLRowQJ9m11EwZmTtTZFrOPTiVqhYLOt2mw
J2aMFyRXSJvojMQP47GBw99u31dDC74hTUolqcyBZGM2Pvea2otQXPb1wi8OE53Z
0hxA3c4sACJOVKWJkOWPk7MBRMYgPnHtOhGX6/aG2ikM/Al2pyXefpe1MwkSVF4c
QsbjcbsWQ8zSGGMDheQcCCYHxd8Ez/VKx0bG5JJh0sIRrZcUOTLiI5LE2NRmn0nq
8gLItG1XtxRLOxlcLVviyr+uJVJr+khdwmj6ta83JMcD7eUFcdYvB/frAK5lEDMh
Bqr+ZHnl4MklFnhsGoP+p6lBzPZBs9bi7d9XEJQC1cKXWReQ+J7uBR3hXhE6Asg3
YyoDoNUi8wth0suySUDLjF+/yUOyY8Vfv4i4rtKMR3qN3dODESgdPdYFK3DS3j9q
hBClI/pdgJexuoDgo44WNr6dTjA09pi7s3PfSVWdrL//tMrw7IN/65Gvp5C0gAox
KHOvM7MyoYnQw5SBurcH5yHVrcykgdGtnXaM5FemYsZOlCQdMSNzUixQ60ysEbjd
OjINYl/ScsWHkB+Wng2lqJGGg6MRWCe11JHq5tdB9sF0OeTqy6i0uBHpKiOf+prw
zRhPw8+wafCyeyI36gFEQ2aToOxxSOsZcnOG9XuuXQV8uOpaVkGF/1rOHSR8TKxF
/YXkO1KFlym6pbuzJ+dntlzxkmqWHFUWUTFD40/JngyCKp9ZIy+FQKUfkctZeW2R
hhaAIK16/Q5FAyDp1Y9BC2GqzSuW3u8RyWYdHHJY/QvUKgKXhdwR+TILtev4UaEP
InAwTieKAqeO43FOxGnagWtB4+8f4HI8KpCShOh7lP0VhJQtXXEWu2NB3Q7pt1na
cAU6uG9lVZ0m3KlxrgxZNwbBMhDFS/eFiG1uPIdsjgNvl2U0zpDa7SVBIQc59IjV
9hODdbKuy/BzkdWh5QjsNq8J/BhvaZpv43pubQU8PEP7um3SXYdnQGRMjhyThwPm
SnvmtJNjTJGpGgDCmnL1JjWOzfwCFKfrOJjZq1grdDBtrA1OeVKswdM3Lpk9oMZs
7X6RgMYnN0RV20vxHOETgwUVE7tY6R2U7l4vYKp59WDAOywGr+A8YI5mMlqhK2fE
fxO1uo3t8anFVIqXS8k36Z5LapiG0WoS2ySfKNAkyEacAKaTrH5/Wxt1jRZUEFaA
ssoowppkSwUBs8R1pTs84nuurgifSo0MDt4fkqJKqZbWjjEnLz/Aj7mEKRK1NYzx
LFtkJEjEukTggluStVaeoJyj7eueRjxa+MMkq8uM4TQ+zZrWM4rI3ZosTTBsr6Tb
ig576R6SVKc2v/VkYNiuXUSNiHNQ/ttsCBlKGyrOfjNOiBYs0E6XqqL2jGQoK/ql
Z1SvYfwkUQWo0/0F5sMOceOPDVoJP2aXo0wjmszkdn8X9283+P+oFKviltlnKo7h
Iohw2vds8lKb4Tb+CKDMlDgri+sJ9oYY6LjsIWekbcPlFr/mdDXhl2TYcsMIwYxZ
5Q+mi7WnIvLz0MWOePU6pIRbbeQ8JFjpDGIeuBKlbz9uoWVk9qHKWBf0tNPNZN3m
zVnPis/sCmgbAt2Gxxs9E1xjxqAJ47NWlu7ToGAEU1Ikq+dsBHG7H3wyBe1zqjfE
fS5kh3TjKm54KRt1PAbBUByxM0pwK6C5zyZS6heIkCpb0Xmch/rvc49oh5phE51d
zWYpLlIsYTq+krYixJBnarFRvbvMGfjAx60cKm0EMxubR117lIYmvBBnXA8NTMJv
iiGmbirXGiTTFL+2oTmt6N+5LsIGd2fs/4ZAnBP6v4AYqSg3i7Qdf3L+3/uCEGUW
rhcKHh4ir64cbx/iP2tVYY2RN1JTMRsPUvFb9rON5AO1AxGvJ/Vlb+r7lA4Y9Q2Z
t0aN37PxSajCdIAb1iInhDzhVnE6xG72LDReMZkLMG8Je3QhIJ7TzlvQXe0kyRTa
gvcNZz30wniFqbyVT7O+z54wiOQg02VgZ8E/YjwBYSc6mFQVBcbh7ewhVGAdTrW8
WDRGc9cos5aD0KBHay0ue1F6tzZo3CKlgEsVXzG2i+uW9gvw3alxQECCnPrWyud4
tqmi0rVkFYOAGqjppn69GAepsXaaDqbP2+TQk5ttTio+OnuDW42wPWxx84JBdcm9
ClDJquQbyrrGt2DFzmRdVKAabTWywQh+YhO7mppptpzh7ZNll/+t/kl89J9ywc5Z
73TjEvqqyfHGcnVLod2ICq23NC8OZVmtR2vi4Nya4X+MqxxfXPvUJ8aU4/5FOLKN
8Z4O9oHpRPRDLTZ7w8W4XxKPNP19Wsqw4NouKTD6PWXAa2SRDDy1hNtmeV9b7dhc
Jx7UIJuG9/+zpMmSHFH2/1FIX4iSZMfAo+kneX9g2YWW29KinGOpghuZuy0oXWG2
DsHI71j3coNICeR6rQ1NvRjKfhar3Q5Il0gSdUuEeM/XK8CqNl8d4VU0IwOvFZsc
l8sskzU5FzaMrHLhTtn4Ily6YqJ+9sSa9swcdQLMScal2LRVKXpE/nwIiWpXb/ZD
1mCYAjtIOHbuB8E/NKuDj5n+7MFcK2/ZH2sJh+eAuH0TS+rlIBvCMqifdLtlSjh8
CB9fto9d3EcHdxK8FmJg7NTI7V+7LYEClOrKZKbz0G3wjCa/xEPNrngTwq/IkNiZ
RE7qHit6dykuZcr2K2wHyTbeH8B3Am94hGKfRbAxyedJ6yQ7mIyfMnC7tJ8d9grj
grh+GWLhf4avo75wnvwIlBWPJuoQrfZUhBuq0KZsjsIQQidRnoJvAnuMfQ+bIt0D
0acWlb+tIgiAXkvNA+Lg4nys5ARy+zrntHuGvpWTx1VGC+9ciUjZCpIvw+ZqSV0B
1oHnLC4+dsg+ueaXkVizIL6f38jq9PJspdYgIcqh0Z9Q8cglGvGgdmXu1UOuZpiv
EjhoKbe/HgL0i3qQGT4W/iYRpKJVh+rEYwQAf05+gGTVsBYvfTaCs9YX/wflOGKX
7fIrI8h25l2WYF7pc94CG3zG+K66mL1fLQLa3VGe6VcBq+R6edDJ38ENzXIq0RUr
bIVk5uV1k5725kuWaww4t/dDfQ07zcR740KWnAN/iMNlVmnwVg7jWGLRB5XDbHnN
OmF4IQEWNNnw8qsRoTBJZcaFlIpSyEJn4EDiAvmaH1SKXXFj/Rmf1o4U1dKth2Da
n7PEgUwVS++4BMZoRia6Cjwk6UdISLbrK3cV3FbPumTrQoEntehqa1UGbZaKejv7
K0Cnrg75FpoIjgcmGedxHE0bQ2sCLwiR7XVEi9ocx5o2ED6GYSLecQi7c4FCdsZa
rWq5UKgIfqBzkhN7mbm70wYueMKjpEi9e6KFOr/oFeJEXxcgQi89znnEa0Ytmlve
9SpywTUhvAT4OOnSfESmNnlh4sl6wLqAl0I9ScJjk70vEI4sM+EXAk3JJ2uixz0J
v3TsS96JlP4A/pTqq+9s1IED+ho9tM1gm0xHctwNuqYJxjTMT3CLWQX7h+9z1led
mNkoZZ5nCHXn1XkuHz5EqMSUfG4ciXpTO4CFcblcywxk3So0VYh4uAC7XzwIAjOz
VUEzpxqLETd4Vy6BrlFH/pyMVHTVIXx4BLG9VRtfaAn0qsmi2HQHD3FGQSUSpk11
WgAhjkb/7AcHxnnndH2iod4OYKsIVFeM8EKbpFnU4VNa11fKCXcoigWynpF7Ek4P
tXnWLf0sDc865WmZZMAyTq5ufMZpnJioajma5ONwjhYvtfSE4A+5kGZohMMays3/
8DDsqiz4JrCm9dVHDGcQxCWfz16W1Qso+3nDpJDZSjdbOWclFZBce9BsCm212xwq
wGXNAR3/9RS/t9Z91vmhrvh2tQQk//ukwZoYlbe0PqYj8w4SA+aqoOoRSpawCTy4
nwNXmPfU2qcal9oEQL5kdQHxaJxbJLpnfpDNhARGduobjcWmrFfTw55h8Fa8NuYn
YEhdXYFE0h+UA5gvnRCqAwNlSR8sEasSLeGkcQNjhKhHPgPVjgDaBoxh0xXtGfTN
oDSMTJASNF2laO/HUK4Ymqvicmraz2eslB6CXhZ0wCoEjFllQJsB2qnT7F90lxsR
sI1F5yVesZurqTNstdwVLx1YpSJ+Q6dYcOmoPhRgzsryFGBjBUpUDeEgFHwSDR4/
g2O02ZeUzh+US2s7d3Cy4SXgb8u0SRa7rRnIHCb1DGn+1j7p/Y5cOniYUXD3iU1s
MNM7mqh3o7YFp7XH+4+XiflUcmON/9iudIHGlkwERAQxojJc99BQcVm+hAtvCOni
7equdziiouqpa2x7md86vQgU9OrI6916q/m6XDm08jH/QgiUpiuKLfQ8uSOQYm+H
pLaJYKebxh7mkcs+9FPKwdCvptGf0Ybf2bI1GpY804V+zDC2YYoMrI38jKfApUba
tEYTptftDLv7CZuQFM5pZpa2TRgUodftS7vv5aZypSgiFSvF8+CQAHc3+g5VDThD
Rnkmz6DwZ4BlWiS6v52c51YFWMuQto9OiyObl4Fq3Nxsl15NDThob5d/jkAu9JxB
D7HLtKZRejoipbB6gmG2QX9n9UDmHJHeBu6Sq9AhWFPT+kOaIE9rgIFxG4nEy5Kg
r8Rg+BtR3XQbmZSL3AquahvR6P3Qk6wLnTbiAV5lqZk0oO/lQ3dFBl4tmePgZ81W
mbl3iqelYOtgQi3pzSm+5Th4lFu2rAIgmcz4q3Ee/S/ZWdJLFPL0bl2AXZ2rIk/y
LUdQdDaYcF1m4uGB+GWI2X3WoNOgmKNpwg2DDETr1Dq7+fPiY94jVjw4uKqvqQOt
xbLu771tPqMmanhIij9KPY0GF1y+OzASPznM/wQ5yRsOaoPooiqzt+r/veW3bj07
2FbgBoKdsKgdEoGgZ25roMKu8rdi+219wl2FY8CEcnfEMuNHp7k17VQF9EMU+6VG
usUP3ftiDuRbmk00iJ/bx5BzZgb0CTUr2PWmWFXjKS1YYpaECyzF9ZJShnyZ0p3X
d8ukdQ/1w0D+jX5LgcrKsHZVKyUZTi9ybsz/E/BpXWhumxAUmSbJj9DBzJxL4kcr
KROjBqA3qt2ZSj/fhPIIVitDQObeeqNpHkFVKquvyxS7MMK9Rpe8Z73Je8f600mc
uieUTSJE2/8QuqK45gA1bkYctc7puW1XJAOhMAlj1hBeERiByNN5th/srUhThtPx
/3GYkkL8NvwiKmbp2oE32pDRoU9XqebYp6ZosBPxJVtfK3JYZ9J6/OD237hpivIK
s5Hcl6+oOH2bAjcuC7wLuSNHOhjj1M+eDFufmxWKTMIqO+jZAkIVxZjZhwi7c43M
ZdOazX4MSZ7LkpxlEwSl4M+G2GShd+9prbfxi+k3lU1FOmspY2eP2UvzG3ABE4TG
8CqgwO43UqNOyabcCxQgZrMN+hx/bH8iLz01sHsPEvStLJ+hhaEcN6jFFyYKiRwl
AmV+PQitEk/xgt4nms+/kPlk00qXzmF9QIgssZWaLX3Y5X0nr9lMhPDwxD7fs49M
9ZLJb8U4q+bsVDAVCJhpQuGwpv0iQO65Lk4d73H+Vc2cHH/hfpSrVWIw4125ywUk
IVERggJ2HL0jpu7IYvKq47qzoNUd9IWlOy1dTcaVGBO+fth0KYXwXy1wPW7Hd16i
w7wZGfPvb3EpnepsEVGMTwGhFg76vBNWPPfrkKJ5fO4Ryrmuz/XFqAkvsbH8ImxG
M0+X8tTcxpfC7LtiSxg3eK+XzLKf3CK8Ll0votG+lpNGAvTzLdK5hQkQ/jkhPpUF
+rGEQWy4s0BYZQHga+X3S80FcjDrqB5zfzJRbOnYzopUprNf4O34TswQ5bPJoYzH
W084sKM6StBZp3N63KeW4ELhtEy3CKdvqs/AG1l5lul+1igUtXvyafgHu7cmIqu+
gsUw0qZ9pj+SxSUE0tnKeejR43ugKXL7YSQ5xgF6uzQdNE6hvN2cyBqBnFA85YXC
n5dLnguhMXlDsvINGw9jAPicZpjFjMqqZOZ1Jq0EmN9waAEo1/RdPfyNWxWfcU4w
YT7OEMYfUh7Nu5exDek1JH3iGjjSLE79+tWFwQhcbP8IEe2jXWRGVrvTuakXz2w2
4373HqknVH1LYv9y8GyKutdjjHwn3KasXB2xQ9mdZbfDOn9voeSkGFHKGx9HRrqE
LfRUfvXjn10m3uh8HiBWYtS24YIY2JqUJcTNgx1dZ3Wa9zUU4vv7llCSAdRWDn+K
6Js3ZUHcmm7zz/wrPSQF+W000xYwvOJclE0Wnvxuvj6sB/fO68vqkigp5PP3V3LR
+O3+wT/UnsMGFa5PPppcTthNBbqZd7QbdV6X9LgTdQzqgsPfCO2fP/LF+143mCZx
vzXwhZBTRmyqPPSs8RfoaEc8ex4aerH4XrXdPmkNVguChXJM+ZmmZH/jJ6BSW3k/
inINtIISIMEr8BPpMye1O5uHyLd3v6YyEH+8nalh8ysh5vrRQrwQIqSowf2j0Aa0
JxMNFG/1B5W1RBzPwW5olX9XCkQKdvX0+ow+w8izy1nMDgDalKH9EBzdebog3CFu
C5HOc8CpRGUSjih2bpC/fpY2Fs+GjNo6/5dd5ocyxitiRxcgq/zt2FFpnPsQnS9i
l9Lxt8XXJWwMnPeU7VeuYEIl+u9KItjFlozmG5Hk9fNySgkGzAkissNqTN2gc/rR
+LxB/AETgGXnX/VmoRviFxe1flPJpkVSju4hbGa7RP3seuu6PKGoGdHGp2cUhv3d
FHT2iM25kqp0izYNrqVQWH8eA82GLd591QWt9HG3mkV4WlkEgKhJ8QMy25r+5Vhn
mP6X48LvwhllLNuMKkp3/zR9lcvXxBPZk7MElTSeLz3vHCcCNRgr+BqNt1fx7Yyf
zRk3fN4artuu1q+iufKxFSM/hnPd54JK0Qc8JKdGcxPO7IC519r/9ispYvwJ1KhM
mr7q10WpdMlCOont0sLRvdBRm6XgF3E3ip72kqHhhKyc1qGKXK0SkpmUZUBSV6wI
Et/XsvUUvaMutagDeNvrz9Ht+1W41faeS20I1BitT9FuDWwLPNU2sgSOQ3RY4gzq
+lOfThjL5ImJTb1udr4DvUY5H6lApTHiCvhcmy/z8vF0/3ScMiWXGJg9oiV6qRL+
T+IVZIL5oLNDE9+H5DUUf6/LMZcFwATb144qUjYeMwPdWB7TFH8V5lZsh0rabu/U
ZySt+fzy/A5s8MjkHLbCNFD61W2GbKZAshf9haac05zhozzYD2EsnsOO1Hx3qo1y
m/WYRXpGPxYGQ/wg0TNnKTd4W0FAqCr0SBiT/2KUu3hjNYOIvkEhcQHUc0WWlItO
QUwDjgXyH7XdFlt1Uw6OvS6Awnj9ymIVo2dqOsMqpCqwb1lxgvNhOFvlwTEZVxeb
2oOfIrE03XuRwV4jFTyzZq0nkNc+zjlKEDwqzOw0vHaJc06DZ9pMBhivsQnrg3/B
lLC7u9FpLAy/ljCvLmc8UOAQEmO2CS1JOvR1zEFf7QznpyKMJZrulZ/brXGrvRbQ
l0Twv4BUgLc/kGgcMJBnvxcOaOG2pUJDyyYGDKk419enf7bThomonw9vb60wyPcL
ZDXxkJAvNMUxGzfaUnbQYLLwhOpCzUKls4ZidFGbja49epclmSvJbk1j5qpMYPfO
yfoO0crKvVoNVuX7ZfIkGRIV/3b+SboMFjbTUivTS7zd3u6yz3vSOSsfqZV5PXcq
hFM5y2CvLlS4SJQyBgxmFSbDUbmYNpllUcFpTGVgjjgSZM3e8i4zl5BTV/B3XX4k
QTHC84jBz/9EiRoJkQ5zWE51wAMBrDoXyeYYo7YZVwSp9KUmFIeZvuwwFNYeZ6Al
FFezdolGIBlxF8CpmN7L5BYvO5RgsZswDxy6DAXKW2IyXwSp7xroUHHMdh6vDXmy
82tVpcYRgXi7jMLSydnSgGrIZQm2GELMqynOVIeAl0eh2t9UK3c6c5Kk2yI21UZi
WWcc6o9s08s6B3xWxNneTzSq1zHB9NXCir1p66rCYWLoSTBokk5Nqn7BVtI3GfgV
p2BxC4JMIxsHZrTTL5ZRD8GqCfTUu9TJgjaLatks8psUx8swKQ4DL29rcYenXOKX
KooCtshDksRaUfw2G61wvqhuMGY2t/hOVWSN95SVDTRZj2+zTUH+GS/8tAsI/cAH
izTyEIne8He+goq1k9EXyHNMrb5bvo0MheJ9MtUuJAkyFnZoIPeUjx5eLGn2AghV
lOrbcMD+PdC4IqpB2FRxcY+xXMzM1xpme6h7TZTrZoka6LLxv4vp+FiLwiO93trw
PyWQWMUyJC921zFK3JUHX0bBj87HPwT7/9OsHrzdRwPXkzfBOzDqLZy3UhNv8Vhe
diK3ID0d3uWsJzt/FRTYSua24MxHYQ4edSfmzG4YU1kPp9bDAaTdhO82LY1rgfhC
Ji1R7ogGiOGndIMqCRrX+Kq94stRaNWwjOeBbwriX+fe5z24KF2Cb2wiwZAVBQyz
9NvxQ9RKXXGW3BccjxCOcCFLuIQxcrJwadkk8gOIfSVaXFD+D6WRn25llp7Vkb+u
l5o7M2SpBWRsjzjRP55DxJB7qk7f9i8/4fGC8BprJXNZtFJNr6tAJHeTtu3hcgwP
orxwb+YyhjVV2DT63LGgGg3u9jLd4ykBeM+cD1VYLXlEZOIIrPbY4Q6A+7WybtMD
DQe3taphkKE34F7ObWpF02GYNvXFuLSNJNmiMgKrOZdAqlpWF/3WRyGfBiSSKIkW
DtA1t0m7wGLpxqLRWwimTmW7A4Ru1roujrJL24Q4RdzAemFx+pGdZ3J5oF4GmxHj
J1i1wk2F2XY4ZeGJMP9E1o3xWAUSRHU6c85acejFGTShC/0V9wkH9FKJJxKFvuRH
EmaqMnW9KuifacrCx6SFt2w4NYC6PoH0Z/Gb2fgvlkwThOo28lkThFUr0bbhsbAs
1CzxSeNsHOzeoi43hPwzyHjXt/3ouzlxxJPR8HLq99/vTixNUVNOghSfIfS0CJ8u
fsKmS8UY574K3tdskTECrDoog/10jzJAGPCQWcQ96CJ9cLBvEyeRA5JuD6rN2rrM
ZBOXjbFYVMkpSYA7u1F03kpcb9NHMTdIAeRL6giC0asOGH241T1RHnH10zv9R1Vo
QQOmosKP2mT5LdlVh+tWlgdhcUjbwfeaBOiYhxqTbAmkYLxJEKlLFGwLKCCvxWJQ
A4QvpHT7GUvsqOQmWze3UvZVNVvxxDhQwpKaVn9D5uCT/jYzgmzn/uXgPrl5jrAi
EdzZqdXX34o2JmgOVBzUKPidFBeEIhepffVF6Syd/8UUVrUIN3dd6WkKaU7s4lfi
/t1yTOODtR1P+TLMVw52Azpiyw9dePOA02n5Wu8PDYQIUP+i5tK/Fu7ZVSd2Ywjn
ANbBsd00iP1vGKV0xbdzljgOc6CtL96L+MMo/yAbLh7zFat74ywydgSWQ1x+jJPT
u5ps9p0jtE/b+cKNUYgO6KcQDVTkCQVcJqlN/Wfweie7kOPegEkVSanpDmHarLEk
SosRh/5qxbFSVCW+sC4oSMnwvimoAlijNZSiNyZFtUllIsgUCYOWAzOttb/RKpd+
YBZZ04fFyfZ9Ydau5ATBKLJaMXUScJPGn5elDK+HKfeowY9rOzDumhQ2UmmVM/Di
1RpXga7Dxahz8ErEbAEUpjmXAf304D0+PT9RlvH/rUKm7SoqTEbxYGhDrq15OBAp
KBAsML51/Z7NLm14kINTOxljvAsdNYF2hDgRlzMfwkEsAv5OcUfHTkSW/bKL4oLE
w0xSFGU/1PE1Ao/mo+TnYLZQKT0GRv55MaKp+4O0NhKThqAad3hix1CuUdzQ2xFs
tlhAKQ5uXH+i/ZxEXFZMHdW4tAg29IW7/sr9BiivgzW2R1R3n513MXCi+42EgbBE
vByNS+imQ0+10ZL3HsL3llsd89s7kgw408MuY1bp1aKO+Tx8mRhJ+nycPfXD5ef7
yLQpltTTqnCurV9Yo7sjGNjWbwwFhodvJUfnbYqjApX4fXgFl2tzxMNp6CNbxrYM
YUh/TGSstFEM3hhp9kvMDm7ptI/jJZBHf5kSbgLwmgrVs4ntKBcQoKUvBfmLBi77
9zCsLmts5My3+RKhsL7W5kBSFv7bQuCFZJoaoDIvKdN6tHMba5lfdjsSVbdB0qcv
GR4SA8TUVwRbBEljjyvvkCcXtMvzsnJDY6lQEmdNj8ksdO9C7EM4LkBVgU4flT30
6V8Mfo+eiCZB6NHr5Nig4w57XDIK21pPiP0VSGKa4zs6IWrdOwtW5LHXA5sbMBur
tQKeSCL621/2AfPiDKmAxgguvUa/VxzXfggdMzaG8s4efozhKiDbkYFkkOj7emJ+
oby2Rlp1brvK82Vt6w+6h5i/70Ex9P4aNUEuEynXn7SWo5YB1/M0XVu2WJBaSIcm
LCnNtVYuaCLMREK6ZNBtsuRDaaZSJvp7nr27x3HeIwwC3ckfh6nNZ5i/9QbUGKRY
FdI0/JaC6BQ+lwXc9ovomWaGe/JazD+5NIcMGIzS4b2xdljN9G8k6taNANwI19zv
jRD1cnHutakXZLvQ3gxg6pPLyH5lMCE36bOOShpL3uGDzYEKFKcilsVm0FtDQSzr
VaT1T0mEPwexT3ohJEkjZgqJ+N/FSIBJrDfU0oHRWrHQVV4KGyo/iTqU3Oq8RQVd
SDxfMnBZPqa0yhWFTlOq4EzgyVnFsaAT7J5uduz2B3gSNnPjZICZvbew3FWHKxvm
OMR1eHLSIIcuIbaeo4uAGeiKuLYWTzS+ZQ1izWsZ3cMVEaH4+Y7c1JMvF4/foMhk
qGdXcb5MOv3IxEDdiJjRCqar35VL/wbkJCGS4W+tmHhucw05RJpfFAFXD95T/U1c
+N9Zx+rTlMRFBI6sWE5stQMhkpbm0QsxGhCj1Rmog4vpc/7y24t7MKNVVmA1JDN4
NRuFHtBYP2ENzLGFfDPBrtAbrrYg/WmM304gGbBDFKk2muGbQk6PZy9p8uoBQhZ5
ldEpr0PY1Flc+sZawnoWXCkQFI8FsptN61BmZ9lwFh5zBjpAU1gIjQyUFdVmaSwZ
5wy2bBL0u5Y7zTWWHORYagKli/r0g1EFhql6ZLxp0LQAXMl1aqXWjUokN0+PLHj4
8+noKjJ0aUJRk9WEm6NI8om2CWXYrPQajeSbpxvxtPQyzvL3vTlS9ApFlLdi/O/5
EiiQiSrVJBgZsb9isx49ImOFEpaSzfofDApLET2PJMb1VmxBW+b4c5sBz75xiZQK
Ln5i1KCkYL9F127Kag0RrSMfjrtRjoLwH7hnqJSoYFk/1JJip6ZboZIv6LhMZHMB
PYdwVwbRkUAwdSO4tl9IWq6I21gCeLIOqlVQQZcDX9g67kMWJB3T7NDBVTk34kNC
qwVPUARBleSkRHr/JW6B0TNVuYqCpUESXhZHaapju/Ts3Wzcgd192i1m6E8A45nO
mS1H/AsRehtt1L0zffGwI7Y8ceGdW6JAXgzVkbwH2QZ9X2Xi/0Q2JTUc86+JMIoW
vnVKJcsTj8ym+XeMaaj3gRkY0+vvZLpK3nBxRbsSEXymo8npDVFo4VGzZDRMNxHL
LpIjgcl8Wn2s10vcUj1T69XUyEH9CoJUbQTfDB7c5FZnavUtFiOm5BYe9smSlECd
ywvdSSvlID8E19B4AAT/UKb1cwNhZnd87ZMzUDFVQft0CKQSWk4K2CSzHMcpIn+E
XVW4H5aRn7s9Hl8Ys94sAVUganw5tXuoogW8iZ3/DVpBxstpEBVpt+/SKmHjfoiv
bofqY3+Ha6CUBzUEAwRs6YR25NuBVVHv2rPPZP2CGD8PUkcYmS3B8hZdl+VCSd2B
QzZvswWvcASJEnxR7M40B7AVD62YN5G/2cHK4qBV7XedZFoRlAAAulT+DIumY4Jr
e6C2rQlJ5A/ReDnZUv3tDY0+0Rt0SmpsRlvO4CtfPLfKna1RbfvJVpvoHARWAMYR
xwPWMsJA2z4xk0TqtxDOtFp+hpYoVVKxkjwQcM+3RoIyZxK5win3cWSKELjILnmU
sJft/cYYGTqTLXA5E/LQlS5Eb497vOe5rYuRBlY/ZwxIjHSMydNlwaOa0Zea9Wca
djYiHk8VPI3IKb8erS03GE0wm8nYEtHOBQ6i3FytyCdMRtXsPJktTyRMw7LjbJdi
EI3PrIrz3eyxKme+QbUX00dYy1lEEbaOlcVEZd8pBCm+QFfTLsfVufoOuuacF2qW
V+Ml9NqtAuw5irDI8CXIGEGOzrrpRKZl3OzFznJzkS5iZ8Q/eSDUmRL2XEzvZNNQ
IhV6Ov6q07p/b5Kvk8dyfkYOF0tWJULgY9KxYI/0XEgzSpZ7DkZEMsyMh21LzU8Q
rXhloLCmHngwYBBWpkkgeJFrj+w4Fi/kjAULepW5d2lyVfgZl5mU9L/Y/HlI4o/F
HCW+Dw26CxbolCCk4Hr6Vo8GqFkapR+WTkSeuUAH7qqbdAlml6VePIXV/OePLIwC
OWkmzZhOczxpCpfP8S0Q7Ew/y70zPUAasEZfto7ZU1Sh73l7KBM//MLpknlSmRJZ
IB8xbY+6Dy54paUkw4mIsEqMDtxeflP8bo9ekmFhjYSJvX0Npk1vw60u5zHIpaPP
TCyChJW/OP/4o2VQo1y+uV/6ri6DJ54W6j8io0iCORNNSoVEgauhlhbkOxKXUTwT
wn9PJyOofbpAsrYZumREOOu9hnMjnI5Nx7BErVrkZXqeDiBv8AKZHJZPyqKVPRwg
cmWK7n8azvajM8kBljrFjO0XCZwgxxnkwtOZGyUbgpRt17hoIa+a3vPiD/RBk8oy
/fXVbFWrzyU7HUtatNsSgEvp1poJua4qV5EGw4Xk76KfPq5s9NuU6SFMqa70gwyL
Yvu+0eiCc8rW+5kkAJNjf9Wsajmj90FnavIX/MCbb4IbQP6yAjFvexWCRJY2pLUO
7fC8p3Ob2bAsbmZgy4C1dhtK1YBUwRJLDRZBFH53U8nHRZkGTx1LIE9NNvAnvWXG
Wlo1H5zKEHF6oH3s8XKC8w/l0RX3WOdAk2fjNnXycolhCUEXb3bkU0kkRoqcNARQ
iiaheLrFghjlRnQbOxXMLIKROVN55F2AW9vp6K4tS8OnX9ABXkWwxpDP10C5Ku2e
ltpZgsRvB5T+1Ogn3SRGkLC01PZPWIn7+4soC8/uyFQW8s7i3dnIoTIvIEzu9aRV
QbU6YWHG1jLPshvSrWdnEiEwMlP/tdA+nZmxX3zKk1qMoavy0Ei5jR1LTEDlcuiL
cj8odtadg6/F4E7u+d4mz9nfL79ufESPpm31ne9WkjdfyIXinPYYqaymk3U66CI9
AlLZBN3Lwx7Dn8ZAJ1YF7wME7XCLXq4yIu6qEEKhx8uEdqvBByuh3jh+wJBidssY
FprSwuTqHXnfZeBGlBj/KkqrtaQA8ddyz/ZJoaR9K7r5NH3yinoN7b4sz7bqOaW3
Df0bL2PrjXmdO8DizohcyFY7G3qlzNJnf1nVaDgjc17181UeNiGUNenBfVgITCxt
CVL9i0R55t97n1G3eWdyGXjm6Ssn2zaeB0t3ACjewtjupmc77cik++fKKNIjTW2j
ePcShhGpN8+yJgcrFcjofVq/Fdz2Pcwv+hrQrhRBxHf8kZ2lR7cGJiEDrZE8CRIC
qiBmYGBKsVFa0yf/6T2PXQ2mwKJbbiB6G11XejSngf3twy3saMRHpe1IiIpnrPHQ
fC7crr+z4YYSM5t/BBFhr8DfSZvP2jQFADQoufOBY/PIly4iX7RyhkN0VgEG2/+D
bI/teNQJXGZNbiKuzPKi9IjJ0du6Sit1Y5N5w3VYndsQC+Mfczv14ti6Riw4RVhd
/GE9UvHDRI1clSdrQhIHzxfdmYcpFzeRsJlH1AUbF3LuZaS///EVIpGr5Vtb7nry
i699sHhu4eN+D7tRrLPLesR0B6AJaTIWh1lJqYdkUYAEEUvP3/Ew7yh2Dlw38cnN
OOTDI5XDgnuSW9oQGVUoOrS/Gtj0weKAs485bl+dCfmVw90G8SsUC2vDpyQJKLvI
sjsLBc3lW4mfV8Q/K1ZugUKoK4uJpR79UamzelwjWBr4xkE8T5LcO9FOpBVm/aNV
nPKNt3i9nMDVfxHiGbAWR+XufvsubiDFJMcPmG0ncQPw/0ipBlaUVFHCshtqD2xZ
Yjzbs/SIh/N0ssYawL9wPZmk/PZtr+OuhtKpZDF1F3pUMAvg0Sj/NHYRk45rLUpt
dWxdgKKEc4EGHrX9OA39w+qKef81kYTA5Lsn0MNch5FDO+Y5WPkf31LUqBN/Bm96
ZqvlUlCPHH4kX6s6HEMvdqm7ZOLL9a78SiwY1FRNTOKnHfCj0iB7mhFvX0CaWWdp
nD3SYDADafhn25jfBltBvEzAdEiilbBehIao41cRmwxD/WXm7E6p6bZtzTdZcLUW
APjEHWpd2Ik7f2AdAgJblARVWrkdwXblXeQxBCN+WupXXpWn04/uHn4Zl0iAqMBH
X1JEE8xV5NjCZTaAzwwvSvxmm7uyhit52JWGIjh6a+HgXwczQiMQPuPHioA+3WJ6
9F7Xz3Fu0nMQ+mLvPkclbinB5GUnbuyAnSS78AgbvFYONF12zXEEWZF6DzjLYHJq
mWuHl2Z2bTSeUpsEBr2BU2FG/bpOaRDve55010Gx7amtsdo01LfoHU9kMg9j8AUc
Hct0OgWj9GWBE+XvoLDzoSZh6AIpy33VV+0fRFDmY62hgWe3xvgYlZCLqfYnNG63
3sO5+HkoYj4Thq/tWLKoCVPKODjG/oRyNFvF4Ey4TvbN/2sV07MNolc1isW9YHsg
nZUCnwxCzA8eWgq0i7C4B+EXSuTGvAzHRKCjfrKNsZaSLcLuPIHANKkfFjHv9eHN
8DtPaD6E4kelLQ7vuCrAsXWD0BGcYQZOhIKN/bCnoiMxaGyy74lJo+uQEQuaJsQ3
roNHjZL4+7KSNMGAtnBUIX3OWbab9BYGURIs9DQ6piM4MsBqD5zigSzH9FP2XpCV
z7EhNqdkUkhiiGF6PXfaqWNbiLJ6MWeRont6e/CFLajbjDYAHgoXDguBjt/kS9ya
du/2h6RfSKenP+xUjLpPJ64utTGwMHYKW4BCwS+gGkFRO540rHteOCVUXj1WvJzT
CUaS1/R2Qy1vbbaTCkVWJT0u4cJDQwPSz7DhsJ6J0FFOz636i86toFYJAW+mS7Y0
Jk50e6RzP95Bf0/rayE0yrVHYZyMQ+WMR6averbxmgi3ZOzGERqT2n5O9c9ceeN6
Ekzw4J26Ord6bojpwJH/q+PHlf0QUkSltUhls0nm43Hon2TfH5Q2j9VQNOIxNaeS
J1E8iSfVJo23QZqya475Cz0uBVyIBVbQt7RTkFpdmilB9Y5CI58VefxF1Vm61N1F
EjGAT0UpAVrv/dYixhRiWPDNGS/9kkl3F5K4jUHIkfTDVt3LKm0O99F+6RWIKDjv
qIC3sXfpREszXZzX9cY7H+scWKKcoqSX+5ydkP5Yi++oj3oMENbiTS11jGpxKd4t
Jlx3QHF5NHvirhR+Qb4PlqdnILrlcMvhWlbHpNr8BOtp01lNxwrZW8d71PEz5HiV
umr8GMG5M/O2jOZ1iBRdeJ9HqMFCSIJQ8bPhAvk+rYqY8CdlOUIMKBg4sFmS8sG7
+PZfh2kqrLgM9BIZjYPPaafImad2uxh3d1b9ars/lcVmthaYq/Wj25Jblxc9JVZP
UA/gWHaD7I53y7XEAhytp+XRZ7M/i8RyCDWdkN5YB9V354r3oaMZ85GVsByLuCov
cRlkO12ioMe8plHoecmfRq6s7xaBaZBATzdiu6a4EAONRQoN1lqk4Dx/T+YBheYP
/26DnKTb0t8WGFFOCLvrVwkWP0gDooSVMPX7eRjgBFclkmz8ncx2KY7jEQSWp+LJ
B3Q99YyNYuQJB7UV317nL7MH8weE3hBkG1yZUzGPA2JkpOu7hk7hZIuma6dunKGZ
7e+Jii5BQ0GgjAbtbsV4TrD10dR6YsAI74qCtTYDxoM9C1lG6/tmKTZl0kAtoegC
WENAeymrURzwC6VwSWjDbauyETKrdqNFrBOGheiU491wJW14kc9ybcHtjsEk+J5L
SVwOuFKg8LHOs7HtIKVv70BQW0YyOxx4IUpL1pLK/MvSXxqXNtlvVqaWeTgbsE1W
IRi7Fu+M23BEC2CaPqPIJlqUOyX03dtRpGsPTFajg3MzVP5MKdkEND3C6ygsA7gq
Udn8oXWxWcjwbZYrEU2X/gGX/rGXFcbEs2ognfD5YDjVyjGlBNFwK81L4CnYoLzY
FXXcViWJxU+2QnUnSs1KIAjSPrV3OrByNu2xwqK7wYj8dsnksqsjhAS+6PDzXuaT
3sA7SUAHqdRp6F0pc6SPKXg36o1IGi2zO2MgYfY0ZPDuXkv668DDYvhonOaNfeW1
hSQavEqS0qE25N8ONB9Peze34V9Tp1kHMvwsM9o5uP8de9jMYImykDJW6mGyZRMK
WFSF7E8VLLbMYCyzJb/4n0efkeFoXJ78vl9fizy6+amJ/1YxgIH0MH8Pfrlb1PkF
2avr/hb+t6U7P4JsJaZirRQGRdRJaVyQ8wudxyp/inLk4uifLOkQ05MOHNPfPlCB
IMzkPzHUfex11bUsb9EmU6LwRYm0jvW5JrQ8OllegiZOhHaK9kCUX+cgjpaU4k6X
mAUfVUAFfU7LKTks3YIKnpvSxa8syFYAK15oacdE4j8QxLki415tQ/bYj2XLoBfl
5FYlobgi/7apC8bl+pMNnvRplYjsf1VlWYduTIQN/KD+X9t0LcNzImfcFAuSmtM5
8YADRICH3XprvSyIR+kbrk9PHPmGN4s10hPw9/DIrHG/HeT2TWaIL/vwIrGv8G2L
3lpBW/ehd9FF1B0y7l48Mky24hOUWahd7QFV3ms0y6AX2yHhpvsqQ1h5meNTXqux
5XRn1Kbu6O0tnMZYVu2W4RJpBniiQfYcjTnNaFLaZFP+IJkpzAQqX+kyijLNp0IP
BtEBIC9cmWx8RKP5fYQkwghWXEZlczEezLplc7VUrKf67Ot4GR/CJ7Yhx8tr0nhm
oY7iOei4V9iLzH98ztH7KMas6A1KZUyY426URD1sunQ3Wghahazm1fNeKagiLNc/
O83USGE/VmizCjeCyRL+/adOxVtj32NUrMTQ9gEYNGmf4OpJ9iuLFhCkGAdfkBWA
Dg3K8AQ+/oj09+V/WTX+BeBVylyi7H1V8dJJBsY22l9n0HI3CcYBca+BCNsd+1oO
5GAWSwwruJfIpdLbCtM/WGJo6tZdws9uRRvcoes1dR/FtS5bdeMXvfeXlFviajl/
OL8ARid5+mliTkp3waxjcwgzd0Q67w/hbURtiVD4TmdzYDefaMiTnBfjymoJWq4D
zo3IyZUi8zKNOUGhJJlJRc3a8qUXVRsDmiBZfUTv+iiqUYgLsXq8UJOQybXSg3qW
i7K41OhyOcQGKOgB0MICZBwYZxT/xSjDtA5fosi4s0w8NXC0CwOiGvQIOpwtqgNC
trB35JquRswE/94wITjK03meNvbFDKHNVH2hqEz6Zn+bP9gsYr7rrd9br7u6fHJE
9f7K59Bf0cXSZfwUdUfWAovoEVcfXDgMl5dpbsbM4+0TICyPwCuNOBMqEd92G3xu
yVrQHTkCNSaDGKUcPmqbvjrgAqR5NrixBslrp+s8Bs8gSK7nOrr5DdqIjd7SQPUT
+/QlPhj5D5PxhqGnDtERtlf9y2e7iGbrTlMj+cTz1uutDizFK/yTEOii9At7Kz2B
elJJaw1Jwfjr/xRe+PX3JQRLD2yPPUhlQbtLYx6PA6rV0oPde5i/p8IxiEX6a44o
YLpt7VLX+xkOMHMAsObJnV6tUuNChnYwNOzKmVTvjtHLuWNH9qV2UADQclThykcg
ngCYLaKWw6LrXR8OB+QKTkP7iwdLkFYFp9SK75bLQ2o9tYQDbzlJVerZoPj+MYdM
SxSFdwR9PlmyaipWsn+rZd/DUgPN/yQdyTOUyM83W8l9gM4ox+iXTVqaTH9BDQOM
X7cdJvePJOJBCBT5A8yNgQGk9mbpefR/DaJJF0SFubR01dZtM7tacrIrhooxqWHu
O48l9n7u0deHiB1Q+l1cjQXLIcLmS4q5ZXEhb/TbD3BPZlAGASTfWnmWCwTzTjfp
DTBYCKUEJtN1eo2BPSs5ZbWIlAxXJW5u65iG9Gf5XDWAukreFLXxAEVC4deObzzL
0C88G4REZtFrmXgqVqqERqDe047PAn3N9+kVQYEYazlC3lFPEqCVEa2p060loich
TXtdxErnrK5oiEmahSv2v9vnguKrRBpRfdbzSL8pKWpMZOqSdSp8N3h8vKhbXJn7
5w1A0SVZaSjfgdukwHl6OvM3hkjg8lp51KhWE/f9nOCq1EUXTmDzIaxs2A6m1BC1
3jJKbzbgpVFqwg9yhsGklZ1lF8SUE3YkbPksCZW8QbxQqGRM77+vbMaxf7xKe8Wt
/usELNwMcH/Zy4scdpq9iZ0eIorn78qmfzNgTeWAB+ddmX827IFEewlfpTfr+axR
IP8Plht0ljdbd90dduz+1cqG1PdZZ5P2zKph+QWhyhlnNLWFoItAygF95lSezku6
XxuN+rObCO7NQtlvd6LVNiF4zTlztQM/OV5U8S7UAHS8U2Yr6Ply8x9cx03SFZTY
Tf/PEkkst6OoXapWIiJ/AxFaZOPBKw53nrspwgBiNs+wL0nl/MpUn/EU1jI0fuPh
SqjnZ0S47tk7RkMKZFtI/SdmTExpXqgUjtrxrYSQQpQ8xl4F0akFfwhC1AZCAFIa
3cN3mocr+NraVG+BWHcXnHtBMJoE4iCdh/BT/uYusiOkyUmCRF83p+aVBC9JJOWS
s5V02Ddb27iwPhx/446wqakZpuowjHhGmzwNuGsUC1tzp2QT5r7kFo7hwTiFkJl+
LIyOollQzfN72xrsBPEatIdXmvOvi/dcR++DW3Nnl45JjY91NiRIrUdB+ewFQjwm
lwif5Pzwqwq1ROBHZwVZuiVABYoGCBk51Y3pQ/p/UMDTW7eKVoeH/3UFBzgiDt2H
0vl/eoZLhY4uCdmNmd+DFgdMFxD93yjVBpA8wNXgiKI2d9BMn3JN7ZO1z+iTqc2/
q2l2BAWy0z7n/3pjRYuAYWgz6t4NA+M4fD4Vn4YntARoc0zSX+PrqyJZar5MS9m5
UPC4EmjVmyPDH//J7cVsxz/o8vrRBy4zwGSvS5gxZVf97s1zV/6hsS4kb0XV2yC2
+1nONT3uM+xgODmJovTiaqGTx61Mmq5j3V4yd8EPrYlzojegfw0UrYs0fHyKe6Qx
rM8DcTPcxM9KpiRXedWRVqWl0A/QfoyNwsTNb23oN1cjC6M5JUx7slvKi62cQiP9
kO8OzHEz0N9aQyNaAUfjL8K65ynbPkPamQjqAbknXiJxvUasVZZ1+NqCeW4Hj0/p
2Uj5gFGENQj4FUAOtbyg0EC7QjghAwLB1NJuPBfSX508qPGIIl+4nfOugGtRn3ZA
04QfAVazhPfhLjZPrNS36kKhnWo6ZgBPNSdFf3RC53dgtvUJ7DbcZ+PjEumTKbB/
3cX6j0BDaZGbnUt0QXu2S5B56/21P7ffXXTSFNLDC6cwNRAjFQ13BWxSGdislg69
E6s6PubXcG2+P+HnLjsEm5foRRRWRGPYIpcUYhr8ogk13Wa7DtVzme059sZPyt45
ZYg9DKS4qMTWIkG9amlEqp4ArmjrmgpqOi2/Vv75bCdMUVxzeLSntAMYVkpSW7Sx
WOPkQwD/J80tKb7r9ynTbWR2m6NoCiK8tLpgVDGaKdhjtpJRyBSrwXJIVlX/8Zj0
gSgv0ZiolwvI9z5aOnykrQYZocnMScjtBg7GVAjhH0MMaJKLkrmSZQUbcF//uade
QE55ng3++z9RuC92TxsW80/oXHuahTtrsE9Pfn/dUaR0+sVS7TFiJ6svFhq79agH
+NrOYV+/DC3XS57MNBlb182pJKn/6vKCBWloii6A1dO29oHIX48WRFmLCMETdM+k
gT2nZRMXXJ4FFawGzia0n3mTrq5vb/3GzwHU7HqP2k3vkpYV71TxaEIIOc92VdDD
n7Rd/K0u3Udue6ZllgYvEYU/EmNs7H5D6+ouDkWYyPqjbNwXTycblBrx0ZTEQwTN
xg0BSDCuPRIXGMLvaYboshhuGzqYVkd0PBDUQ2fsDPHY8J2DqRP+IXGhmwzF5+tF
1zr0Hv64JmMuREuJTvXixCO/B6F76HiPmIm+XnwcWFM8PXkZ5Mhx0MoTHN/efTq+
fVKyyTZtdSxU1KnoEp0+1eKYaPYm4ZjLc/Slk0fjFRt7DQFd8ogkETWjjOQL7kyV
az8g75GLHC1IkgMyiCZBsNP37bkdms9QN0smp5qiXbaBj4zNe/Rzc9S2kEilXbdZ
wZYgTD6fPIREx5pjoNkjO3XD8iG7YoSNfrvDmpbzRWYEIG6mA7S4edLZk4yVrAwn
L+gQG8tuIWH5eaXf4VZK3q0YmIsxM1q9JQv8rEfiFbpd7UaeRUjowBYUNWda5zfh
6cnA0QSgXqF8YGRF8qkYEyspWfwhmeY5usn3S31RPPsA/t9yftwGH1JEuztk+dZE
JI8zyQ2fREk9t46dIDNJNWrQsBR8TPjxS4ztzgumI5czS1hq77O8rP2vB4UKeOgk
9LLdQl0xxkOyNh2pK0GqMJiez9v7nUbI+QI8EZ3LV+B48673nB+VKq+lB9M9bW3O
F5O4Q+FTMUGbG0Ux1gjc4ZEIDrxZpQ9ke8rSApuA/gXhdEoe7Vqoi9lL1YAYKfL1
d88QAr4mrDLOHj/AMn85xDpeclwxHlvV4UYnLTub09R1OHmLdduCcT6bmCQfXR8k
4ocbO7pq38sDS0XGH0RiiBfV4Sj6HDEMJ9+MfxkEveRklbG5YvqB2yJcjuDTYcSU
PUd3TXEhhihuTBliU/hE/+WiNtyTcY0uOsiZGqi8hnVE6FBXIOXaIswFv/fX4Jms
f8PO2Y/NN1Ps0CCr48ydaIOTUNTBMSa/2XK5n8YE2s1FtgEhjvQnIb5Pmcg/n1F5
xDu86cLWsIWainiePwUuOwpu9QLBf56Nie3W4eRwt7xVcq3F4IKnFIC/3WtLGbPq
z5OX28exW66rOEWQ03hDyHYeunNN5vEtl4prCvAADJc7oseEZXjQdXOtNm3YQwln
52HelmV7F80iYMN67UQUHr4hVSnP8XamXrYRqdFEqxZVQepolFDHeZW5gSCMvl3U
wTiGGfo1WBJk2GoUKtk5Ltsdqznw2vw7CE0kMxedzD3pSMm9qzVIPr2Wk9UqF59m
RNKir5UHeGo2uXhhMjJVrsrSlAcsqJmgGFW9AN+DxsVnjCBKjM4SgMSWCZ4Qs+P6
O5Pn72yU5UvfQ8g3lCkv/aReq+xpVcd4QtVqiSm6uSORE+8Mi0rkLPKl8dRXSWlS
rcXztuQJk9wd/2DHhTf4yyM41HsMfRr44YnpcPlhMtCnZDwJWFZo75wX+gchdYIY
SCMpvj8orjaXv3lQDa+s9qTSute2U82/UDbCo4/4Wy2hfg/0f4MEjT1u+ZT6cNWN
U5E4L5JNjffEN7WMXGd0Pw2mcnZkSdOActokMtLG0zAyKE+1HkfxRKiEwML0GGB7
+BeYavfKJDYt/GOqqB+U/GhMVvMVde/nNbsJE9Q+CCuDAaPuLgwCtvUiWn07jE21
pzBJvrBIMI760/Es0wXX6Koo3sKrPl0OXQ7CklQFXUpwB1BSgonW9ebBCu9HZrJK
iD9bIWCjghoOG+BmjieXat2F/qvjOS+6WMmaBxq1O7k+BUONBI0BhWh/TxdBdSl8
v6ouaLLgIagufEJHLJWtomzBvEM2kqb0XvxQ0RgYcpeJR3J5+bCbv6sidPlpxqY+
woEwSp9HXB9i4N7zf2yJoe0JTjX/phshXqHhlFzxBdBAqu/UYX3y39u24BG+4I7f
xkxqylO1+tc6602Tzi0rbaiyH4W6xYC9F5YMaq1lbcKGbleOPKhJ6CE6rNO4xbHv
ImDg2WjBhGiEoILt6mx7tJh/ypA8zprg0Ms56LeSCHo92YK4c0orIXIXYhARz2mX
esRutym+sETStuoPva0d7KKxgTH0Ms/SnDk8OeJqYTRjmJxNHCCeebuzfFhpSr6N
i1UPPGlkwLu0JdPhr1b9L3Y1DQ/7H2dZF4F3SHRSZeC68CmtOVt1vlHe7IaQcgbm
8CmFpGPkGH5fYXf61eWLFxAgIdoq/ym8IhwBU5dRGOmnwwfzjJ6r/+dMYx1+S98F
MQH/0yehpTMK5uqbtBM0gynTEphMJy+lLfIXmm/TBdmw9k0sJZMJbe7ezne5ksCe
KV8psW0Kl9o8eV3DFWjMFc3zK46bodKbZJ2S4aDRbwQGMO24REV9wbf62D2kpwEj
tbDqdnTWiLoWitJz15FVrbuqkWJnCxliDQUcxEvjZHzTO/31EOn6v8IdpVQfcF7C
KW/9GaPSqNmjSQyMbIa+Myqiflfn9Gk/YeaTcYxZ1s9e3zdoH6wt/Sjfaw5hZL1D
lLIqezeL0zaV+Q2yBdPZdGYkhCOD/pNpwUEH36hdohALTwbasJBydrQZVCp1zmpV
dwies14c2Ph2Bd5dI7hMv78rOWCW6zH3zCrDCKZfOhisX/YLatGpSH0KGgAZm+uw
Od5UrskSSdz53W6SpUew0eWLS5g1vtMcAikTBvSFg3T6WW4CL4LWRapSJs+goAXi
b5R1ZmxFQ6GTZhGJaC6VsZ8wFcZKlJ4rB84zWCEzAR+jQi9TYLn1ID7Vy9SJeAT0
8sShECdcOqeclWMdu8b0DSmSRZXo4r3ybd3QyelNvXLPmz6XyKhCTkDA1ysU+Gcx
Nwsf5+f5L+EKX+paVZF88hkmfZsDxIf5PVHgfG6gkqWyFUwFYr9V+XcaYku/f4D5
uhP5FsJaybYuQzS10eW86TwmbopfZTGtPuBPUl3s5gJavrMOmbfOVCz9QZtIZfmy
/xUHQAZqynJHbAxyK3gk9TUvmENJn4BTNgZyruNWY66/H1gkpfyRzx33dkNhpEB3
8CUblxGmDVChLIT6vB7DNvriOx3RcLsuvVJIb2utqp8Vxh+xPyS7V3RauAhVV3YG
uAX6PFFVc09dFByab7MTGB48+LpsPE5SticJQLHhqzV/+XzzPh7WvZ2bKQNdzy/u
6q6195y1rcUCg24VuJHBCOffoudgO0fqZ+f5sqb3ZJtBF4cW4RK+YvgQK9FuHxFt
S5vnuj6Rs+DNXwp/IvIAsQgQFhpmOFZ4TKtL842Yrm/22spfaMvVcc3jKMTTBJ0O
zfWbuxyktn8114uw4dPsdHgSsR56lsoRZ0ZXJHOjFC5o7EOyeHV/Ns88Jz/+35Ui
vzfsvz1w0M5BytgQTn0Cwa8sQ1xOdM5GLftUpxKRTCbJWdQovhdIDOWagrfh+Xvc
T0xOEzs48lku5vRP9Pzk+WPDgBTe5sxw0m4K826Izu2VnKPIZJkUFoE4s/eO60+1
P0qOjoDybgh3tjB6scXnvO4u2+0D6eEVeHsWD2VdEJ57gp+llhpoISaFKWZInJW2
BeavAbZ3z0TZ+PHVCwpaNkNymN7uREiZ461Yw4d7erUTkIcBu2pOCEljXh0xUU8I
I6UG6QAaclzUxjp4Nh7fgcEQb6Sg3GPfxvWY40p2JTuqszfftkAON46NZh04muhv
Ebi/F297LHY1TxN310tSpfFp9xUazpDCZ/MI4NkRlaj7qe4Ms16CtuLyOKm4wvv6
HmXj/eQDK3+h16dmgwqN5Zoomwtii7H/kkNtYQwba+CG8Kg1FEUyRUqJkR4NT14g
BkXjI9Bk6GWyrTTOKnd+m6crJFKutkNwl4ajtaTq+e2/j1VyQYtvFO2FZNP4DOfi
y7spPfshbU+hOZxnopjf06/1iVkEGXb/kxU738dWwEbEJrqPPyYe2Cb+5b2BL0vs
FoQMaGDgedV5tDotBqs6vaVjLDgu0gW+Teec1J66Km6yRdj2Hq5wgr5A9qVe105s
D2K4b9swzSk1qunJQ/D2nXsWZIlmZxC86tRSaJd0FrKhEss/PeXa5NwB0/SrEFG/
1lth0kJJx9Lo2BHFFcwxtzNfF9kHvDR41ZYp/QfVC5fnucxQUFWmGS/0ZexCEtGB
2wQd35dkf7H8IVa8PoSAdDZyQIs6IUoLgrZUlz8pW2DR1lHPvaO0t+/KM7xwfNuC
cKy6lHE5OmKeDqTvxjwwx5xKvY8farD7r0+K7T2Mqf1VnTUmTHGQaEGAyUnmD/zx
uCom6LvbmRJC10mA27ysih5AzAnr2k6hruond3WeGCUYJ7SYOj0qS58QQobblS03
xkrXJeuf2wKcI1Wf8X5mJvld2hhKDBanwY7gbRU7PXp1DkSXkDinwZS5qf73pHa4
2dPE9r+Vf1XZyfO9DL+w1dun/u6SrCiuXj+ZJz8aab22vFcKeJ2THB/ScZ2XHz+e
dVLOLNLablMW/KQyxpHqhhR+UPBSCtjL4fI9/pfeQvEFtuFL8KjnMyVoVsEq+IX9
atjmAjliyVNGXh1awAQUgb/JyRpt4CesZdRBTFZgrFpKVRhkTqqM6RPJ7W2rnWYi
utHnRA3eMQXAtYjo2sHzD77mU7EggxWPyZ/B9v1OvUrnFGpGCFTgJtB5vFhXNRVh
98WBCqTNiphdVNTVhGch4v43D845j72HKF9LHg+m9fDLNGJ/u7jOOrmjzAxRK+oR
mXe3N94HTZkv5VZZHRnob6WifW4qP72OEQkLyAU8x1Cgte+2ZmblvdcdqisTO5rf
cBHwBv20ulKOpLZGsAfYbCPwNeT0Eq0U7uKD8iKZj0fGD2/6wxhhTTClZvfl0Lzd
7AVkBRCexA1Um3lKk2ZUxetw6gJuqtWyaU2v8yGg4m7gylugxSBM9HgjfBwp/s/E
4ACQibvVnFsUaAYzVBD3DS9SRvjA/kQilAJ2vsxn4Ltbvgvm1PeE8wyZ7v4RaHdG
5GmcUoQTEksipubttFy2DvZ2qk7HOg6famOEfktrZmFXRoYpwrdHAQul2yNxY+dt
5xZH7T1axFQmv0lGDA6VjFfRIOot6JWtQNlgAYxDumUNlIt/DeMKcxj9xY/Yzi+P
JMcmTK5B8JD24C4ZdJVqYNruqi6zMEFLElMxvFYQiQsYLOsF/PEEZlXXXgjnf1gK
CZ3IKOOLO3YiZz4c2x6QP8GM74TITrWVe05/SGJ7MSFSzhBNfRSFEXYAZiGWbCc9
/QDRnojwi2SsfHTzEFe0c3F8wDL4NlPP9uPyKwCcak1xJ2TUP2+Oexhp+B5EooVg
A2GaswdKQVjQYDPCGoIxLxKKBOzRoFJVGH0j4HFaI2Y21jW3jCyFVCNGsMAf6vX1
gNI49xxQd+NR6DGzLmIWE8vEs+a5y8T6EmJbzKHnf7KvFhDou4vdzKCih+chshlJ
BERW2av2whFe48H06FodxicFIs6LwzWkcJmuvoeDkipJm7Iw3TzbBYomff/9HOCf
GnxaZH7gGl4GlLBPasSB/0VhahaFQIorrLItlLol9Jf5knQFQya5yMwDslBwIF6/
AEauA95YqFWaeoIDG8dzHMa+EAGgVAf6+amGNAfqYvS50wrLA3BXUjRxglXoEqoS
S4MA6LRjNxsdu42z91DehM2h82HiJg99Qrm1WUx16Lh3nvPy6DOS7QES6WG4n30X
G93V81QHnY6JH13FFy0IgUgMvT6JYOOXgyEui0L6Do4qYhXrMNG+0WVn0QPCJRBp
txamiDE9u+Qktr42gnNi59CA+jbgus2fm8V1bHM4eHSRtQBbuIzmr4Yt8RbA3LdV
ZaSSNdvqVkjV4jEmfcOVYq9B67qEnsQx9iDlH6xnZpTakx3S1jX5EHiK+Sp25CEB
YS/FyXbw+xpKRfVoexsnnEgOjl4xiIBp7zq7+9Iph8SqpS3JkKDtBA9OaK98og+W
74U90zn2lkOMdNneoih7MHoKuB4MAyZscCK3SQaytQUeqc45bufo31wfyOE7oV5/
GzTMN0dVxmvFr5cUS4E6mZsIGQkE+GaoXj0H9/hDqbhR0RGAwFRIS499Ux6ct41b
+/vmlWx0XtSVN5WmzjqqqmXsiadNyvhyrmXkgEOiB7T5OqX2Hulpwj2p38KHG/No
swQX0xlPx2Ketf82u7jnu/lhA5zczDYCWshAgxynS+Q5HYSpYe/g+/rGtkjDymEg
zCZUbEdKkbmI/NuNhZ3G9MxPLhf8rZj6l1JklYAB0uH7oft40g4M6/M7lH2AUTeI
SJ9xYltnHDs0iO3zo8iMe6Mly4olxVQS58Nogoea1CMFyURagqIImyBq75crLDhI
NE7MJb+XzOK4c3Hxepqkadiq3d8kyOuy1cOg/81IGVbDRqfn3JG5+AgILaMthW/c
GAKF0OQbEgLzXQ31eoOXGW+lbX9LW9+t0eZNZN5xgYuWWk3AwKvouMgXtjOcyHN5
EFwsrbwL98O44QMmFxuXpxsJX1oeSlTwv5Bz4WOeRouaZMSOoYUvrMtnC/v7ydeH
4ZFlTmdmab46cc6qAVk5nbPqr2IDnJuaPeQMxsUZykoU87stN1sGCjZB1kTX63B6
WsJBk9w/3Sgfh1ocQ/jhjCnAVFaOG9G/SacmUoZtFVlpGMTwkPufj+R/4UtCWJg7
Abuq9uO2qxcYeAglE4ZjeDIxGctu7mymT9mC0Z4I+wFJb1fmESuXDdceHXnbUELd
q5nCLBuWUuS5tnnNcmDJOy99CgShz9o/wQuzCVu/8NXlBPP93+/r9JNfIBV1+XQ7
iKdRDYR0Hm17s9k8GtqbxVMYKCYV0G4BA8CGuw6emaj6zDnIlWTKsJ4xT4ZBauM0
ZkzmD8DyAYwSjgXo+nNkGXwUYNvl6r2V6qddlYQkh4Lr+WvRAStbFjD1S7q0Mso/
g7nbpWX9Nrd4re0O/7RBd6AcYlzTgGuRnZeUKjHxBp24xdlUlWVErfRRS0tzXSQj
oCUJlImGuoKuq4oSNuc5cvUefVNKdBv8sZxd3xJGtMxqxyVodebWCeN6S784LVha
wKyY6hnRxMjoQev+ytQnhPeI5+yH3SPjTFVwbIJfj20Xj5+KY/zvM/5s8s9CmbZh
fhX9ZD1Kms2UFybVdWD8lMJvR7Xcev9i1GTsUB4Hye9x3onLiNjHHbnHwgD/vov1
kiOpZIlhNwXGufZ2RSZ+i5uF0gayYPd8BmnKmNQGp+COdH08jxUfe1KENveouDif
L36MttrZYvU3mJgjyGVE9qXWhg1tx2oKFfOt00uVIEnxhU/zDCdla2NtN3RQU91b
9EQkYGZz/hu8EzBHaiGR971LfLk/YIJqZvrQpW9bJa0Fuk85JYqsYuDqb4AaQYEB
kXozqNoVKZtarDg8psjfTvCEn4XwcLV6XLuXoaUrskYo/JvBGUF1hPx8HALmZ2Je
PZwV6anEo+qVKh9jcrcHohjIqnLkMCYpcBH4QyQa/7OIUtZcLAP98Ow8l/ml2d4o
ku35mloTjOuc109z6p7S3VyNMm9uPMLFJr0NECWciNZfXdseZfrkvSCoCpt0WoxQ
fy2t7Kz8P93PpX5szA1L/Ro53bnmo+7QvSpioWMBpltcSwtgwOT3glLtZQv2hOjP
t2GjADttqdlhWMnD3Lu/g/+lAN+zlbRVUpKF1CrGtzYlZrPpvDHFQ/AI19ALeFy1
mj82m8/EBdvRCpCN+FU4Vt0bMM/IN+1JF4dG876J2CDtksTg9AN+gr0xdE8tSHB/
HgZhMRGnPvf5EamIH1SjFYuqFNT4llvGKmCf6IwjCJ5mLXvXdZsM2QUTuQfW0DZ9
KrOL/mFkv8gO1+vxSEo9wE7mMbv7DAlU1JuKvWkODTZd7s6xHVqyHDOtwUI/LTi7
bbu4t5VJUqSHBkPXL9nzdI6vd2ttrV4H+UAygcnNy3sneSo8G//pcMnxqKhBm/U4
WEJ2qsIXYWcyRudHmjI582ZQhgpicSgEaakR3dU9zbdNMGeE9tLmefUCRM44Htmb
9aC3/Tg08RPkMOkXnFXLrEtUfbynbBO88TkqFjV7YQ49+MuVI4jKUYmb5ckn8gtX
ogegzdjrNXH7/NQLHPa46sBo3FIKp783XKOmXtundyf/UgyPphpffLS1HS3WnvEr
Iwl82F+HJ0cTTMfypNcofjThovB++AJKR6QtlxGoopS29VU5ihoqF08rfxXMIqy3
k4lJ4Ap2+n5Skd+zLPmP4exRLhGehNKxk4krkHG110t0u8C2ceRwXZ01XcNBVbDb
VI69X9oosjFYtu6cGl14aTZeb7Q4gpCSYwIubY+yDIrb7I7wRxBbiKdG2vVSTn8J
K/608BdXxuoCi9QsECHGBXfrVgM7hAETWefKp7xeij/qLIspiwLufWSotNAkr4SQ
9gWaghlDQF4bGxCP9cp+pDwgYVmKloX1z9vJOISIhjYfdXZAvZQtfWYLZ7yziz0L
QRnyG8m9r1DB/98cCkvIlIP/qhLl9ONXb5vz8pIIQkjz3WvP4J7V/KNaA+O++oZK
ulu9TslL2pvvXLZK+BhVJEvQHLlFAYAwuoimN5cPW4OFfnLquUm+kkXPNaP9CkFv
sJS2Ll3+UnVnHIB7my3H6ZvLHZI9MhxIa0sK0iq23mQU9SPE2s6Z2ILM+l7V5puf
hKBb3xqSpHlaUv9eV/1+M5kBgAYUFgomx5VW4XesorXbDdgvgBVfUi7w5If4fk0j
p+2DRPledGViihsZEqj0bVJ0R9iNlk1ERl2vI1eH4NNgGtAVzXMh6ewpt2BhZNeU
cF860BWlqVd7wN7oELYoiOBVQuTueksDEdZB2Lkn6SFYpdWZ1bmv0yGru+ppnWT4
h9h0+bcvyE/1IKrSXXc+E0i7A0HTWtZLyrflQR9I8AlQw60ZrAMudNgl8lVpDiXi
PrWvXxc8sdxzWuEotiy0CAsrXELFQadS4jaiezASG0OOC6dhL3JE1rdsPzk8k4bJ
vW6A44xjc/Xvx4MGUBJLoQQJbUILJ8Ohof31VUrhW5+7yNvTG5J+bSpDyZ+49TT0
5K4b4xBcT+d2TG1zKz3HX0F8o4m/v9oFyQz11onxMBxHsiIp41fuCfWMZzuUOTJs
XNb+jvyDxuG2cBRfGzLOy3B+Tm36yF11staojvNaENa9eeoCMWGjpyl+LMYiaWYx
aexjJvFpa3/lfNw5pAEaRZcM/fZLvQ/SEbevnBQLjiSkGdU3kGPnX2+ybCEocN+U
gxU40uZmKVPnGdDmZUE8ooDlLQ6dqc7C3FBUUVHceEdQfOzdD0J/Km6EJm8zFI4n
M1ielKHuGmrs0h/pl6D7UNANf8EeEPXJhhRCnJ1RcGdwKWnipfSnCqGRwGO6BKWh
6RoQv4wLAkv7jckmZg0E/8nrEIvFRB5hsqLSNvYwGUUDRGWiBhy5wjSktkpxNHZF
zfJafQBpSKq1DB0uaRLSbM/FM8d6+4eR1LL6LCmZR9XjrL+L9KSHV4C6HMbPYBVk
PSbV02xZ+rX7RV+WCbT1WQbgRpmOClTdHEUFVC0y2dK8brWPvBxdbQQgeNDn9+XV
hp86yvPEDTXNSVE85yv0zbeFP1N0zS3t3SqPNnpJ4IPlr0bP99+oF7whR2u7lYTt
yMuldefmQPoYqHe02nyd9NCnPtlaP6rxG/tuBso3mGhqj3vKVOWswjHidU3FmjZY
iT43KX9MtDyqtH4wFtkbbPKOTfWe06jlNFkjuTmPIsnljPCIBdXd9unu6I0Bz5TD
IxwlKRplQW3gqgWHI3Lcmyw1EIF/TXkOY09HG5ket1HdVYQMhOey5BRCFUvIIjuk
ekGPA13EIQaiOyk1EjYnm2ZBtMzlet1vvtoVRryXJKlFqScraoZq7PFZ0cIVbBG8
MMQacPEEym9K7TJQgjX7k/BFa8ROPXpky1oe6lL75b5ndcCoG+AZoGZKNte0apGd
2aVn43ABWmGyYqpPM8UKiwvJF3JBEzMoQRCEn98IKH1SjpOpBZWPfvp0L5NNOTTH
QuyfV/iMLrgoMt72azF+Ed1c65XgrhYA7xEr2lViLiDkEqHTsdSIm5EU1U5oBl8C
AObn72y6VFSp90QBV5/PdijQqfAkjefrkX+1qOqUzSqHceD8WSBRdqhEhElGsRtq
qI06Fy/ZyY3zWUSLOQnYzMMdcih9K9i2GHPWhZmW9J8HG4SOQAL7y5kAKLclKaQ/
U0G4atckD/8KKRTesI5Mcq9CNF0Cotys8lY7Xu4GdpV4ah2F1g/MpGSrqxWTwaRJ
izVFqZphgQW1jNVA5HftGhmSQnc5FJjxIRLzAwR+4tT/2LAmrdpiS/S4eTG4PiGr
mr0OCIA2B6B2WT2BabBhdEw1DjLecVues0w1HDQaLpGjlmKw9uur8X7rwZt3kryO
kMCkSLBQ4LHDHoxYvyaE+spYUZ1pzI0i/7k+/Em0N3XAvrtcPLO/IzHbv1p1okCy
8XD8fKar+uNqgDpfWumoOz+/KA14vyPgBbGbiEHTs32+T38JEP+zgSdVwnMfgZpL
vNMaa9nXh3ZS8WsHPMcKbpv00PLv/onwOzodD5LkmHDImt6OwMFFTYM6xaY7ZLWR
zOLfYTup9AoR1PweTSbUvmiwQBGgISjd9knefs/nqZ1zEO/bYOCfF7bz5dAufV9A
f+j0PasnqwGy+U7uhgdi0Ae80S8ScNa00PJUbAZ0a82L7QkUEbQdJLG0VHUIzPyw
ihemcTcS0Xv+Ifzk3yRQtGuTuHYRgelNIt0jTO6VtAegpcst1dyihkJxsIb2tPZV
XesOnezwdL49kF/l6so2kPwSzluIdvMb5RRanw04uUab6jwTJx22v/MmNNOWy+gw
IQ3WSX50Bv28jXspieR+IWZQMKXlse87UDuBvfTN8QmQGxrXXBzQuV9Jc0vyjuj2
VFGeMOd+N6iR0+jrvaFPDJiWJ0ugRnQAQqR2JspmUf/Za6SrFvYExRqEBjvEhknL
5b0FqsNlo44N8RZXqAfsfQVvY7OukcAUCB4SB8YglsZSwOBbpu7xrIxwEeezr3ds
9bJJUST5QCqjqkv/njJcJt3IcZmRqLT7s2SdZ42rO6kpGKG9GFcK7SssZIamUsws
Y7ss0y88bjVfdbkLn7L6M7LSc6nDkUF/zeIqmwpBkcdyGtmuxnlDrNVXPvIezTGq
vciYCzT4azjKM6eJYxpgQl4eTKDU21Ott/6sU/myIAny+5C+Zl3gkfLgUNHbubw6
Pw0MVK91iwscCD449XN/dZFVzuK9XtMCvhl5h+joKbe9VFHubCVp7uPLAxM/dWz+
hi3xelqYdS7QZy25Gkl4kuv8uRUR+Ie3JnEPORJhTQvlHjPcwwGz6Y0BXcx9x4sa
9nTAf7E6NTFZ7spP3QxfZwGrRGg88yYvcnqIDBT5SgE83Yns1xlB5mpbXwur7xoK
+yxzEPhKNBbtpDT1embmdrXnrGTIMXLhXY4yQdFO0FFs72o/ghduOoRwkWIUGlbz
KJneGaylyujNDg+yfnb4bcBkhKomYnIjqEOeXSMLzsJPXCUUfczyTf6tZQLpV6xp
qivxYX/BEL7N8pSFzLeXlapsqq5CjFtXRlVjYAuuJza3TI+/SSCvPhOub6yevkHk
iYhKGcvriItozIEKe/IlegrQmyWOj4kPDUADiOCpIJea47JqBQmYc17pGgaOIKLp
Rg4HWqVMDZ1/AnLcAEGcYXhLkGIH7ADxer7ABQlZlBijvlM4FaVumzecn74DbF/V
X15Ij4bjtaATJzSmipp3CNEhC9KbYj2eNoS0EqjIx61V/loxzEI3OIHqq4z89sEY
Zdw6ZHq48J5RZUgNeSFeYUNij8JAGkPmwNVvWRQ1CpbDcx8CpxzWr8t2G19HeUIH
moAFUl5FckqCN1TQR9sMaH6ctcc8u83fEs5xAhWfwkErX2aNGInIGUEZYmzsjJCm
obU5RUxLIP2uSMS5MPuD3bm9qpHelML7HkPy4z3aJM5pJGcLIVLGzWVsf8Zg4Dn+
Sy17RMxutOsendi/wghQhSBCyVgr18M2Eax5K0h9NuTnUe+8gsVdwoUKxH969vsC
wYAYQVIEbmcjXr+PnIEplQbRXlZU7wBow8+Bwg/QfuCeJRLf6AXh9ZPIFds5H1SR
s7Mc0QT0FobeKoStFqKxwqgv0EyWX3j7kx7pZedWGoTgmIe244n05V3dyUi7/rfs
WaZws66Laf/p0Z/CrvCtzt4M9UT3U9oCJFfJfQzY+dNKp+i00VRU7jmg2i7PDZJG
rIhB2lJ5ohVEyrmMxhhLGdIQR+kp/irL93dsD8rI8/1uka0Wl0cnXqfNzVFxXSRp
jGjn5cez36C2P7qf0LCuNzsIBMdZUYBa1INhGGRenlU7Th+I9Xufn8408UciaHrm
Lh6qb9su4fjiJaENffJIQRWjQqHM3OsDaIrfmj88/fybpLy3Q5ULWWCrUBtkjNKP
bXq/3hcHjfRIG3bZTVoPOowANRp4gsMYo6FeF2XIVs/wjcUeQrO6LLRRhI6Asfhw
LmvktyRIH6J/T6ocej/otfuSRkN2EBkTS4inLAJtbI+ImBl++7A0JAc43fif/5WA
IspSjM2QEpg+fpDoe0WTTP4G4aW/y8dV2jo4p7mbyULc64OFapHyQ0K6U8IQr5aU
QBiZpzGL1O+Ty9y9Pvfersd3zLT2ZTWWTDQfhrFcLGoi5z8hlnhIFuiw9fJ/iBX4
IhWQF0itYVNeDEKHn41mXIEnMgEWvn6zCDVTCJKEHmHcvD9i+/xpWwpBQ5s95rIG
IPpjcGVaz2I8i5Ztgu4dBZzw0q5thFIhh3soPqTgE1O4MoSf8q/rvZKjPC3O2wPR
urGGZlvydlBYZZftm2uBsqVtbLfJV4abBs8228LYi9Zb6OEMLooZYLpv3bCGFuVC
2T98vH1n1o100LXste1TODZSEIUxNJ7ctgdndRQjrXD4RSkjws1b+FKYnRWJr9Wg
H4kc5KM7Apa+2n0LZT+GnBenlH90HEDqayVhqiYzQMnwSrW8ZVaM5t1nARl5qeNz
zZ4ZfiuAJfTzm64ndkBM+2dvG1hcgw6+i6y2baTrJa3v2bl0DQWAo/UZ4pvwFlvm
85iU0q/rRK13ppOLFkqND6thOAHvp2o7EFNyp+PTw2a24OsoiJxW60OMlmjJnqnm
AUfHT3tFFULy0Ji788XcFhC23Kae09t4E6KPNF/zZISJB4fQrEnQvJB6VHGbKjst
MhpmcMf6NtDbGpUCKEGbLQI7n2dgUWXQ7FWTRDWzhw8NxJWubsPc91cYVqoU5Yt8
acb8YirWbnkxEnx36/aAQlIYOKqo3pAdhA5km/rcB9d7+zODJAfVkd/7qRQrHcpf
PuL/niki1xWSlQENuPoF/dY46mfUccF34qg+Y1xHoys6nCbKhATcZmlFeNMiGxXq
9MPfDxM56mV1kfz8NJMxyhhjyOHcO8BUJXnuvfat7A+Rr6jfp8u0PFRdOHpLmCn9
pOENW6xHYtb+fxz1bR/yY9XOMr7OCWvFx+T0osdt1P5XnlxGp57Jfiy2e1ib5WlT
eJdKMUDUw+Kg2SG53YQh5xpqVv4VCj5YBGO8iTXQ9Ybb/XDLN/tRQsDRDZw96Mbb
vVlk5BwaYTBA7N7A5dBNEBNYVIiueAkgK9Jd+gbYQM6/TqLOVHoQFk9kJ4VDLPPA
sU8zgUhKWjSmiofXhbX2S4PuE5gmlBu8CCHBERUOkH1eM6xXpiibBuv1kHcBq289
I7nJU+r4GDp4YuoUmn5UwTQuF7SCJw+5CG0VPdy7+/607F9fxGfFNM4Phj8n4ae5
Jspar62ko0oRFWR/6A72lNtG6eZwPZEyoVQzqho/aT/tCuhCezfdB4DjLE1SGi8c
T6G8nu5fPxvyfXCHvzFz3c0VMEZ0d8APkYhpLQ1pQpjMwmaAqGin0l+OaFlq9HXi
OohxQLJCsxQ8R/4nDcDH0ZGIDsnJYL2HQnnr80v2OjgRTWMmPP3dZLrBoB8vi9wL
CTsqx/uzqvp4bauW9mIzgG/f/vPRY8FOjNn7aXIOo/jzFQPf2iVbwhCMFY3qUfod
f7c3+XLPYzY7/fQZEEjkxrmq94yM6v0u3iCPpbq5YbLc6CfhH8J7DzRQdKM0k087
JgFFjiaQC1MO45GZupHXGwyclI1Rh69IGmPLruqsdlbULGGTBdvRZdH0wYwJbgjA
EFapVEgJ6GhcNSbkA3IdyszcohXWXDWXaqhYHjP0Biq7etgXC1vAqdcgBHjxsaMH
yDQp/kYFIPk0Ht4jAHR0F35+PDdNMoRRTZ5fcSJ6B2z3hB6ZBWVr3uXDsgS4G0Ta
sSKttaKJI6m7GZQRtt+U/k2bR/VcvQ+F/cfr1heQK3/Jl4P10BZ8WIOd2wWHa4dz
pdEQZSbv7CNqSY7/htiSoDuI4i1DlpwprWKFHbZJfMzhIwBqz3HrgbMOY6bq30ID
nMbLo2wy8Y2nkjuqn6MDb7SBlLdYelQ2tJ8i0XjP+WjPnDIKHsBN/N26XEjv7nGD
x9n0iXS2TRMy/FfLPlNbUxk3OiZwvDmtVua+ERXQ7DvX4pOVsbJmTqkvSCErtY2l
599WhSA5k9TEfW+CTcAoFjnKq5S/SdgW7ua+RkVTuV135tMHBWOHxmd2NtUgK9G9
oAQlBKXKA4SYMhWlrodc2TR8f5TTHPEuiCLYvssQIlJg6KnVCylCw9U6y09NNOot
v83xrtcXkSrcCEUZpvoV0CdVItSj+IbE21ds61KdUvm7Q2CXA8qrMaL38qy6aMon
DrAxfAvl6m3qiuJRskW9vtE6lo8inANclouyp58OlGIPHg2GiBmEJpkEczCoSUGU
5e/FE9pn4jH/S0/j5rGTSVBSA+3XbjkQNauboo9ZnAam2PKr8uclP7f7Ul1EeuSd
RwcHwqAQ9whpLadX1vobnzq1XRbAVE3AXXhVY7Qvewtydz6+fWAQW6Y8p5mEtB0W
Hus0HjtlsnuFHVKESJ5cVYwaUYmEkBlMvBidXYqYLEhuiyIZbT/08nX5aYDONukX
ErxHl6fDuJw2oubvy4d7D+sxAg91xrDyhNB/SGZ+O7cj4o9ZSbHPM3yrko9KEXNK
7deSbm79UbeXDO7kjRbSaTLc4xw2sgZu2gnXMk2DLhA+jV1T5ES+fw6SMNuic6Kk
sxkCPxHz4HZML7q9LCg/slRviPtjSLaHOUBytXBjJrY6cD/5+fhsR752urHzKQd/
cAWN7nj+nysCVKmIVMgM2pc9k/PNqiJ8lFyDGe4UDXBFPZZUs8cFvPK1xYEuu8AD
f3HqYm9KUAyxO6+duj5J7LQNeipxltt+bpKKlu5PQ6SEUOmpM/mkdfC7cFq5nPaS
5sQ9pZsVzVWvpagL/s1nmPlGWtknQiOv3tdOnZdTRl5TpZdNDXXBIl698xv3EIZm
vojURqQHuW1OvYZaCm3/2ybeLzI+DwEc/iZ7QM7r/45OodMCXKwCP15kf15tM8Z+
Ra2OqzlAG8+dMMqIZtSd2q4/5wj8gvNJPKlip54Rppa/Ri7opMZKE+S7BOHsc8OF
X099sUZKo1lG0F76NksmhpXdsVtrup16yEma8Rxpaopqram4rbAhXtTdQx3ZhCSj
04/eha5nuXyN5Rqagr/ALLG+KtnNyoZCm9HB9gGgAUbufpUk8qz2aW9HQ/vgvv38
M0fTYO+hN0VdmHgRJUMjhoqsmi6NGKNDdHoWIBPcZx9LGvwEinGiFEdSIVUMju63
jpDDLnxwBYbpqktScEB/K4M+sm/dsaAokDL8p0ZWcTOzVpH9INxYbs1YgTTTZMZf
76VLzeTULbggZH/yH6bGe2RsHb1K1wdzrmMhQj2u2gG5TqL4jqSeKozwMMCVLjGr
rkEiY9UzAd2gpwIKhKUDXUefBYuXoY4n1QeldExAzDzxIqqDhTLrfmuxC2EyYXZt
QCVeRqM4MBUvjb3xuCtXkk1xBHq/YQd0Sm2ULdMzaLrKgNaXn1JvxDBrHebL8Bn9
qPgU/uuchODMqcFYweIYe6XXeNreIf7YOJdEhtcoXz13QhRcVMqWZOnnASxECr0F
3HWBwPSA+dONZ32OIBbtG0JJKuaDn5xQErIPZVGmC9ph1gvaVZUXnaroEEkvIXB6
eE0/M7IWBhO7MaUMy4blMOdzkSM6KirYGpqlkh8NOuCZ5kMrwiBKEZCFUQEu/LAo
BRACeph1IcRRS4o9Ya6Xz+XHV3L47O3qL0/HqJywQhgHaM1xKsdJAOdaxh6GzGaj
3M2mqccMjgu2jIXCGMI+qsGT5uEMCTgFk98q/Ses47heNQFyt2EZ4H5M52fwz+vs
USjNg0VUHNseKBRAuVqjsHKhEpxFWG1573lGmrpE/Igl+6HO4s+2bDkObwnXkSqe
F+wDCDN/rF+ZjhAbH3S2hk2lMjeShjQSRdj0xeO2j2aaCcEomlrQn/ywCTCdcqPQ
ZL56XG49g167/Og5mJvlcvwFl/CXAXSYZKa4bS25EMB+OSx9q3jTydDkX1NVAdFB
cNlI/yVEjGw9+KS6GjvDtJpbg5XiovQ8OOuceGk3cnNP2Tbb6HSY0WOqewS3pUUJ
DQmEmC/P7O+SfMw96TP+HEAugHPKzhRlZeBZOU9YtLZBej9Sswa3UZGGetTpexUo
oYEAfr76KkMrsB8Ge29weHPqe2OgwwTdLXUoFk18/4DneS0H/J9ZvZtZZB7esb4H
3NfnHZEDzm5/O5ZRn63Dy3wk4NCA2p80Hnanujlba/HxcneA1NTh9QB+90ikm1cG
4c40TA2fvUKqUxUyTWad3c/x9zq80VydHjnMNKpqpALESuSEKZdt0dRgLCdQ5Wh8
fjoj92yBRWb++xT6GnmetRAnUT80D88VXXk/Ex2sNwTm0kkgNn0BAxEoO34QKSok
ymlS9Bn8zmvMoDsKQw8X+uhGtfcpbEKH4vyPozqhiN0rRAWXArEx9yB/rOWolpHg
VYWAEwUK4AVocjLhM1lK/eRylQOxDT5yUrTvYfjke3WLh5EAgljuig8mv2Y4CMCW
FPQrKkAbUWhE5uD1a02YNrxQmzME4Rzv4Rl8Mua3JQcToM4yAHIQn8qFiI+h9UI5
lHDDnd5cxWZkAI6l9yw65aYaehJZNIs9ZksqKZSo/OhjdBQY4O6ydGozph3TYTGt
+xIEjmY4bJHv1aaKL8mZ7L/FQ6EMY8Re1WF7M6cKFUWvOuU8AI/jWf/VLtsuf3F4
ahCvoaFitg8NthQiKM5OgJlJRWIW6PG3ILDbe0N3+8hbveGjpl2ATJnDqnURW6KF
Ytg4j6C7ZlbCDU4D1ZmzgwJpPNakv2MZF/o5s8capmLPcuM4FdZKo6FDKVBFG/QV
+DFeqKrjc/aWKMcsyjiha0JkADKQLZWZnKLEvGsORbEAHYOxTcyLonG6rTWtXJv2
WW5JHWCMrL9A3T6XiQfjs/klNf3ZMhbVlHGfPiGJd3JH9J9KXwUhLs2GsGUrHAey
NB4EQF+86B+VfeCgcvdjcBkZIBbd77rgXvoWqBF2z468WFX5raTQfxH1w4zsVqsQ
9lTvTzB0hYnvKBCpai0liJeEoWwmpMcsb/ALgIFjQjpykPC1F1soSaNZ8CUWBYiF
NrqQ/S+CjQ412mr11ohjZa6jNUQaydzWXQXCdscC0J+0WK+EUTjO2pkWjhnvdzd5
WrXpANeJFX/QKEE9AxhvOKXxULD+agPAekmbsoOLJP0XqbAHNoMos16hPxmyUJgg
76LDpJMvxEuC/uLKhwtZpJ/LIR7xmhAGNWHde3fVob9r3nydE2ra6P5Voagn+42Y
UZTzltYiNwPR/TWb6fU6DCkBtvCYgxadj1viWQL15d/iFkMPYLY73HSUMb8/2hb0
agwoZR6zkyeNKoS1GlRl/yPYi+/vitQwuIUjcN6Yvm7GQ1xP0Nj5KhIdu4Pe/2dZ
2OLgS/muq0VnOt/+BoBqxljd0qMU0SFCGGHxl45FtP3BSZ1UC1wokkNR1OnE6/6y
IPrW91mOCTk+qStLuimCd37X4qqLRRVp/pAWbhi6eEpp8vZ4HB1QIeNkO8w8tNCY
bzautw3keEE7GmPXxgcGvRNDxw2UjtmF/W9+M5TmEBRP6/UfDdol45lAID+hTS3I
xV7CvnGiTGchUmxH6RNXIHFZDfkXcpnEBCkzXVpAu3EEp6SEUGKxQXMj/Dk9m3qP
BZl7BSlTQU7NeizEpirUnEhgLPkrGAUxlCG48fWJMJl2Zdaz+LYV/CfE9mv8x3hH
5UHDdkzlSwffUYSK4alFiEqTpfsQb296Fx1PjS6Q8vgoaOBXbdo1XcaVT72Vui9y
CL8wqMUNz1AHTimtg6Jc5a5uEHS6Yj+SvILeIGNYvqMpEAQz+3tVsf7R3WMTJTk3
mtqfV77tzaP2+NOCnZyRCEKIZsxdkLzdatrY1AWpUdPMZGnG+KAz+Mpoo2V7XLJp
9H/k9crgM8y2k/MPf7tYu03xZIeF7KFkpmnAQYrqVcCEiYZUnLwvAFrM0qYi8hBa
tMwekkLlnujMvbfQFaTOZ5RMivUtDmhz4tozhWEuYDJy6ExyzsFQxwQzVlRBs+oA
2U/LgAAibCWc2rxDfffaqk1ymhWv6pwwLOe3E2jsiVYh9jw3+0rvvujdXap6h/3U
J3N6+HXnKDmZTNYeKBQgiUEsGAm5cREefv3QvWcfRlJ7jXzASiA+iOscnJZcE1D0
C01B08HjC6jo1d6ZllngclhHffJDvEOCpsG1KP/2vbF36SW1QkjH21CuakuU5Rd2
+J+N/5t+PXpKfGS99D0s3VlwlV4bGKcj8/wKDc1cVvBSkykmAzs+MHeE029Mjh0m
uy5vIexvZisSHoCgun/eit7o5lFtKbxsabS7LDaJYlj+3ckPDOm3gijtKjFKx2fj
x0EhdwDJdY/nrAwPWDsciGTCtaQZ8gic56iN6HG3y5OS1jVQ7G4vb/AtwJctbCoK
OEeu7oC2+ahZ87qbcUB9gYnCQgxSv+0CrAKAu9a5Uj9dDwsIIwRH9qKpR+NSo13n
upoTnDy9IQpBxG/ubxV260oKLc9Zm9IKFrzobNoprYF+stlAvcpHhajM8r64u8ql
G8m8P1j/siBH+vAKMct/zr0HLHTm17rVPY/iFA5VSvQ7lnVcCBcQ3ipFRxLTSLDN
t75PIHxDf8lrtwCmnood4yODVkPs6YZ+UrEGOmBMyOnd0W06sCqFNdJGwyi+veey
w2bTvqlUnBjtn1LDjZU67zFUekRxPV4sJM7jwjfJ3M1PwV/dqBRQiGUQhhA6tdon
uT7zuAmMzP+ZDQhgpdYfcN4jrp8FpViclnSiobU9Mc9iuVEMUg1DDW1s7dC5N7ln
c0WICAg4hwHUWWev+ToJIC+qLhjTl66yiC28ioiPJiLcF+JqK+xRbrWiGQZ3W1QK
pBZ1NnZN34tuHy3tnCXCy2zSdB5TP3hljk8n6aC7v1TxXDUQwrNDqBjnZ+QbjfzF
X3vFKGceBGtBJu6W3K9K/Pllz5rXb6cHktjxgvlehlcJG9UhiZ9Jiup9M3WinZBM
KlO12Zya9heEZnBDQZKLw3I2xcVmkkqxczoUZoTaWoV+M2eChPOckn5gax/g49mu
z5/HyXoyirWdwPEsOPXj5sFMND0nDPd9elFTGtbJzrdWDAu9xkNPFi5y3znW2rVI
u4bQpK9wq76hxlvTd5FQsF24p2hXxsyTVlCyLOlpdIc1O3tNQCLbiMsBMtBfskjw
F4lNTYTwZdbhSbfVHmVAUcMrlJGiIKpp7KLDevp5rZ9dYCTzJkolkUEgKq203uyD
q8tx7NImHM9UwxvCuSlFAaqQisdxHk0p6zF3nkVKlglHmCoO0rqYD30LNvgFpMUS
uPVfK0dmshrtRBibhXzAbXV+mnHKpWjbjrFNb5OpQmmJG8YB1aQTGO94ofmP6dxB
tmsvfsKTejmrWRJgYVabTEhtDSLRUc6hGbV9f50JKnyAX9QqJ1FQdhoEvxiQPHdk
hDo60z1KoB6BY1coZDG7bEhA89Unu+NggGOMfPD9zHd8ZSilw1GrAvx7ORl2inAn
LufPD2y4FyyTmTDnrW3bFde6la/Zpllf4/we9qB4QnHdYv8tIiT8Wmd8BnxEVouP
Xn4b7IwSJhYaU4jIn/DHvXaoaWWc05JnDMy+5DeiGGPHjJdJLVIeYs72BBO6BJlV
r4wD4rk9kRRk3GmbroPs0PPqMVVf6LJplHfefK+hHr7Daaawv9Q753RidCm2SYYs
W8BpsXncpNkXib1SLnJS/1L/Hps1RGDGl8kp9SiZElaLfRm+O65Dl7adqPoS48dK
eUNqqs667c5v3Fsx3c/SsYMQbxYf5a6h2E608PeykIM=
`protect END_PROTECTED
