`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hFN4muNztO7Nc08bfuF2E+2nsDJ5qI5bwlej8GCA85U/2D1vg5N2/+Eiuv8dLdUi
iaODIU6riaTOTJAYOjxiFpNLfiSlsWp6H7pjv3r8wLeZaVdiTrACrWv4KdBp9dZQ
fOn6dq1BENfEyFQTmGcwgIPDhgxQNS6ApvUfQXR5tLXzZE4P1jlTLvseP5EB9TU1
AOOyWVttbFK6sxbQSy7fsp0MZNG52CCAqV7gAeuPPRaV8FMJzFL0Do1NwPNakEPY
L7ZuBk7VYu5J/3JoMYhoJ66WtckIoLyrW3eCxbZYaVLmiHAp+NP3tNTSb5GWPMPk
dRWOCGEIhj4blpc9PBkoFGdKkrSBgL/1dc1NP6txr+poxKVUM4yOie34DTgwBLDT
BUyeqRFUh5ULMjZwbzc7Er3uVhH85XHAVS1Rg0BUZG2dl76rq849KKMm++/o/vbq
Ttoc72DZMZ4Qqov6BHfMgQ==
`protect END_PROTECTED
