`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mxtU9afd8ANEvXfy1ZIIvAWUvUy8yR8Nu67qEhYVIfYtFpGwvyWdPg24eTEd7DWi
/Z4aaZsuDcy9btKrMwTXqL7kqdRml2bcK63E6PYLDCZOLOLqEmi/yYRfOOyyH5Ve
fms/+vpe9MPheZOMf/hs10cJNBwxrxvD316raa7WJPeQAB+1s/g0rhCHzyvqn4sz
seXHZVK4r8bm+qp7sHGxeOgubToxyksdjcjUhqY5ZQT3zPVTMbB7DVPFNl50Ow0K
c0aFzekV0vG2j6zP2RSz37B03Jtr6UwDqMGSkplrxvlOfNzw++iJOlIfxU7uTj2C
bkr6MBT/FMYI6n3FrBbRM+/Vr+GLDU2jBL57M9ByTfqX46WlAV6j/w62oSF/07MD
WafRNdMb99ptcCR8gpkYsCpA0poAtfC67xarmXiFnk0JQOFX3DTh69zkA4pozhx+
3sAlPf62j6hldqS5C4Rf4If59PAgzIoYhEW+fCDW2eQLGH5pF7pqTxPR3gq4d3R5
Pi4AIgPWxn0qmFpTBbQKB27DLfBIY1np69hNGsxqyD89OIAMwn/vVwgp01nuHR8y
L7ir96HRPw+8Q/aep3Tmq8bc/1GKOk6aChtMaYZ/w6gHjaqJQt19tYVoSTQNwZcq
1H9+BZOdHIjJlpMaP7D6akvwP4QSzh7zRD2lMrFu30DPb81V8hmXIyZE80TVRvEk
U/MAR6Tu+guaWVTKQdDR+buCCBhe7TeCPjhAl/WnWK1A9ps1I3BpyYBIALvfDOLw
psXkFbx21aEOOmhCjt4DrrRXij+fivoFw+tAYbEVO7gKpxL7YkZygKpbb4Tg0FiE
dcBxHLD6uAARac1igHSL9VHLOMK5GUGfKroEhqUD41mUARrX6jOJ+aRKmyZwlLS8
NYWhjeeAbtVKiQ0IFpZ3nY7yTm6uD7dGh0pMnqyjm3eCnOLI2+4MxaFq7+W2uChP
af1kaBn/HzTA7f9XqncSmmLsvpXdAs59R7bxPCFQng/pXXNRABL76dayhSrt7T4s
S/K4f0yV/JU6Hl+oUxBRUOU+7pTcumJ08Ry6ziBMLxBCICt+9pj1c4wesoEAwHbi
TRdzz+vPdbOTQWLbPTwdEvhiGsB1/4T+ngr4aLmB7T3wDLKGo3t5sAy7plTAgAnA
cnO/o1Zf3CvFFwb3qvOpo8aUqQ+HS8ek74LbtVJghXg5EwT3iO/n5CXahn7Ql0IP
SceD68GQwYOyONPvUyg3D14gwRHkfPorMCWw8GyF/eUwKxvjrs1NkWy3MDZn74zb
RNUchJnTz6BwKQwhzjWt3DbYJp9YK4WD5OmNs7usLxGm4bIE6SZL58m/Aieusui9
YeqgAVox/KcDhmVu5B1swyfIYM/H/tw/QPy1NPylSzC8c6xE9lDx4Q+izqO6IPcs
3bmVK2cmOeXLrtvGVarUmi/zNNM0rhbdfIgBWZ9CPRCDRcsBlhWjs8iQUbPv6uuz
/lwVf35pLgWWSFzdVieqYgnBDS71ZNqGH4xYFmV9aFuKNvarBSPoPKsk3x/TA40z
07lGB0Cp5Q/MwfyZG3HyzBD7giX3nyWyTkUTQ0M2ANih8CgMtsJ5clx/YIi7RUtf
ApOA2GBRx3vD0uxFr9OGRMlKIY9JHByBlCeZzQXAoRF4bJrM3bnLLXJTqp4wIPQF
vTErE3dHKZi+P7liMyTwH7ZM6+E0a4S0eRhEr1Wtndw8POvPkTwNoIsz3wwH1L3Y
GaiAishs6/6h2wHyZmEzs0bZYD4lhfq0V/dJpU6jW9hId4m5TReTgm7WWIZTGiop
XFAivcIEx8qa97GiDWzYIyZRccn5qrIOA6QjQ1zCcsuFFdLLs9MkSI8jO0dmv9vN
muNRU3hyYyvdAHVbf3zEciFT/4YomXahORlq4SfhbgcFH/GBndOVXM9goanC4z26
0jpiG+YmRYrYfRNHV8ErCGWJwZXq+GJKnQqQdnyZnzJCwwfj7o/ZCY/yLyh9JtVC
O4NHHVFQuAn9IkFGXk4ZhfMy6OfzeU+rC2/PBZe5fJoEr94CldLrmieOVr+/biPY
Efrcpn+56/MbE8Q7Iuh22lz9G2QyDR73VEeMfzxOC1rgW9OZecE9KdaaIzT6s2pX
uOVOc83RhSkhBP97rPeWW0+cN48sLHyN7108KkVCKA5XoPaGBjfUb6lQjFrR1/tL
hrmtg70io8rUev5uJE+YPNBNw60BNifdMe6Qq2auRbvDlSv/tf9Oo1t0hYIGQ6lL
v7MIcyCDgV8EO/jwa0Tte0vqwVbJaqxao5f0cKecyN5iupwtkrW2z7sZ3/uQuzEf
7daacC8vmLya55lkpyZPAkeZJuK3aJtbU5sr1SLIBrt/DnG+1IiophsSRjc8kZs1
eAgm0SWkL+Zyv+ZQKmjYDEjUe3VyvtR3lMlD5XEQZOyMNOV+aTfGi1An5IEi+Ob/
D8qeRt385bQsdqB+41R08zNCMLNADxpNLv8c3m6sJa2zBsvxZnXc2bjEsQV20WiR
Knx8/AEQax1IuzXFvbBOGk1Ni6SfnpCETWQYlsEiWHqiHUUSXZb9czkMSjuc9xkM
1aX6wDlcIzsDidKXFmfYpHfHLa+OjVLIPU2VFy3z6/SnGSGhl9HcV10CFylaW6pC
zX9jZR+yvSKV+uxOm/pSyiM1a0nFHuQgm4Hqo8Apko1lzrUbCqhfM+ysVvPV3J65
sICcCGGWmTF5xO0+zHJswgvQCWx92EZLnYlGn5pur+KYWmTiQgbL0HutcD0p5q76
ODjCnpkqL7VK67Ys/7MKA3VdYznXsVCffY9LXrPKMHG8ahXHoHFPora9IbNivobZ
c3wIwWvi8ddAgTMutcvW0kn67zEFvHRqfPCJS9ydbBdOR0Ko7ofuNNGX+Qgjj+fC
QszjUZ+zVszn34W4J/ryUZmCby84phmH16BPVP0Ni4e42bxf3zC7HCZA3/15AbXc
F4ga5ZDtNuL2eleDUZxKlvXWoalg5ULZUmMDdATJX8ddPv/I5hZZkn/GG8YbdyWS
ymxepaHDoY6ikA6ArQRxush4eFTBeYSbLTfZX40W/Zb/jHFEip6g9gfdYLST1ig7
TbTzJfHVQiMuKo71pRXmYgBfGyxor0hmq7x/kO+jEyiY1tQNAH5lxi5W/d61zZdy
ta3xPwnTPfQwa1BtNzC7oF47VvifWVNDcccteS+KdHMvYSpjrGYV9l2pJfB2pVU1
5zSTUCem0pPiI7hWXRQR+mlB+dJVAqYqK2jcePNrkDaq7PjTmKtfXiNDCUfxVHFf
ROB9lqsvghALejhPrPySc/kVJuyYZ+lf4owbLqExEGXwOIGvZuXWqFm6kYH9nhjh
uBjuM+WZbnd5dabXazr/5lk/7ylQ88zAdT07SL9/NlCX8+xCD5fZI0az4P3e4TLc
ORN0dzfGyJf21trM/YGNfa1GRT1h2SENSPmfmZkQb83Xdz5TlmiAYrinSRhWO/DX
Zpx5N0n74seBK7/550MM+hK5mq07LdUpjGIQ1P4id17Ujo4hI/uY1vQpigochbAp
fFKkqSIlA8zMlG53GTojRhjwQElGx3WactsK7a1ArHM8aCznDL72DyrleyBcavMJ
7QU0tGcoERSeVRJ0S45ydCMIxK+j7A1yC+7ch+r9OyiVHY3ElMJdKObDM7196orB
fvRHfqiaVpT5hJov/OYo2+xsTA58qvygAKjMex8mn0Okda6gvO4wW4gb/fZ52fu8
MWPz4H706Mr6Rk0LUj2uzYB94okV8h4mcRNKWAHbzvIO98QfowL1ZxnLza8cAe4e
6auJpRq2VYegkYQrKYAhy/Sfhhy+oxeqyuQnaJ0HfM+4mujkszs/1bxdqCO1Ti44
8ejBxt6zvbhFmuN9OLCR7YXZfaI3pR1IsG0ZEZCVO8Oc44WjLVo+KqfsE3pZkLGY
97Y8RDWsH0X//qvQIsw3VDt/SwuAeO+k6i2FagDXiZK62Y1ZPW4rLMGwkI1TzI0Y
QHNAnUWQh/RJgRbAI6tTNP9Ep5aWMCtBklqkSUN/vvUL7lZjyhCNQ+kkbFhVr3um
No3c6faRAeBvXFMVLwNPlNkOYokagP/uSmbJawkz2S+MiacD4eZZNLISTC2sG70C
FhiZrDRdruD3BwIoXBKbpi5YyixxfRTzrNeuBM+Tyt7UmYDcVx2p0wG7ZYRf/2sn
k57Ha55DCO3EukRkDu/v2zPhIAzbziwu/mnXnz8DLEHB1fYwghQ+wL6+78uW37yw
ti3bscjU38w0ueiFzirgKDrPumNj5+drnWRCyu9qrZ7uP7gPzJqd1mBfmDVX4QwJ
H2XFaBbF6oTR0nn3J5hIcHdtzNKy10+c9k3SXJRv7qC8+2wf88jjDcMd1lM96gdx
HdfPe4Wj2AL2g+iWCMf9HTuHgyaXs7P6rXSECnwSomUMCHjP9kPNTUv9DES5pE6Y
vUMbgRS9XPyY6uekAEblkg9/MmJHOqwkikN6H5+r45WYiSoQQ7UUjJfjLKs58+AL
bxhC5nnyoyPW+UOcSRvaOBsO8NPNAcwcAV8Up9G+Zgjx1aGCaE6fWyZNFJGisnDq
XoOfJFjD82Ts87HAFc/2J9r5tXRaQRfpTUwa3Dh2uO74kY8lH5ZaDWzJOOWIk0jd
`protect END_PROTECTED
