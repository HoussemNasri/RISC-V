`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/X6nDNMU6NGG3MPSnWR84XZm1N4U3bJq3UN+eGbex0FRfcX9ot97HnWbg/+rtVO
p+1L7IM3f67MKLSS5E0qYzTgnifSW4qVE+VRCRznk7si9+INZBHNSsyJOJ75FwvW
5dgs7Zh2N4atpKDQN7Kq9CmdUSQx0t3Gy/h6YQm/62UAAl8wXCCJ1si2Ih6V1tEL
pm4tgzf6MxqKED0aF1hRyKXPxX7Yrgg+juIkSFbFBfsyyx49gct/XM/P3FWDLHfU
+l6465k9c+89AkrvDz0d66PR5IveBqHmbJk2MpZ6g+jokrt5w0OhUmkJtDJtdiWs
4KEYDPUol/3/trJUT5yf4GPzTYuk9h2IwgSBKdGF3x2ONpAodJZ0OErbuH/jAjzY
H5nS+byqDXPQnuaPQBtWHt3SSg9MkdQS7Ba25xUGfuNkL1fUHC9TF0I3wUl6bgpB
1w61KPWaHS74ZWx/QyjOSHKop7/op3gNivYb/tno/RnQj1t5rfoPYdkXMecogT9l
roRCEJS29zdCH3/qpir6WN5dWXPvEolvnkWZ+fpzPWy9UDU81hSjo5Mvq7rMkgSw
msWnOVk9PfdGfP59Fy6LBgAc25WvkmM1jOIBXAecPiRyNZmNpwuDGzvi89TsyuOa
TuLtFyK3294vcDMgCYG/aDP6VZjCUD4knVrN+sWqizQoJiWiStXj5houj9ce4omh
vXKPW3Ag//bQEOMK3NSfhisyKt4vHKvlH13DG3VLZrCmPJtbxlVLaZSSr2gWXpce
qEFeeDNdsqRbg7pQdwnFnfiZJ6t0Ta7UCo70T/8dHpV29Pt/mPk0VDpixo4IAJCu
o7wzPpHPK8UkpzBfUKlLwkBphJF0bNCkO6qpliVJRRVYKpyhgltQEC4O6g0aX99e
wyB0lFF6K4RvS2XKAfwH9YkOqfMoUpQv6qPi6nqZBC8JfbUaT0EFu2XBaFe1tgBm
O4I+6ewtBg0bx2egeq1+Inv0IgrEnadFI8eZH19YtBZFwzLXK01YQFVSVTEwY23d
wJ4L70V/O1FUQX/cLgO3nuza35pq0/VjqTzv+tobLbJMArZ6ipENpxhMRIom65B5
O8O8WW2pfLsxMa3YO71lD26WhkGAjh0fpLAUNp/uw9e68XB8o6DVbHRv/ZEZ0B/4
YxneBxsBNMqCGIXbiN/owz2S0YJFTmWR/ez4E/EEjzqAtsP0kPgSCU7ro3VdusZs
0m3H8H+MnqUBXNquSVB3XoMp++ykQkVgnzaufVRa/pSpXzgB2PZDRxFavgshJ5sw
rMYsmqawSykGIVNMZ5aO/388xwIePLDgfblT0/sOyBmQJR/9YnE77flQrNag1kwu
A3k1ypglXDKJnD62Q4iX9nhOqK7NJ7Hwr6few4SvPFrXwi+b1rlrcraEP3pWCgLv
iK9NsxLJdaZAb7xvYLmiyIC+Db7uPSwNEfaXsP1ldUNJf58koqGl6GnCmWldEahW
zs4BO/Z3wi2OPl7YEqe78c90BrZIg7ldIwgGuvtVXoFQGFc49oTOLhGIc6lK33kf
v9xHVS+5T/35/rR8GytuGT/9TKs4i4y9lNg7/8aeHa8p9I0TyiB2WgHinNohTsa8
zWFzPh5cWOat4sKtLcSsHZvizGebMPt4kEUZYMy6g0kr9wWp/uejp4k5Whsede5r
JAesOuHX6hDEwYigz+eFzn6WFfnawF+vibirMqlBIbRhoUenKzGfpNIp4uIl0vNw
aroaN4V9UdLLFZ9/T36Gy6ZJb/e7uNrx4M6Teowq9JYDu0pIMH6yqCxXH798iJbY
Tp5iY30g8BCPrwHuoWTMmPF4DFm76+vofT9vCeR/vu8zR66SXvc/DjDRXbA5C8yU
L/zD12wMsUI4xrZUFIqTDFHOyYuZyY750bRa/3ebdmucSM2iQn55q7j4t7BZZu31
SOT3hnRGeO6z7F9WbwgfnyE8aHjTVl3KwEreorQ1wwfIqs2nXUgTK9/GaOYezViX
7/qNfsBqSm1NtEsu+CLSwO1xd8Ee/7LIHVuI/SvfjVqlhhFDVMmEcvzcuO+JXn6e
929ygYoGHrfYA4FRcp0w2IsazJfcjFnu4z7WbO9rlWdkMg1lYXko7bXYItfCczjA
20zvYTAoqgYVcJCDQLHoejTLwcE++ozcGx8PKRddnUUvatrAHB8bknQo1wU1txWs
rVffdD9d8SouDz8zS1/azLIWSnnhDeqxOBHDB3LLwKfFRIz8QydDKyiT8yqnlIX2
fGotTuVbK7nqLgaUghCUDfeK0ssk2hjs8cLxC9zlHvfS9ngQSmH2L/+q0rnrcEfg
NyS+6RbwiWXkMcRSjeo6nlsQtrWbynKC2yuLxYpty/8fStcuMDaQKYGXzEfOMFeO
R+qt41Seh1+HYFStIDrDIIHvSyZ15sAr2XPQyJuWQHStMWk+TP8o3jWdPoCignQl
t/q581LYjh0MzF0gWp0XIcFK3vOaOvxzkyhDEjC3Bv3Hp8o2GwSdLigP6Jto98J7
XaCeUIVr1V1+v/pBaL6QpfxoffAyNWbXJ0LKFpmLRqV4tU8G0pJ3sz3QcMmALain
1Yeu27oZ9KiEXXoQRAvS3aODP8p3u5PhBt+LKDJDoGoS5Hjkf2+XIpZtPDGZOFPi
egrJcRn+XPeLIe46viRShJ/NmEeS2FJlxziyAguCpPuDE5Vfjq78JNPfjYzGTaMv
N9cViQIN8F4Ms3IZmsGtlK2biECCGVaQ74Z6u2QDaLQDl+FxCgvoMf3VCuv1+seW
HTIye8WOHU4Q32mPklVPchgpHhCSRGPX78GeHYuyZmDv999KHXg72/9BUQ0LF9hU
P+e3gtX+S91DiTKXYBnzi25qbmWSNgLsa/DXa1S7PH0ZIvPcDBTdSUfHENTkXxqB
l4/o9zousQHqPFTYNPz5K4a+81UJMHfbJbN71WRrw3OR9GVj2VqVM1y39gCtIC21
JjvB/3xxSqq+QQSH3v2w0d7Gn7UWJ3BC7GcTXhYxpeFpNg8PsdLLsawh4vEH70c4
IdP/J+EBno6tq0r2XHgBSSAxeRMycZAe2hC4Y2mEzxMBfBC29Dj1ujb3RxW463p+
6HaaIHWso8o+R2KZpqHRmRti/VrGmO1C/8PkcyrOEsGYgR1CBOjqcMSS/aLS3g6j
SD4MC7MgGqX/jwwd6hcbf+A7oCXm0AcnwNzEjHwC3j7DfaU9ndelRhf1Y0AvRTBv
tvdG2eXqlWKa+59j5P4tMmiZeG9EugSb09nUNAvH+lQ5LU2jmh0vqWsJI2HBaZVb
NS4t9Skv1pZwrI3tIxGINT97KB5/L4TpLJrAqbfIMvANEg8SdFO5SW4fn3u0Xm6x
gXdtSenfaJO7UP6FgxUayOfSkt3SXYx44Lt6UjLe8YdqDzZE6M/wCDxa+vjoItKH
YAk2AdCy+61rEup9g++1ORNNlMf9YocXGngu+JheW/wixUik2cWFncG2xz6SZGml
rhSo1AC20805C7Pl0JGKTvNmeQREJG7LbQsxbQ+/sVzfKuockrCOJre7I/vhb0f3
EXDcVmNC/7fBroaMHmSs7y/gYVderOeGKrd4INiSuBm50pB7Yw2iYZGNnjYvqw+B
5Lgu55JnQCOdVQiXJ7x9Wo9Nwgv5aWNt5KfgLdIv+fYR7DNTW+uvaKPxODrSaQna
zYoWvlV/KP7+RdMoOtbsuylHoec/HqtmRXv5lGuZOCMqU8u88ai1vOE7YT3kLPD9
54lHT2kS47l/xdTIpIKuPgviFJ98xUBI5JpIVo4uUDtB7zw+ByWQGntZWF87otPr
sunsoIgh9Ht4Kv0EHwVMv5WM9A9OkR7UN3fs/VQI/ppXXIKYrTrR1hYL5XbrYsBp
0+3rjtxaORWft3j5fKlWHd8geG3vnD9Tl/Ux9NsPic6IDkrschbyKfNNmhXYKnnB
F7nIhmndVrWXJIh/t2wUHSOTm1M79kRrqJPwO44O6Lgw9fyEJDc5bejknFg2ne9b
CmbcqaEGNkmjY7Q9YUFEUL2WNBgWJcSKqLHITJHI59fWEn+q+DUIOgohC5bCtu3D
gdyq66tgU+J3RjgAyJIPnYKL/zzH0gQiEhtaa3xZMG1PFXuxIB/wAjkkGc1SUsLA
04R6NCDxpynTEKRbPt7AHkIz4XbWa7jl4usybNdxd1ZEPCW8ve1szyNFnsGQfq6g
VzSLqEdB87yFXMIfaRm9DUzdhxOOb50gNlDjqs3HY4hx6cLQeGYz4joUT0JvCobs
OkIR5NY4lGOasqPC6vGnREJJG8QhWG5DfJxqCuVDF/MkGngn3yEo0/hLizJq/5ik
4d5ROUvbuSjothr2QENgON72R4BQHyAicej6cE1i8siNku1jLGOPLBfI2d1nOYdA
3R6Kstt3bIyNekwTv0KXbayGuFMVCSSVIUaK6p+AZrE=
`protect END_PROTECTED
