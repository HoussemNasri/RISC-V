`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8i/Zy8soO9HA0pdIJ20LE01zbRDa9gNcbxE68NB06xrabYSFwfJrb9MkKWnam4I0
UzD2cAXImu2Go6FxwjWKdnxnGIz+yQghfqjXn2UTneEGm2DxZeXE+n3HtlEX0zKU
RVyYtL8h4nj+WoiwiQpDGdaVqMwZmUPia9hyvZelhRCkH7U9sRs3Nvyff/pkRx3I
yF/E+bv608C12LS7ZHi5JA==
`protect END_PROTECTED
