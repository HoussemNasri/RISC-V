`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HM/kxt+ZlsyhMOyARHTd8uLpylMmgLihrwrSr6I0SoJg1RFls2/EfTKrmebK+SwO
MRhlmj+lOVR5ddjLb0MQRdQYqtARr4WZNhucmHT93VsJGA9t2crlFXzx1Xcd8+N9
JMHPNlJhXxV2yTLmvKqMmDuha/Y+WYal61LyJXqw/U7xSBVlNFHOWDJQ4axdzkaG
k2E0AHDe9nu7XroZjsw18ma9/K7y1gKfwi0W9WhnkG/SKlOd8/tcv7663mSpap0a
4a8zUDZ9fWg/JkKfIlE+IEjv9UztRZ8WyOXEHetG292gsO/eLwb2QxCxMqIu+sNk
X6ZX0IBhWU+kLVAHuog7F+pB9b24hmh6ZaxOHaata1LMC+monb2hFk5rW4XhjTy2
gj/G7mCV5YLB9azBkIGA5y8iufyxubvEweiD6ANzIuVBTII4I6Ye8w/XxQD5civd
vEMWmEOCA6ZYCbaw8EDRJinIPwBw9PV5g1tFYOmsUZByBBYsm0W6rBXAeRts3Aq6
M8NhHQJPJHK6z4qCjZAAlVVDZkhDIP3uCcahWBMWQJ4eLBdJwrdz2C6+UMW/5iop
/g413B9isS3PxD8J+zT6VqXBBK7unK4ycAOgeZQoSl0hmsvfAEhyR+qycVkUHBi1
hMfFxRSivfbG1Lm0GZ4rfZDfYr8lfnZKrF/CFOCPEM6QFkkl9YsAdPKCGD7kFPfQ
MSgg0ie/9vkrcG5XeDyfs52sc2ZeluFnfXLDmI0m6om5o7qNo+Hq3NGQxiCPCILw
dDNYtWc590RQ4opLmFmSymAxbekPhH6Bq9+GW/VT4++7eueCW0mSwPVzPO4eLVM+
MZ2lNwKLEBJmKrZGCXz8FYEN0rGZ00h9cv1A4Nu3/cn50mlxTGu19Vy43lKbHy2q
pTqXdl5x7Ni6fjqHgk5J7fqgOIFpKpQTeREac1pjHaklJHwIn8k/qNtRmsfwoE4R
oikttd77tHJhww+uQWrBX0cyH+FSnJtLj07r4bsT40Wp7NIm4ae5iRbQuLDykbTD
Vu9aK7Vh40RHCNXt/FB6UAlShmjs0S16UgA9PmBXnQZzarrDTvA96MMjnu7jM6fM
v2L+D3HOCaIKOVPUcBoJcKrzfMoZOZ6Ho+6jQINagw+ktU3wvgjPyR9XxxETofUR
XfoBTlFQTwN97JxnfghyppyrCaf1Bmj4NRjn0koFpTQmXIMokaQVHt78ssRYpybx
oMjIIxQGLeHZgz0/M8KAnKexC37Sq2w1TW1roHO2IgV7pFkpzgmjPt9ifd1U/0wT
Fl9dZ6Tz16kqMoy9vcS3KY7OlScOW8LQRakn4iaHcGtT6T8n7d3cTwOJWFxUT/4s
S4FSLlwsFp8UzFtZEvlm/ctFzDj9GiYQaB+vsfy6q/BBfsUVBaVH21Y0AtP99k/g
BPEMNd5IwrXa10OiO8HNiYobRryRlJBX/PplkM2Gp5dJj9hwvKZWj24u2mfauMl9
NcxrMxqCXa4GzTxDTVtHK4+779MJHSDw5R7SKx44hyfEDbjfmaWVbgO9lFaRkbt3
F3NEYQ05jGikWN9dDmZSXK0mJOATcNojoedKw+VzIJDkWI0cFad78CX3OPjdKXHk
MawVd0O7lKfIEc3s/zLaYEUh0sBKwOdB718kUskhCpDitrUAifJpVcEOzPMLAYQk
REMR/SeIp074F8AGBYpygzeLYx45yqDfRFDMht5gnR6dbNSLVSXCDHq1m4eVvEHh
pMTG/lF2+GtMdrx9PIag9CmyfirBxCErj6DF+opzAjFzm6NiKXtSpJeXVZtmUZlS
KY5Ny8cY+Uq6RTD2dzrRtInudK3CcGf/o3s8emTxM/MCC7rtttRSQGxG5QCZ/w7F
Ib9w2HnQyM5nYnk6HVDF6YplE62rEzRMBXyueC2GYO6T+oSsVPgS/RSAGdTjUOu6
8jG6Z/7CIeV587Axmb/226VQ498ciGQVJBA/jEFC/oX70tUee2RAdozbuGfLszgw
vipUWnt3x/XW6gLv8+Fcs81aRwGqk5IYibPMrN/1Q9xngHxj1Y4at6zx5tAFEDbA
7kjDBVDM47DkeVXFPyceAykjn3AH+hfCCNjrWSLEVPfZQsQdsVt5kUzOycgGBVGd
oogo2LmeMrr1tm9g9a4gUuO7DYQT1V0o/PQWzUClYcu95WOKVXzId6nLjkZ2P28L
YqZpb3PIWPgB9NfS6cGWqSw2eYSV/L+lKv0u7P/BYNVKCu52uMQwEa48bsoVNZms
E1cyK7F/DteEDaJU79O71GTzxI+a0ZCAWMdEPvcCnQDMUBApK5gjBhWdCAoGIW8u
A/ZqtjQzxHL7LZ4YKCk9CJpUYRCFhnzr22aZM8AbJrSimXbqKIDrdUB2Eo3Kezrm
OCxZEIdQIHBCWf+kD0x58qXLNVkXWUFtSpL+ZjK3mh4D0lBlMWuGnN80S/fTuD7H
qyzqjwGgZ8hklJV1VEO04J9/0cL+HePkUHofPq7xFY6CWKK4AOeYotcvW5qVqgYJ
VsqhToIyY815NaoDP69jnJEJtWQGpR7AjOOh4SjFqLPOEnuFHcm+MNWa0xvZIJJK
VIBeFAMW6jAM5LTdflV4Nbe94Byl1QfrMfiToB2xfe9itmeeJe7rDBGlDddHfjpQ
0C/8FXe44XoT3ldy3Q1Y6L7K7tVXCHp2Rx4sOWXDWsu0lcLEgXYWjqrG6a6ffZzW
eb7PrsIhWtoUGScnKsttpqShp6Fvw9LRYyWnwmIuUm8uwL7WO7Tdsy7TsX5UPEkl
f/bPfobMdphzEVh6Rfa+DeQRTp93TZ7fjBj63O7x5L0XPqdutk3TpehM1VXbL6fY
tTIzPccugH0m6mhFys7hsfnRv60u5WQOv1pjHITUO8zYxej09yEpSBKC2tdaUnoR
PjZHWH8Z8bP8GRDwxSp06zuI0uyaSwJMXwB29AQ583WjBs0kLHwGpCc9uRZUKQau
+W9F0ae8dzp8rfhi+NvdAwHeF5TEMyrt2o/I1bj4H0WcTcTj9y5Vzx+evZdUHgN0
vCLGYT3ph1ucuAZHFb6Uwn/ZGj5p+ETp2c+syv/ttxYu8dhwfW8dSJ8TAfn7Z9Om
yxnzbfwaF3VRXnuLPut0vbIy5cRHdZxKFq/f8IssO2wP/oCaUYvBUUgp5pLzxFwe
y5S5qXzguZbNBhHKIlolpYqyAHOY3WQoGJAu+ghGRoVt3NQtQLmpRxGWHfvuEr9Q
km+QP/Ii6Q0nlj8ZVo6JJZ1/h2qKLgi1qk1vtMFiEa8xxEdj2TNypeDUr7IAJflz
zK8NZTVzZWlJG6ijA/dA9Yx8bxYoTS5Suxu9PUkAZrxzNXeiS84ftyaa1Ui3vT9W
u3Mr4k0UW5XrBjN95bH5FSK0/b2qh+Gz3IJlPRAcMp0Q283/niTih4cVxu1m5874
k4vINp/HLY1hvzt+6bRuI5q0xXAvoL6NHQbJatnrypHH1zdxtZMcz9oHdG8mfRBL
o3av2xP8fb4s0iGGGfu+BEsox/DG/iup34COfwxObmmLiHSEwjUhVLUWprfNm7EQ
dQC+fpyit80+RYgJ6OWnDw2SAGZ1AGTITICBII12u0KMDQtWITJHR8+k1CL8FzaD
bd3yTv1/itOt5AmskFIWmaJpyB2s/CyVOSdZ5aCl3J+Wzp40BbTTEuOmELiX2Upy
I+0Om+KNQl5kt2uJ2MJRTiFRa50NV7ct4f+L4/IhC7EIgf/MELWc4BTxBmzIJCrE
o/C8yfVfR3llTwRghtLIrytANDoi4gVeQvrAKmmhraJHzA5GEMWSSdBMASpgUvDe
ENM/G29TtwlbY1YVRghGGCGMS6zj2kzes9r8Pze+s+W6AP3De+TNuiSqg/zMtlgq
lDwBaCtDFAMOybcNLld254X+E+tPRXuzN0dOoTU0R/ZauyqBFPxsAvYTVncaaB+S
oMgKAfVUFdsqNUTRngCF6pRCNikHSc1OkHTow+wRInYDD+i16XduozrKAjRCn7ZQ
6ngP7uGgigrcrbD0qN2BbdH0VbM2U5rls82v4s+ZQ7t8gRmSFeLh3b3dejeqXknB
TRpWp1p2dAIu8Atp9CxB4HEGVyxYeGH3aQGwjpRjuACYrFfrLbZwcNtFWzM+Rusd
v0UFqC9jX8bvkSM8vY0wjUhmifTV28/LbWCC82ljYbOmQmrDqGMXha4zgKrecA7U
YG6YDyOJ0iIgw/+CBf3pylYzEoQxvhukuswscdA8mtLdBqDSBCNr4hTF8iVGfqJf
/y4n7pnCgGYSz89j59anqbwt+sc1J9Utaf2tkN4C1UMwM/Xiygj8LLbvsxXsG3ls
VFpDtX27tNuq6QjdqDu6VPBG+PRAGts1HFbKmKBGGRhX7uQYXT7R6LsVSQgFPKNW
0M5dgunntGKmC3/Sk8gU+5uZjhfuiBai6qjeEZ9joXXNUNTywNc3uSsK0uPxATch
P8na9sQSeak0SZmzR8O08dW7Fa5w0GpO90n7RcDtXTSbTir2mFfakQSg1Aivek62
s29eiWc4U1vfge8RSyF5sDBpAjZMMVeYheHnU7plXKPZ3K0QaTMbzhs1+SvjhEO+
KnatN6rWGLoP5vHUWc2R9WFs+9vnQF7UqQVoix1TtcRDlv81L6WmOKuXobyx7Wn5
17wl434OwJb4WnZbZlui92UU/ggBYMiBqbPjC6bW3drGVyfSXLJ0isL1zi4ayWlf
Mm+GcamuT/KifNjDsRkOEraHASq1xl+clJb1rr5jasrUy8pwNQ0n29DVnUVqtCFU
9Z+AkTc5hRgWrdG/ZguAJY9TTWnOGSTkaGl1S9GC7uddVj8N9YMGPZ47MIBKlr/U
0DHkrhngN6Ksn78SsI/Ivo1SE1iJxl70M6vxW2uXt9A43D3ci6QyfRcS4bu7Ktxz
V+HMgklfqRLjSIe5ubPrLD6wUK+ffoWUOfYpNBRx61nsBuTX8rDr0lgLgNhY8JQh
2Ecm79f4bQ7X5LpUn91EUEr7e75sFdHlrHQbjAebOiDQ81UyDliDAwodRLTA+2RG
XOQqIYSY+k6zCRK7bYSPL8YdOwjjxh66NK/QJZQ7XZwHV2kEZJH5DbdUsrsE475E
q8c1+X5fbXE5W1dHdrrYTV/CBcsPejwsW6bHZoOpq7SRep/gBhWXe9ubdIknQzA+
Xlys2p1uALDkj2NWpfDPrUwJVpK6/jmsqExsfZ9cjc70Kl2uPo+CYlDZIToUdJ1S
0EaIipUqIiw3zmqOX4DYEmrNkt0h8//xR7OPcftYWpIze7V+vnLjNr5z6lQ5QoDX
vGYsUkuOpJnfikk0NGkcfweCs8T8hMICCLM9rZF1IMzQuK6MtqRW8kjrMVhd7rQ9
vVyLt01iOoITZIGzTAVH2WakzZ8ZiGFSDzjAol02e5KjtxsEp36kqq7aI1m1P2io
nw1Vwyqqm7eVUILfPCzDaUEsC2uTTcUEEUJVRb/WSRfdOEgNU4+wUxBWd4XmQZ12
TwPDiGcwfRh8FSltoqssj/Yh6dEHeRAadyKFxYzFqYkFGepx+YUYYxvePqUrbOdu
T5xjFxbbfrgTw5KjtD3+samDAjXvpuv/mX4LcnEGmyeEim26WX7torSMf2Jm0LoJ
iMhQpeafgvffdKtN/xauSzxch1iov6Awr2zAKCCFCOii9MLz25Ecl9gnaSldTU3b
vsC5G1Ge45KLcmV0cmT2kmuLYFyDN+kAa8LzzFAZ7sTODoGx8wPexzgAteb90NzQ
DJeKn/OIimuPmT/d4bnDk526Fi9P8i7t1FU0dnpb1AMpsPkubEPKG9zHZHqKhRGa
7LD+zsWKpa34+OKjpGO6rv18X8ml4p9l8FKD7/l0mVdD4mE+o16OqAW2DqrfY9R4
wRd0Zst4LpedbfxF6/E/BkkPzWRZEVCtHC1Tg7HUDGV2Shej6WRsfCkJT/s/MPAH
D9hh/AR6iFBzCHv60M8B7Y8LGVs+7LrNZJeRwvMrA6UURCm/dyqUVihy4rrZxaGR
wyU+tvIUEJCmRKu8zluVSDYo2W3mtmG1ojMvP02yEvXumPvHvbk3qy2M6RRQumgH
Vh/1h+dZqTxMWdQFhuopNCnf5WNWgNcyrFrRB5AOKFphz8diGaBoKYd7ekMnhDwx
qMKcVP6kLV8mr7064FjadWn7SdghwLL85rJCEc4WzeVxOREdJRdGq8s3We4DNbAP
ZFSocqkOww5IhdOGPcMsVnMkxGvJnJjeasfDaUA/gg9+qnc4ainp62CY90gN+fSo
Mtd58YjPVwIfSMN1a5Q6ZXFqxX3thL1ShSNzsTnhPtWuiwM4/oDq6qRQAj220iJe
s/AoQqpXV1iEn+H/g+2lmdoXmKMo/cE/xQfLZkZ/IVHyPX2hmTo2hHhiDaqhi8Yr
TjKHFy05RyhyFiRgJH+sDF218MdkI+nGpfgqtjqlCE4xFc+VZR9MhaWI3xCkUdfq
lWp8DiQnIwld4/PkXqUX0k0RJW8HXTTqZirMM/OUxzmXWpSZ5ibyxN4ps7R7++81
k7K7keVlgNtNiWbxlTZbfpod4pyHGNeBY6bGtgbUViUcJsZUnitvuGRkDI6yNctF
pjTzeA+IsRgFmHkmynZIu5t4FQhecvftRgVGd3++/+Cm77vgDR9op3xdFWdSxDYX
9JuhzJTmo9pUgXC52BABnbWFLqdhlWndTzp5ZuRsrzIJrDJk8XgNr9RWPZMnSwDQ
N9O14ra9FWkz8onABCW9wzEkrrYI825ieLKfrFN3FPDyytEgulr1En0Hg20HZSyn
X4CztlDa8bwVO5PtkMcvWSGobKUs6I7PTUQ/e2uPRm1rZabMpKE0cHzCLpjfm47S
C7c0cfvv5gLieZCfdbqbWktvtTmD+GDn3bOm26K0GD5iPpmEJHpZljadQ1zNpql3
3YI29GrGwW6Cyn8AR6kddnXIunPTQwxFlbHTHtXRM2sO2B9a02L+iM0cz6psh4wg
dvKogfDygEsOBIZS8E+u4JwN90zdsJSE3ome4aOJRAVshJ74cLGgOTDUAhJwfpVk
d5KbZcM5CBqe/BsmvmC1pG362cBGz+OBg4RluF/nSJLemtQUuY+ZarFNEvbhDDDp
xb3/4bPpBv/KmXk7phOSkmx+KDTtOcGzvkd3FOUc170C7sjMS0RhqF6ITUlTS1lu
aSINo2aK9ZM5+Hwwgx6Ejbre9mtHT7FJ83Tv18kpJOq7a7HUEM+qKc5K61M+qFY8
B5X3/eOXVegpyqTanCtiC4Tiqkoieh6Jq+QamkyBLYD/6ztNdmLvoHUXg7Rum7t0
UPk73/7D2HBJh3XZ24N80+OvZOKWXBn9yxEKFNno3ZUYOt3kXOEUltyFPyL3Qnjd
JFTjsdGULuKBun6PDtoG86LEnJk28FGgNuPuK2kiGpqg3/uasfD+cS2RF1LIMO9Z
Xrz5dXjBR7Qq2H69cCaQEafXxVRYS6SUWmsFyFJDpM0hQpihErxOlXp1Efb/toYL
VYofbSkkQjih7S8/A+5zw4Xba3XNrkG+LjtPMngqM+K0HpzgZF2LL/ZGmerrh4Nq
9SkXT1h9h9H4L6V/d1GL/7jF7EcR5/TQruCdaNBJ6sMBy7y/JTM7Mqo1cTgO5JKb
qj6ohKOt++ZJF432fldK2gjBU8sbvA9hbdEHuuC35c5p+DyvAn1MREOocF8yNWtl
QMItKU8/71beBn33P2uDF0Ao2CxddfrmjRNxNm6KBljMCuyrm7NiTHT3xoqR1YXm
K85YCtW7xJ80bxKTzR6ZCEo1SS7WaDP9aZFMcRPtHleY7E06m0NKqIjxNqHwXQ6g
fKzXE2fNqTuMcOgBSHFz5iCUPPSwSj1sJGwvxyE6FnbvOfsJSZXrcfIq5gwLABNn
mKfTmdty0Kqul+uZsbrqfI4HuDcUU5dzvUq02nDqJeFohaKpXq0+/sYOVz+uZvsq
9OnSKTTXgUSbRae38RXXwJDtvg6doqPsgeWYLI+UdslgWXPWsjoNTZ9tqvpbir5b
b+jeckd2Y4hm4HR5tHExjqgyFtYLODbpbGfh3gOJIn4qrrlMz+exndEnPbY8oH9n
4wRDjw3GwNcXNBAS8mhJT/1HEJpvqm55eSn847sty4gpvr7XXSxZF8q/aLkZNKuJ
oKTfsXZzWl/ZXuDwI9PL3RL1DuqBgrneVvlPWgQqpbS7JvZI70sIbycbLKF6/keb
v2TAXd1Buf5ElMyXOGftpeK0h3vDeV/SV58d44ytqCMgP42+kX5U9iH4TRC10ZD2
I5U7VPn6WtnBkqI6gUYDsfouRyatbOKBwdJJwwwcG6L84EhioeyTeOkHDjRiNKpv
tpxQzHV2Qd/xDIXVv1hZFi77IykmcZNzEcJDJQBl6WeWXevWj8g1qXjXd/qFe6hh
3cKD3dD258m2VhSsXBnwckQvCLhDu5OLdL0u13flDioEIFWVgkWgsv/PLsC6RKMy
nCcmbv0lmjvIbdNouJw4Kn80d6JhGNYs51KHvvDTBEMVjvaJmaoVrt57OpSFhot8
QdLfw5UDOq0QSeuArAtvRSf0QjRzpuSCMb2LIr6hQk/O6PC4Xj9crQAv34GNsy1B
r9YUHPbP38dh6Ml0qDcoNSOEG/RsHD4aMNysyP/5l5GjCi8neS6nDM98Eiqx7J4O
5tKnlJVfQu8/DkBw1Z/mbnDR66COQOkuJo38kbjkpVWNq2r5N2UFSX4NzXY1rhso
DSI9KaB9ZrYo69ORuHwPD7BrQ2+tvDlUEO/KxDDfRBer39GlaR1CcJr6egvwrij7
4mnvoFwEuxhT45Dg3Nayt+MiLzpJCur25Me5ZFmKyTq2FD6N3yr6WAo1Hy0P8ftm
EfAbvcix1/PO7D1jqfxlob2Y3+FXInm2J5q2n8es4sTQJuPh6NxXut4z3aFXRd2Z
d7/+2psBrJpUAyipDgRzTqDjkkTEDuQmHaetDmJjw+af4R3ZK9mrG5ig0+ZETQqZ
VGUFLblpiUNmHDptLBPzosbOuTCXVTCHQlWBldYiuFHTC3ZTaIxOs3HcT7acfWhs
lw0pAe5NgHuAnHXpCXEB9t05bgfg35ZkHU+8Uyqs/ceD8hyDMtJILBoyCBFPXp3u
yD11Ysw/rIZvOjae69D/aUKiOoQQnzJtL1YgLZHA3TXiIF8TpG65Kq6Dsg8kuUfK
cGDfMyjvhC3bwFFox2uacSiYa/BxgqGQn3DYajy0LW9geoMZ5Y4mc9n6yCY+VfS9
QbqmizAl//W+tm1ZBlpgndDfAoZ/sxoiLcWUTg3VNxdA/ZYXxQKkSlA0kxATYeDV
LIgac3cC0ERDEhc/OBe49wWI38SFdt5W3y7DLJQkbMosMZzjHH99lINF1s9/vUmc
Rijhyln2847EFI0zMCu2dtVVkaZ8yzaeXzRNRIeeG6pUJ1E/OGcR6667kaXTWOdm
YKr8JmlrkkigMCwfuxdP1CxGiBuZz1rFK9sNsjmz7LI9WwCT5OH8CVTy6MVNpplR
kfRdId3NrFw6cE1E5zPe2pMepSNo3/Vgc2FSHLJRw9HWKEHawZKx9IhKdBb0M5Sr
qNn0QhjMzc2kG3d3Qp38e7MSWaYJPb2Jx1MWqgSSPQYjEzSU6D/3V70WifBK/iBr
qdl7d+9+tQtZPFxj8a735wZR9I2FvaNKDjPykGrX+eznp71hYt5vLt1WKDhi00T1
cnL1lKb5D9Es24t72gvtTlcGvSqrdUhi1Rz36dmsJbwDFHYtvv3SAk3zz+CajmJn
JOCMZdWR5H0fpOrhl6DFfQLKx/2WR2bWpNU5AUygJuYOqQ1Yfrh9ag24VnnEI+Cd
gQeFnTheYcoCcE+M7LKW/FjsUOCnC4FxyZ3i/qmImb8C+LfxDemx+dmXzt5SmGEJ
qavv6Avf7Vdr0tzAng98INcMAGUmT8Vn1cgSRNphIBkwYFpGFdzMPeJ7XVhhuwPm
IYnSXPDaeA3R+OzqLSJFMigwKT0EC5dTvmrLfylBnv1eYRgVKvemm7RGsRC5cP+T
RfwqnRa4FdO2LdpMxfaPtYjqO0wh/YmT9jQwhGNrozCqr3BoYSn0THZmLO/uA/vj
g2qbUuFCVw7Ym2fsahV4pUlHtwfYcnx92uubZ64Bq3hAR4FiHX9QYSWEXB05C/Kc
q33OnBknWhvEUlYm3q7YZE1oPWfC4qdJbMyMRMJYz3vHJ7bvvyJvsCcX5Pm4nAyR
NXgRyMnzzVfZgLYLpVvYYSM8fLTkjZ37THoip8oiiuxk1Ft0kr4y5jIBqc6Sd48A
LD6DggrmTVqnxl98LjSFPbikypx7Dw5rkYeZUHbxR/VTriXXFC26+aOzE2lhnsah
J3yVnvPb7KJlhcWB2UCMUfDBUSUBLUcfavPhhm5c246l/0BY590NS+xAd34a8TGP
vlBPtR5hpqr3vjz58YYYRTb2dqjYMFJgY3MBpcoEGYKHes4gQCkMZzrCZstrO/vZ
Gty6xXQboDwHySZ2JUUdaHvVVbd+VxVt1Zg2QMvKGPXttZjjlsNJG5kmoZMUpfHX
5uFFvx0USdPJIfG8th5BkPEMcjyvqrrd2Zeh2WuPbOMWyWD4YSabzyR2EoCFlyZV
uXVdlSxyPYvnjBxrP+SKcVpuJ8BYp6DjCGF4UZpYWFYWaCa/Qz5AkG8QneHZJWcq
lOV9p8GpORfQlMyzVljGzUPPg5duanTp5yXzoPMZC7Ode670mSMG+/5Z34+dyN/e
uZ3oWIbI930af3zQvCISBQGi3k19Rh90wFBexxezALOgFKfk7UYsOK5trz8ElQZK
OoxanXJRiWGRJH26RXJxe/EUP1xKvycLj9740+KO8XSpJl/I61SN8GXjJVRYSqCf
BnE4MUnEZIOoCwqICGWuAXGBfll9yoKQwgf2a9sYQdu4mM6rTKopkkuVaiCOC42p
UP3nnfFzxFFcIgSWWHaFsmqTWuIGmDjM8kgF40B8cm0CbvizGefiidDYlFO07+r+
adAGgmlmFysW/snGH1gt8SwDE5uId4nOrINVPeqxJwG/cgBTTSpGI+Ca44yYHZKT
6wqh4x49cYeqKgf3KcUAOHjMMrKbxjH9X7F4gutS1aZfEMqEL3HtyZy6Qz5w7izF
VHNl1jInSERkX8KfSgIBiAfrtm1+7WXcuEPMku2yewrKEYocmCTBfpCeJhoiywVz
ohKDL5GeovdL9GqAmXLVlNJXTIZc/6CODmjg+ZMg14ZJxnliRiKFxll8PH8KCDkL
ThwgabJ1GZwCRI+SJo0rT/2BHy45auWaQWrNq1NpwRJSkV9ucRAmlyzK7npvEZID
bchh7zFVNVhclvZsj+uwjn0crSwz+/M7GEr4myY1HvxhmQCfXmKDiqs5G/TIDOeO
7RznoH00noNDoyZb7WahfxbBLG13yUymYhCb3p5A0Hp60rs3ARFuS8iRlZ2gJPoU
0ynYfNBLPkO/pp/iKqk+LRGbPk0DKiFTblcFNoGKu4P6EHBNkBDPJYA7UjIqPzFZ
fzoYnVN9NXzLVzeVgQZOWEzwJYJUtJkrA7KAmc2afjWckHxBXZlxwcXuZgforjoU
W1pj5pmV30hbswgmiITfw38/vwbq4ASaaqubhJC2vfb8/7v8xvVGYI26xiJfLa6e
zlnsKuu93kAWIK+m1jAkTBUiV6otgLN/CtRdgYjsfyt59dD/ApJwEJQ8t/S9t/ux
PpHzINUNOzNg/lcR4cJ8c7M0tUCXth4Oqm8xcs0nP3wlFPDxKFsDJAaTzc0wQkwd
+0SS/VMZpDc8i+n/N4ggvpS4U4RRxhaOZsxxOvJpIVvkCfe7wQGFnIYhJ9DRq3pj
fDBQGpsfepd+cowDhwpcEStRFsp+0zLRJI04ZnvVSNyezpI+w28h89GlHOn2Q8la
tnRXjaUOE7rx8GSz2hSmiXAo034Mro7qQQrQGBYmT1Gval6URGR5WYLcwjwvvDIX
WPm2/BWYtYRPGUWLwSoMiARwxxT8uHzHxlGzpgYw0Uf7RUKHbbg7ltI8iVX+J6fr
9yz+mAHtKb3TXeVcZ23YRcu7YMaKRyy1CzImvE/E8jOE8vaaUV/zn+oHUTsS5bv1
V7qNetOI9TptDwDbKqmVtP+zrwVm+3dGsowFIKbfszJERedEb4/U6J9dgGN5j++p
YxOgLPjaWtu+cZhCMXmhCdmOYElnCWeeFQ80AQw0nislZ9whAE+Q5XnfvCwfrBbz
6OhhyqsFko9b2CYgthkVzmV6iQGa/WPxU5bmE8K6ReKnlBKnGPPgZdyvcRhA5PDe
7IJ4LnIW7ynBj0V3x0H/vstq9A6XeLPP815oupDCAuKzNCRCF3Y0k4JtWih5DHIz
+MiI+yNFvtJQFZ7NqLQMTYEhApBdEAxJ3yPaz0yIjzOndA7TgwEHVYsa6N451Gic
F02xAmJpdt7Qu+87dF8SgZ3dxIAEygSBrihJRZsIU+zQ4o9LXSJ0TDKNIaCn/PM4
gMq7vG1Ecq/vsF0/u0CiOcdjCTRNpVoUMVBZikO492pOKrtHzXXCis4MjZXNtPMa
CAUJMnJ2avWLpjjqOjIqHp1cgCb6c0xK7z5XC1LVruZMSiOgKS0Jw3m4N8yFj6Q6
4PZYL8WzJEzIGyYITLTviWFip3vl3zTrknoD0CqqbQs=
`protect END_PROTECTED
