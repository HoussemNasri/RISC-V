`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEwPkyOZZn7HDlUxDTP0L4KNo54MAsSiprb2t/gyf1BbUUTXLfD/x9+fZQkkVNrc
nIVFTZnftIRuefkFvNNa8q3FRJKIbfw/+EoTyN2WVwXzFT5yydajXSgp4egPeDDm
YEjFo8v0LYDaLyjVRRYe1vKKeVYATXYvM5phuNvzlitiaz6zC4C+6Ogd+qhnshEb
jkvnejRH6DGBsc1YKlWKWQNiu1TmTPfbhHdMUCJZEdkSLsBIXlO59VRlL/TzhjbM
iLkjTFacthOADrvwQ8Hz0MToVDV7uhCs7ukE94xoVjoMmYp9WxQZaPzyXZycHAQq
bO8MhMRMM5ShVx1QgDMXwPgd9G0bDG7VQFE/4OVuoiKt5a0PyH+hJGEIhdu+BL3j
kCJEQ0CS/kb1WAg7BdP2ikkyK/loZ+H21TKqjJuknvSg+UOE+6dzvebkPwOdVsMY
p5kG2wckfsF9cGKhWN6ALkXsf7dfaflCUPNpLeKzPLOEJVWLz8g6oQ8lphZ4nu/T
HUnCr0XbNgWQn+YzVa3iHTAo1Mgnogplz6fr9Vubu0MF7upbsibQ5tDb9e2BJWAD
3RztEY4t4QFO8qmKaFyvAqqGAE5Cii36t4hrV/pGOAlEqAz/j2QFQxWlDLPZrcHK
tSfg7sz19lDmOwLiChuwHiDoWqMlEcrsQuYF0Ud2aBOKruvMjpzfJFISUyRS+fOp
RihjRiZndw5FEDgzaYmQBY/u1UBYzqWZjaNw6B6ZH2i2LNYX/70rXYJGRzs18axc
SZhq6Jekzzyht8BKk+rPTwXeh0qsTy7uUCQCNAXV381q3XRmtmu2/QN6UgLZHj3K
usGg/1ANc/7zEM7a1lUjQj+UeBvVwjqn/0JitYTsqgkGphCiKEEVuOkYEjVIiCO7
dfzO1pAiMPMQECei6/6UwFP/6wxwxn0ZhC6oNxjlPqrtCjE3rdgV7eneKxewVAHu
h+T/gm5CyZAF5Dyby7bekDLQHbrHUNQekaXUqARTRIEpu9EZQ+alV/SaLDdcXIve
ymcffdFe5LclANg5PqocKsz7XoyO+8UokzeHs+SrxQcXYpiU/5HOwcdlHRtGixzs
PVcxlqdIfO5xfausC5+OOyl71cJFNNJyOkM9yQ2Uc6ZwghXJCb1lDSXlWIMyJdlG
ep8wYkieRkSebMfA1VXaxeRZ1RxlENPys4QSLZBRxJj2raUI59s8xSt3Valmuvni
pgxZ6Sy11l82Z/lPP9nVmvR6tEUTQ4hutq8rGguShdtITyA+oD0/PADa1RL1DgKM
2JVH2FcPIpD2E1aH0pDOlMZPYOGz72bKIMIQcNwZuCUgegy553ieCjBOmACREXhZ
4Y+rV1+Z3qjybJU4Uz6eyVv9W9eNO03LPHTIoEoRoHxe6R3UkNrSNt5s2mmN31QM
uU/9n6a0nvrkdAwUe7dObQ0yg0d+UwSL0iepgB27BsGJ5fhB6qxn/IJyXRv8IMjs
aFhacm37CZkQsMeyk7ocz9JldeyeRxc9seygACojAO3SSrk2H/9+cViX2DPcmY7A
6VhMc1pb4SwJoYxbgbDa27IZdg1wvdhLPwsu7vkGq66RzjC1/S6ivSX789P+ZrRr
86UfvRupOGn+lBee9i54WDDKvebtzSGLw+dehd4vO+tTbpLOCmyq7pPErkHaYTSu
WvF5u9dA3wYQbiIwG/LWOX1QNYHEGeAJ3sV/JHVvZvPbZkV8j3vYGXWAR1/Mod6x
eL69TWe2hPPIVYykm4s/6P+7qGNQo4KytxPEEVRN+UMlARD5/iEKv2w5LhBZxgZe
UoWkVml3iiWODcB+oAJq8hlR06ba1T7zj+Bdj+zWGumCQYTTkvuoWiZ9YZk1qXF0
huSvRlfbBWcCmcxznILIeCKGGX6z5SP1chvBUtu7rTW02d+iflsd8A3XFmR6ran8
zHj56PpPDdOWKdfqPbpxjauZyuFAUlZB+P0vUos1TAmQ53/aqxwzLQnqYUhAY5ES
J2GzRby+pUT36cqmkLomNvB7xIzEX0zWm+8h0KtirQyZSY1yL2cKOsuhY2mVZy3M
/NXS2JcpsEY5UeYxBHL6CA3AhO1Pb3WPC6XEgJRZZ1s53cEaOxDc03+x0kRFzlWx
fXToKUKZCgF0JGZrtxcjcuLlttWc8JFheZtvNTjl2NCp2M9uqIHqJ/Tf+2T1Y8pm
43gAfELZStn7Xkb2736sY21AlFaVpxlNiAVYt1JibJKuEIMcD7vcwxGTkLYB0ZxL
Pkea3l8/4QbI+gxZmrPSuiNd+nGxxEF1hj/UUWsjTd0tE+x+8IeEBRvYSKNxYSOf
4EbfFgVz41E8J0673dNfFtGF03xsUexPqI7bk+Lmh4E5tuIi+iYKd+CaipFHxwuK
UX3Mtnwkm4mc4oIUFzPwCUoCIi6icvzWvV7d9DuB+zLd++HKEGAsqS2V4VVymwC+
vk7nSO6UbN1Pvveyvd4ID+xBG3QEpwapA5x+XOIZa6sQjepWzMUs0iHa89ZdJE61
gBba7yJZWHBUnXXKCc8sm/CHDwtopFecOPBLaLTTa37NoElX25DlmPZuFIajyu/l
Mi4fU+8Y3OM7Su3LVvUUNY6bszYyLlTQ9PgCSfvyCmm6+zl0+1oHCi1xriK7AI+u
q0Kn2z7Nh5j/vOHpcndQcCX8XebtI5khUf0mCS6gvdAqZs1Ew22ffASYvpz9nK1x
IJT5TJ/NgHT8Cg5bJ+beUf+SIY6rFpDUnqEnSzvqclka5shwdtTvPEeG8GjF8YrT
xvFCDhgnGr+LPoMetM4BSKua88MeHV47rElDWXprLHV+dMv/x6/0brKHv/UFTMDo
fjVmIXSlMNqZMuelwPBAj6D0irp7gYTbX7e7U63qYQA/OHhGOKQxsbUC7HNQ5NCa
zvRW9DVMGWgT2nwpzxyF4zA4HALjYJ6PSlghK36RmREstVHa7gm8SMsxj0HlY23Q
wf7TJbjSbb3uMIQ2YA/5EMxcduZVQ33heGXns6z9mKJailpL0hUNLZ+3F8KqZyfZ
ohTcVWg0bcp+RX4AOQVMMOxR2xGN0DCvVXFguaUiFyl5mcH1YtPvrt6di2NXvMdm
0UIXTPjv/5fSmod7VkqzHc1IAQY4H+6ITjPIPsnlvciGq0bqLujUT6Y5/j0hpjzu
aX0ZNIXfJgpphT6T1+XpIZKoKny9w0KpaWHYaJGhqh6reDr3QrMKsQJOrJvxtMeh
jlPs26Z8BEiM1REFiBgUw4KpHkNcEFzfwwtKN0v1D6VQ3OckhatQlEkeNbvz2AL+
NrogAAHm4xCbzEAmCJJprN1aFkp8XamlowGuHX2xWTtZET0runqlQamNl1WDkpvl
zCZNdho62QsjmYI++pgkugFE88bP3CzhpE2rV/oJzYJ0cRWftGSO+nIpDmmY9WD7
tOlCRPHerFtt4TlIUb08L3Kuy/7eSsGnzCO8qcM6+a48QBbYf5v0z2L0NfdY30q/
65Gk5aL7sqNJ1cppZ75ios7KCsEpg6vq1Ie5jDQZPyciTCyZHdYBMFReWwlqfUCe
izwz6EDhd2m5mTL46CD7zPbkvZQt5wqd/m1txf6BRXAN1ejdq5xYHrYCHeDQd+gk
UOGKSmQpXEqyf+0efnze4n4hi0lTx1Kh/+zOdHYOEh09hWYYGVwetlTJ6O5c7jFK
3TAl8Xbdk4dOQOtbTxIvulKSNGpYlztPPDP8Q8/6b+n4tB3hYJHJjfEkl9Ukw4eV
wcKMj3yii7U+1Dyra/JRjCvyzp7X2b1Ds9u4f4SR136oufOVNGwdV6d9nFDJsAMB
FbiYTCeB7Lf7itn+4wnqsakPMs3vDQ97djtLK74WRdCAeZhFYpkDZ6PVwcOpU7df
+3neMn4lL029KrV35irrwHZuJHc9qs+L9soz3918BpSbdDsJVqz1JjKXVH5f6zZ9
SodjhTz43qbIfXQ5gCpyhu2v79T/7fDKzYokkcZzRURMR2AKMtRJV3bzGlxogofO
xU7V58hZT69eCmr6LEV03UH1xQTyy6r2HNFATRJs8uXJl3Esa7ea3gXmWL+aV81w
rJbBDpQDTthid3D5GX8TNzlJH9+YlKCHEVFMrEtM2+1uvqOKMfFw4B+iv61SowBA
H1oXBrwtu1cddxIWxfeh3Vmc8fw+fSVhqnXHdx6uWM2pOcFNop2jV5c47uo8dn5Q
TDuFLvZkuHABMw33TLr76yFaNr59lgx+5Gq6DLn67ZTScnLvWHLq45WuonUk3+uW
fORKSH3REVCDSGiGNXZnPYYRMWRF2mGf/nYJRI5/swYZenmJ4D1c1Mat/4A1oqsp
Qhvz5iA8MbUALPWrjKPFYUAJGBXDdXzbeSuHK8vlu8Xli8BwR0W3Z4AFtsm1raCB
Yqr3q34RsryfS8gZoRUBKq5Fa63pvMj96GwGlui36X7L8iLUQbf6PmFmIg/JLjNO
0w7DtpElvCS+QE3UV5xs2jaW4bsPdEKe9t3Cm3J6M42zIPSKy0bYupvm3YKx1m9Q
xO7FDJRw7CD6tPHjSBV2UcTgbrec7wYrT8wkdfGOSny4+hlN/re7H/jn+fv4EqPq
feund7kevNXq+HoeZ2+RiXFEz/P4ZtwxlB438nqf70RtePp+GMB0XrGCXB4Sa3k/
nwVkSvrQzbog/IPn6zhC2wUMsXJfJJ6dkIBwcsu21CwqNxUHYoZ3CipaBqszzh4F
x/rsjxEzp2Euqr7buA6HMmUkAhY6jIIH8/v/v/LUoOAmnDn+vrDRQXzoXXRwsbB5
i1hC1qW1mtxjv0U7or9b7sDtzabi0Go9ODfLv0yXBEo8X+ZcKNBAQzl5awB0Spt0
/HdpFJh8dffvwTR5x8XtA/b7SmmWrJZvdS79hj8LnbMB09RXaA2InPnJxiqx2O0E
49ZB+gs6szM7iGvQSttsQ4vF1KHvdnnEpvnVMB8juB9w0OoCLPSL1dTEusG2DMfW
dkb+xxN2UBLU1xn0iQNF6szbxnjJ9P762j9AjTjit0ahvUmJnTYZFfp4Ajau3JW0
tRsGGVtjmKu3t4JiyUlVhBWzeP8VQst6AyRkbQQTkc8QoX/jBpaQww2KZyOJbeK8
EI/KEuI9kB4Vm3N3EsoZDeGMuy7umW1aMPCYI4GPInz8cQ1Fn6kPz7ptYvyW9wPh
Ajo1H1SyVQzI4zwWtCMU1FU2eqtORRmY/lw2VCnibcHNszZkVzO5IynfyNt0kUJS
2Do1zmKypCjFRkoxJ88gME83Azwo7eDoh4Hk0WWnjTH/g1+Tm4zmbfKrolylc3FZ
EgsJnKWAPMNXk6r26Fqv62K4Mmfx0AG0QSDVSiBO5kftkqBwE7HI5NvYk8O7E51N
MZtOzufGR0rc44yJMnz47BK4GJDZaFLgWJ1JgqiDh21k7CckK/iGN9yzZHvXoSIi
MQ0XDznqs0Dro5bfqNQjZNPArp+Ni4dIuxGRJSSuQUrb5WTn69l13BsAXmzye0Mg
dnrt6nKAOfhkNvJ325QtdC3W9Xj164F9YCMRvdWRh+K6vR0SHeY2WpF22xi2SA+R
YqReat+GVcBwDrFKbT6EohI7KkYsOl8bf4WZNzmKq9KMloNm4DXIxIkVC2fTr9X0
VUXrwzFJQWHFn1qWXfTC90wYJQiN2Q8XLNZJJ0flDFye1mqvgjTutm8hL98P0kPn
6PezrQ4n64kaPvDEMkySWxHjZ8E1GTu6Q8x/moeeDy/NZOvbujWuy1pKRS0yo/Yy
xKSOa/EGlfFCAj6W5ixDT9HEnJoHtmTPn15Jj8hV9BRJOk9Qsw5NPnhvEbh5rdtZ
aKtZ63JBgCelidti51lFqYlMg6zC1DARCBTmlP76KIh4rQM8Xw8DkG1c52xlVibd
SpTatdZzdTK5R5qs4raY/RyTHPWdk9rOV42A3Z+f6htNr5+xmEdBcCX2E4jdUdzc
xStCliSEuYsYb127ZhfwztPjrm1s9C1Uc7yMPxu0F68EjsQbKr8QODyArsR5vQcZ
iGs6YFBtmKPEjfJYSiGr7XT8PyO11wl4nXWCSWsxFO3xH36iNoG9f6VTycJk1Nv1
7afGwrN2jWY38B5G8V6RnPQbdSR0eXuqB0gNMh8vV7Y3iKtTyfwtAw8PtgkPgU2v
C+Rukc1GaQzkEJnKK2xMBif2BOs/cCTM7Oc7KvTgWtCmQXfVeRJ3B35EPCxgtLDU
38+Vn6IEiyuMYLRwsCLUsw==
`protect END_PROTECTED
