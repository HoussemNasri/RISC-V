`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9onuwzi7WoMOjobZOjKZztBNKkVrRc/AIEB17u7aoVvYbB5bK3pbexpoxEZZxd2
XWk60cMi7dZ7+T9UkOdrT8NavqxZFj04NiLwSYbkx8aqAkFmVg2kZuejN0Ol3O0t
PZkBHaJzScMhqQ7Rv8UYPMy11CKlvt2N8L7Y22CIl1HVpOZvGHKJ1PeJi1+kJjPr
VR1ok5WSm54eYQLS57MYDd4zdLDdduvOYk51oPPErwsSofH8wFvkKJVhFJOUZgGH
Dpi0BNLXbg+L9F3fPqkQ7UuaJQYEwcbserWlg8gnW5nh0xD//pMXsJqRNqOganao
a1Vd3bWxyrwEYv6ZLQitGYgHkqlxvl8/FbeB5XUFnwKwEPa3Y4XCHmy2hi5NHOmc
keI/aTd1opCh6ry/a4J8H+G/h9Oxhm0j1L1WhsDr07qkCYcEXsNGUaqzh15Liu0c
wFFljGxzdvfZw/zyUBTISoI62F1TW3475ks9Defw0b6wl+KPYZLyXhg9IofQYNu2
i3bhOKCX3OGZEeLtuxWIa3c8N6lNIHientEHwYrpNM1iY99BfrWrji0iIgapKpwh
Jy/LyTX6jUl18pgSenZEzEUi3lWcWNpxpQQNWXU+7uuKoTFfAfZUNBJQAc+i94n9
+JyKt6PdwPmUFpziK/avu+d+8+30M+8vgqMc6bqu3okZOphSEW2Lciy/J4+2V9jp
kgaGH1PR4bqsjcLDh5v9hsTmM7ID3+76cZ33dl5Sy55XxA7rMx/bYOjT2Q/AUMCT
XBRAnUzOuaa/i2fzrtrQ5qvZLjh+EbAaX+wgTwOhUxM1LoXO0TeNLjfpzWRqEqTW
b4Ds9p5ay/Ms4k1nsjZvmCtE/Hxq2flqjOFO/IoJOBzQn3FMmViwIDF9Wl/vnn1R
kqVRCz0yhANmFbPwrST0oJbOB3yrp0k5qzNa6xUx6ZrmpbgYjMlSrUCobzb+L+6a
GDr2JIfMGzkJkcbKgi5aDvM67CXljv0r4+4+P/LtBzMRP03nkbWdkvx7+ARvim1K
xl6q68NgHFKBAHhTlqN5q2uUA25zaZscF8hy8o4Xzb9rDz5Jjbrs9Flg7DMm3SIw
UTvnoS6T0aKJdNibLKDlHVkSxPytvuoQDOe+J/dztD0TQiUChYQNulkwvM5chFlP
GUy2dBxC1N0B5Iwecl++oGtNmYdHQWkUa2RwHFPUfntI3XVgKjz1lMkbgOXtD49X
SavfWLis4up1Nhzq3PwPmBG8Nq006S3aB6ZmyLsvXiy1aq8cSFJ+2AK4uHqPkg6A
OgMIk2ul75tsuu6lFkZODi64W1LpfeGtY7F0EUcV9CH87LfjY0h4oqJX2EqaphEb
Av+lSTSoDH6awvw1jy7W/g/OTtCJ0s1VGYKtzp5a760njMGTos0wbdMygoDot5g6
kziRgFnSpxFTWSR6SybjsccnyFpPEHmiIsp/AV/cbIrovF0Sj5yL1bMM0qEYCQ0g
lxkz+ZHLc8GR1tafAUC8jtju06f3TW8hhlAnTKUiwWh1WMO4pyvXcTCuRg7wcXxK
755mqFQ4sjlTa0gh7ZHcnQwRcSLAVXcYig765l+gz7Nf8KuIQCwxIEGHvW59QUNk
cN1US3fptFr1ejHbtAXJIQ5JH6pMqgrirSctyDitzTzwtV6j2Wz+D7whgjP+owUH
5ded0gggdR1M6fak2ANv14Oavv/9blLZIqL2/thruCL2dfd8eix0F23DFgPUadX0
KnsRS61X6XDiXRTXLPY3cvuzLSyHE3gEFsvDvUmNEHJPQ2RMfcBlRjful+iALF2K
WBHnzbPpUOPfd72p3gcTtD1ZgHpeJ2q9hPDT2DlPazLDe6BSzuXWC9DYT4zyTn5v
VVoaOEac1vIqaJJtpPlEDp0OF6PqdLGbPpNQyJs9Jpt/YY8gjIe6cjEwPd05Yv9r
GnK8uM4Zs3nS8WpQYRk7JyclMotMqplxcSVu1C9/t8GrNOMUTZSYwb/jbQfBM3ce
0AMKu7r3G8OimCXRJTyUOsbbvCynsLeOLf+3gcYQRhjR0439tPkvmE1wgKWabXCe
5dfphsqM0ESO7baVat3dk2nxwFKxEs/tUHIZi8DJUXumB2QO+aXRrTPE6y2kF69P
5GDFvMGF8XTt+C35sSfSFXsC5qm5e4ihzBqTnNhkzI//hdEIUEFcT8y54I3eXuNE
cflx6clG8BXeVZ1DLOgUcmlgoPwha4tGgcDXYxr7DZ8ZjjIFfmEIRiqrtAKkQleD
18mzzjKbKasGBp7h4MagRXhVXsQJHPXXmPkTalUtHyz+Yf0++zDw+GUlw5M+jCX0
CLlAwnkOMgTUpQon0+YBSWp2RFNJdbbvGg+sWyjCjVhJOWA6v3WIA/6ZL5kga9C6
g8tcEqgS0UdGmmgKwwZTXvZdimPjFuK+v0BWaY19qQO3tRyWV0LqoH8SuYZADzO5
EhBWAOSMw0lWdesevfLmSaNmoNecti62xcSeVjf3mAvEGjV37SrcbtU6jWWmHV0/
M9RoiiO18tZmlfQnHPMNi0KOGZOpdJTXw/a2DEx3bhHwct2+vq+2+6XhZg5UD0eE
yPRRFUJuMPZ3soDp0km5KDzol+UV3cE+vRXJFT71z4nmY8vEYj63wQYVaF1IcNXE
dVmeZ0/p38gCRMTw7lgBiD6D6I/vx0BnsSuzBJ5NeDvUozjdUt+FG9nS7SSAAmR4
3AgQ//yUOw1UCxPX7S9L3YLeDU3j3GylajBPjIKuYpTlMu8d5jIftp5Pt+jybwto
8U0n145T2ql7JvIkqOcymR8hHw6zvxefLXGfWegsK/aeB0TQ19Y4zW4B6w9ZAAee
758bXvRg1QdDTZ6eDM/qsLbQfGKCHog2JmWXJvavYbN2z5ZLaQkmVIm0RmqOSjmG
lAXma2Ib1oLYPFSvXAz0Iyn1RqOXc4eM9Sua84to6gMEkcVQRw8AmmnAHwPnbd5Y
O6LuPk7F0soX4fzFpH6Bsy5qHVVBto5l0tyuPo+uFtXDdhy+lp3JkKRWOkLgPdZU
YP3iySCu1OM40yNuztxYe5wxO5LT0NeSl4jF3/wFwEksQ9D7SwQmInIHkRcAVhtu
l0evWfmieYxgRfZMYtTR2gx1F2Ku87Y0RdeTUte3+H+Xa3OAMDNydZi89niB/An1
5id8ZkITs3edUJiY6cwSHLLVAlspYEKjq3tRacswQiKxKXtphuNOUEM86ehXCSel
GgOy01os1el2NwbA7gvElMXozHlrQnIK7Wwe4udMy3AZUTNIubMD6C2n6oZnvVNL
68n1mAtJlKX1RA0JJR/jcyjuDsP1dkIEtVbYpQLt4V6TV9oXD1F0N6WOoyceSPN5
W8F5I6KAUXuSag4IZDAkT4I+uME177J9KmBaMAfKwxKTBymiuNdY9oKBn5lnBVuE
ejE5/V+dWGJCtSqbnyIG8/iQKGtCfz7ba2b5BUpFSMbbuiBGrR3IdyuR6Da5/CAf
Ugryztz84A1lpoxbcthcM4XLX1KnYtaaCIiNdHvuwXbP1W6ng+8mjN0UBuE/oykt
ejLHHZgRCUzaLLp01eO17ENNw3fRu9/d824dmjSAWodgobmn36LCAIQLkkN7VojF
q7sDUUgI1oaxi7/YhMeNz/nDphKhRyUP4UGz+R1M7oeIoQUApWXy8yjmzCZx/WzT
2DhoZ1hjvF3vVXvN9A0ZSKRiqJ7Dyw29df1YleD760hqBp0irRFtc1Tc+pJdI2g6
q6wlr3wr7EYeKEkvKKMARYMNJBv7aB0RHXm8CZb6l3tLONWqcKzOpjViBPt//6P5
UJc32sJpOvUiOWh7PtWJeYQ4Gbx6HGWdkJr8seivWp3jicPTT+yU763CHWXKTuoK
0lygGNY3UfQh7Z5L4FxTci7ea5L0yZKgwKyX+vMVz86sA9Zq1a/Qg746nt4QKoIr
CE5t7KQlloy0r+VA89ORw4zbyRd5Y+we6P8GB6BUe/F5puuZHtuCJJQn3K8Os4Jf
0FysC3bYw3ecfpDKloVlxrB+q3AKC0KgfiXG0Tj2Rnu3Za+jbg18N9+6TwQcHja1
RJD0lUwoUcpTWpm9hNjOuzBIpefHy+LdhJINTCcxb1IKI1L4nTvtaYmsTb72P7/j
uPoRU0GYWNyFulnxzjfavVU1xjW0FA7XnxEYJSvQNu1JRAtyg/7Wh8cIwqiCN1KH
FhplmSbL8nDBoH8KUVOXa2G/qj773hintKxLHJgVJ3zT2al8zpNNm4xHOEi8bXHU
Yu5nJsa1+dxIv3XR9CRE/l1fM/9DyR5PMdzUyljaoL32DrAxqSlPJpqEfEMerBJ3
P+Z+LTEVk54zLNFwU7QTTUUyoYroL/DXOJPs0cVadvKcOOjW8GRGUzm6adeEoLOB
KSnIsQr7SHRcDEXxLGEUVBxXE7YzSQ8OeaWEjx7tT8YZBhoCM/PtpD4v3lo/lK0y
As7WuxGbBSC1OGfiaexWXh3+OOhd3AvpnYjtlpr2huQ/T7D+JzGrvLmsAX6dcxV2
Uwz8z20xFYbrjU5g3wa/W3rusBo+yEhwE88XSTG1l1md1dD750z2y5hW0sja/DgR
sUpn2oaZelDHeYbUbsDk6bxYtQaIvcTNKHPlQMEzC7rYKGoTCdDkR4f0rVzkhmNe
u4/IHRo3GS98z4bhKWuoRX8MWsMDB2qQNMsXScqfpFHO3ivKIq8V77mK8jsYYcbw
XDg+DGDi37+8dqq4TkMBnYrU3k4lTJiNh7CbYp4vRbC1DwTNYBl9Gb0PYDfvgOlB
lD4Dk9dX8aDx7pNKvLw97ykFLtBnrgOj/PpLweTVB4X3Shnobq3uQJxPVz09fpbR
APNlyEvOjgiV/1l2SqIxlvr2vBQ+cSQ7lzDAoLvAlgsD6tIzuzbz5TDDaey+oOcI
77aP0AFi8ZXhzLBAYpkDmCsn6kfuBbzdfwKPd2hb0YZxOdIfFpZfrWxzZ543B/mO
0OWdCVyly2f/SebsP0KN5S0mYF3TdHQVckVYpACLLkV7mR9QmVxCF9JCtFptZsR+
fE6lR3vw4Kwhwlns6k47vt4UHe02aamhh862xbDLAuf2O+Rf7/6za11sEKp9mVJe
huSm7GgKZkQ6oMejH+pdL89N+lh2/pXxHOWtxyqrtuVu8/1XjExxxyQe1aSUS7pF
/Q3OWIdNc5nm8RGNfG0tIo6FDRCtCyutsc0RTWvToNKfcY1QYZ3Hk6f5/YYu5AvK
yiMsSUThRv2RPIVs5LxHrYBc/BnEWkjjDZmGc+ClVi43kBHsWh/YYWIh7KYlow2u
PYroTFxxOuSIJgOOW54oY0NiKvxwsHy1JbWoDjv+A8Xb41uM3jWJ+KXIfLKkQD9Y
Nna5Uped6vviLp62Ufmmez1BCRTXEo3J9PxDTJvJaNk/CARKd4TeDnTyFlSyX3VB
ZjUHON2UFujzWarIvIUOwC6i8nty5j3PrzaftCKSa6dXfJQk7+cCymH1tZX1BnhX
AOe2rU3dkFldEy/izGQiX/eGBnl/kitLqzNKhQCurN2mF9LPmH06mbHv+BmcXzhf
FfPNYcuX++64khuOPsZ3aw6Py8faAjrCOKAsjSS2HAuF1iLuZuroJ0q+cvinWzuj
uQnTNonrK4kJRhEV6hVKbDxC4WctJWFrRxMvZUFmCBauCZa/NA0AGOuM4dHOCRkt
Z1QQ8Tx9aqkyNXXUifnu/BZlR/3ZA64GK+ua0yk1AhFWm9VEJdDB7jjrmKwMPb/R
guxmGKJmQEiqX9DXPn600GYvgCHwsoFXpjVs0/uMplRuwg5dsac+0V62YlR/fHnp
Btd4VJYfDR6XwLULoT3NRaA9tbrG3G/BLaYGgGqVKkO1V0iNIlI1WvQmfFoPjAJy
agiP9pat85yUwLsJrFRVMKD6b8vNh3SBOEfBWdJF4SNKUwL2Z2uskOocG2ifKgaQ
bYg8oUsoPvZvNarE/kn2DZxwOvMphdOjN/Ltv2MFV2CrjHle1slW/MEdc8LgcS6e
OSJ/FlarfoIP/DHfptNDJTpCm99grzU4Ifx6FnrfUiZy2zTGqDnYKP2zFoYVJQ+U
M/p5ky2sLnjrmEKwz/Wl3namN22bNUH2S54tvoh87pzjnYY+5pstgk0ffmQsBlaU
GwT8Cd408/+mSFUJajwalBdICPFsQX7PSNpUXpUie36BdJSX4UjyAh9PyF+o+Hac
r8hNn8nXVHPk+ugWvhdReA==
`protect END_PROTECTED
