`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gjl70l29MSfkqeadhEz1sCxSBqFIpfRs3foSS7eQcdZuHnbUuBL9LvBBnUMkOkw5
Ko/VOytF+X5zWfxJzogTKOFY8apja0s2WJhxD/6UvaLntvPJ9iK7gg4YR9/1hNZx
4zygumnZS3C8Crc46uTr1sEc/hPMjAN2iN7jSXsAMDvSK7Eg4rZ3GFfOW9M4iF/S
/zan05ChF0hkUS4YdfIg2TzA0WqCQ3hjGQcfg1xQ21Bf+KDfTfCSOkrLMyKBmLIX
hdaHU/55J8uJu96b7NIm5DmcFU9wtuN8MeERz5twghkbqaXwH4KOPQYcBiAlW4/u
p+/X0x7nFqRfp4HBwIUZh2TLEASRzhxsvgFeo5LFWhaxBGcX55EvpO9s3bbywgmQ
8aLrUZAzDg7tb2eTn6wdC5gpJ56lOE74E95g/TTI7soxgDwC2GICjmAIg5s67sRj
kOQ7easwLY8X/s2YotM64jREkmOG34zJokBxiX3fFvuDWJv9VHvjr8vdEEwcynm/
WD9C0paXe0a7qze2JbbAjTyBCrL40coM7KL+Za2RInvKT9BwExKEIQK3SW3tVzeg
z+UhyT96QzLDLQGIxyMwT1WDczP7DZildgskLcrv+GMrhassq2Zedn1KgmtmK3L7
KDe2N7JNhaqZYiWY4jhfDBV+txM00VItxwaZvsNr3k0mNX8yF8eQenr7Rwfu6QiR
JMod2klXy3cYWjwQv4s3AjbKrutMLry7MkaUQV2uVD8JbNe4Lipl5SBTdJuclxal
fwiJbVbdtrPzLRvz7gQ4dUcuLgRs68HcOJCBacW0nMgJcX+w2FiI0lniVpH8Copx
EeVEq6fIScBTaVU3Fg5ynDpzti9dbVvmRinRpt8gbmUz8crUrg61mM3Plt3lAke6
QBNesS+GAplxuIzwlEC0HJayU2JkBTLPEb4e4Jze5KH7QhNtsp2oxsIHYBx2fBP3
7blVI06DjLlYDM4fguJbLpdMX5ZIYHznQbeDtbq82E+RgqcaTo4nrdT8z1NAYBp9
MReFsRBEPclBuicF8N63qIFGTz4UOWCl+97R0CagTOYn1fTgXgiTaNLXxYTSg6kC
IhO5FA74NERRte5EbfcT7jxbd8cMQJOZTSwIVZSvEl9N5POTbr/s3Rhqg54J6nZl
77c98ci8OZ8d53lPgHwhpnj66IZqbVoPsSMYFoarlyig084+c/MybS5j/fUhNKq5
TTWKJLxHXq4KmGC4CpZps8t9NUcOcT2k3kN1ccQTsybLB++WX6YuqwS++/6zHUtv
MHNk5S7ds/mOeLUBMJEEl0PKryWfSMGOp5LJsEeeS9FU8sByPCirF3qZzvQo/yDn
OeoTMJpKTc6tlVmujGBNNXCOTuAnpfFfbKFvkRqrMdSofASBhUV1QuZTfMtIOqfm
/jU9c2l2WZ2ug5/TzjYxcNp+HcxIJjD0QHicgrOQiwmJtEDQAh5w8BX2F/w+TyCJ
UyXGaUX6A1r59dJPorf17+LISvHgK3eLvp6LdOxjyeMrqPtr4MtSXOAl103cjp15
wvYiYPNuP7J/ifr34Htg+BfNosM6K+POK++XAMPs+6ZI207+Y+2K6FBkunJaxdQd
7a7mKxL1tI+BKdbCTOucvlX8LWmQrNewV68z2PPcse9KWbClvICuGbHvd8qRvwOQ
T/Muin41QqDhg7OBTbsVP0Wh9cf4dphCekh+iXqv+rbisIgysEECBuMIWNxj6FRu
VyqabaXHYIM3E4Y9T4IC/WQ0C0YSgNLL2FwNJkd0PvbSgzcTG0lTnFhnDzytCriB
CiaXenDlPxFsp2RA1qSLUhAdZNdRikCp6hOus55aG5kJu8LMn/9aTYECr/IzHXIJ
DOcoW9n7m7fYXn+LF7Edh4E2tzAuLKhbbxPCuGT3cH3V2Szwfx+McvDcWWItO48i
5bUBjPBziUUNWdvs39/LSxsv7nyUWdeZQQfhiIc0OVit9Px3w2ERLoswAU/TYDDn
/d5WGgsI4YDRtjfamvhwQIVrGUjiWhtEp6B4nfbagJbclhPmV7s4uQRQyTqaQZhR
pYxmvVJ1dZxGaZYFPTEUkREz+Wzl7VkVB+xNs2LbJ85wzPTEFWRNLJBz0Z6naRys
SF8OF019TBWqvMUxd9TO/EvLDY5rFoKY9nUq4DuWHTsOaTBQRYt7TShOkxd74L/0
2oArNyIUSOrNu6wAhpGWf9Ilze/k2SJRdA+OeiczLARG0iFZKKFYFPQygRq7CClA
WnujK3Wi4fCvtbMU04ergqpAN6F5Q4Vtt3KB/kuHMJFAu3220r6aU3lgxQfkjJGk
KqBNxiGAgV3ZgRRPWS44F3uuwdaSVlPzedL0TXC04nNqODCBN6ZzjTHhF6bgE6LF
8ZRRMXQ2ly2yrs6XpqEuGqDxDJdyyWYV5Gpey3Jfmkex7xmuu6MPFnFt2MnANDwS
3dK6vpmi883KJ6/T/tMgfgEbDYnxwmzcknv53kc7pRYUSoFsYNvEyAZ7lqsyqYE2
5lb1WYVQXfMtkh+Q4L/GNS8fRVywL/NvamK38MDEsdvRUG1ExxNowHT0EOdqfMp6
Rl5F1DNYBj8KtlgE8AiWzQkOxMJ6mY93NVFYpRA+KkLmU1YtciF2Pu6rLi4UeQAs
qRD+wpw4t2MwhGukBRceq66OeLdkNXDpRaYv9giVMgEB0J2nGc9aQw4+yYeTZXAw
YifmCyQJoL/PRsF+8MPlh8rsAOQIDTXiXOAceU1EjPBLGvHP7Ik1GaZ6wATteV8w
9yycAhT+y0zw3qfHlaAWhhOYRaDWf8WybtW8whTRWzBjaluro5D4uwB3vOADb2LW
nfMmi3hS0m2sKToTWCOTPfGMq6oi1GuYglaPzPVAW9ns8ptTpHRNYtcY6c26w1AV
UPTnKgso6nbn8YFgc6fTtpKBKrEJzUNyXQXWQdw3EX9wUfjJBC/3/YCkW2c5orzA
7iz4KyxKAwB/R2KlsUWSKBoESpwj9lWEmmCY3Q8jZs8L/Eg1t9gaAlhJDbtMde+G
LGGokdAEfa17+blBVMvuPDT/5ggL3Y15YagfvSew+8jQ9UsrNGNkSE8WEdCejcCF
RIAOPiUL26AhCCOp8zOJs0zAjzFx00mlMwq1ZdJ3I7/yRDd/RHxDZVCyqkvX7wkE
r87Xpzv10O+X81tZ3sVAYnA1THNNrkLz2q9U4N/12VMIxUUjYbpEk9Rh546abPuv
7GYxz7X07VUfuWDUQ5qZllhhCxmJ4aQrUe8GiqPIFW2Ky/boCD0fAjIi7KVZvfFl
NNduopUylVL37Kix66/nlakfdY6WNi39gX/WQrb7tFoLCrDrjClC9ivCFEZis8NF
fufSQkWAvizkQGw9jRy9et78iGQiNv2L5cE3ywSzca/cUUNrzffh/eAFrILL+ove
Zk6bqsAyC0nC9hkqbl5ETY2lGkr5zu0zT0aRuCYbxDzUkroczymwgBgJemvcV4YA
l2YJKXVu7jD+NG3Ffa6v8m+uM6y56YQ5WEUDoTdVmevMAY1+93qNjZsGejzPl5EF
24ql1wmyRKbGL6juZM2Ry3ycH4M72HiTbho0sgUIXvdz/4demv5h/NkhvnA7rUuL
xqDByKjYYK7yoKSqlvCEI2NXNU3h7OGlxa/Ik6EVmmOp+lYr8uPddlMOFoTiSkW3
5UMcYgPSJbhRHE5WfmZ1kUrUn0fyzrmcuRQA7qzFfAfuiMKKV3JiYekayp+cE6MK
fMk2d2K9oTcXQxd7GNOD9HldKfdJ/uuUTe6/kELZ6ma8q3HTM9quQKdyhY5sGHCT
VOcdN7dB6lsbjLdxMCktFm/t4gcNz38QOLxeJoSp2iIiz6AxOsbovKQSVez1WClc
pzrDGEW01BeR6QNrif4zOehUwKi3YC1Z0iEXmDKr6xhaaO5CYuXMoz7D0Ojb+n4X
8Wk+gZ9CAUAH70XaQihcW2jH7cEgUw5fwvofQQHIxrdyzHDf/zBzIscjwMPkDI2n
WxS8SlVI9Zi7KsopziJbTWuehCbJyFIKAPyzUECDSrJZQ/ZEvg93Dx1T/S/Z25/o
kGK30H/xk2YChqqU/y6pBE6luq9lpDvUS7OE+1dsPXWIVl0JBJUEosOR2jqMlUL4
DezjH8Dd7FYie0NeNMtjyPEj3dmmyZguLhuvzj3ONJ65iPjdz77BLYs/hkWKM+1K
4mUuwdvvvaX5699k2TTT0Xu9lrso8fgxFRK5Y1pbiBl/3r1v1NVVfyvD39oYQtAT
5FdQZeJSVcYwaRCAoZY+52Drx+LE3FXZqEqQqfYpVZy33tdQe+2QRM/CDVv94JRy
7tkpWzEmKLYOKrNc2qoVfYYzvJ8kyUuvO/zHIEjMj2qrdEH4b8q9U1gGzzWSf83z
kfn9aZlZ8dJDv5hk2mXmYv+CqjdU7jPwQ1gWVqhpFC7MnnBG1G04Ep7GQmz26p7d
0vFAp/WC2DVCqkPTUl3EtHuVZ/dLd7msDJDSgDuXidXk9nhIHO9ysA/dwKL0MMAV
y+0MPS9cqOmRZHnq+L9wNVMKf3MICLzfmWNBd0B86zQYdn7KhGfZ8Bejy8Fpn9uQ
QY3VluyBCb0frLT1+teSXP0868dpqBhLEGQxDbz2JJ9/k19gswaVN+ez1evNGXZE
0AQlvdxN5hGL/VoEwnzpHU0Ddk86WDa2kmylrcdpEzIy3y0lsXK3kRxpNmPleQ8t
tZtLA1df3j1cHq+WLN2elY/PVJt7y45n1fQ05bKi/UXU3NNzPnCGmCbG1+ua0mKh
COoQRYmY8818vCh2Qmni2pT/xaKOzrPmOuM8vzhTVSrgj/uBHvFjjMox0YL8AYvM
YL59QCngj16sa1iWLMqSJiiePdFKnzFHuRPrYce4SAxkI16pRTxnaLE7gqwTkMt+
Vf9drqyDKCD4eaapfhv5WZ81fZTNa6nNaC0MB7aOOZqEWeKAh+IVglJZ/pCUR8ks
9ZQTZYJWM/M/a6qqAzuI/3SfpJuUCDR4SB4hZ1LJUFrLhqa4rkIcwjLLwVecleBY
ij1OV05JYqvkVZ7Z6eB0VU4tk2g5KA9kPsrmwo0gc78MCTjyppBkLWKrWE/oov4Z
2DaoMpZtsxhjm7nyq5mWBTiQCNs554nzVzmDPvjW1HEAkW2XAA+yd9PEvy4IlF2k
okCZ0AHzioWH2BeJheVz5c6bSUyT7eM6XaamZcU8O5SwkgzLdbcLCJFJ+iP2Scg0
RHQ+HR941a5TSVFjxiqDyBSR3FeL+yaBRlxiZso/9lrPRTbeIZ+tWMEv3/8CC8dM
ydfm1tdq0i5B0LXPHXmeVfz90YDdLe71LqTZJLzqbxikNvrLZBSF4WW5qiUNHgUu
JLTFkdt85qF6rt0TE2bmcOAAKf4Iyq1k3Dp1KwO++pRaHEICfu58N01HRiurNsuZ
XpvX8YCg1HKtM8q06Cx51PFCIqWZry0wlVmv3C7X+44rvZjA/Kg/FWnWLtOvsqjm
0bH0pw9XDgFSvHl5pHHPzWUc7VnABQnxHeVJxbdUbS2fUMoD4L59yV6KXpyvzxyl
f9qxfGWHQ3OInpm8RejXy7l0OfbJ2K7A2+kWeY0cjX4vbBG7ylhZK3lmnl1jfCs2
UwwamEJyl55hyLn2LYOGex+xGq8lCx0TKjaCEQe8+G0pQI5qEWCVRc1tLyZWCRdG
w/sM/dd1ypDlK9oMuNa71gE0mDn2tFbJLmM4oaCnPL+RKreE4paO0l8AzbY7e3WE
X9a7uHTtj35y0DpbRMYIAW0hOIRi+ZK5lqDCU8CQa5/xRpN+PqYwSlRoi/V36XxW
oOzkrPwgAFNx+uPnccrOGhEb6xNRoOQpMdmwfmqLjaKpAEEVw0s+RatUC+y3A/ru
lEy2wcolg13KEdtOH6vqumci9o3xyAXNFJGjQsv0bLgEj39H1aP46aH8lucWPXLA
fZq6QU6P5ODUsL2vA0hL8ceu5fEelR+lKUJzZoo4X8VU6mnWnDdyM98Io4+IPEWN
5ggi3OLixWzr5IZFb2g7LM12Pl9UacpiAfx7uBx0TZvMex22LVotqOB4FydQFjR2
KfjvJoM4P3Awfqpul5royV2zqOTTrAJ5cqpFhxH/Onnjc+myea92CrHuecDr+6+j
fD9ZmwWmXbjCi0eCzqfrFUCnM+rwC/zWmKTjQGMWWC+graaWxZjwf01jghOOIwFr
YNRlPL2n5K/MfdvADBYKd/CcjAd9vH/AGh4F4+nC9fOtpS6t6YxawoAi+WjoK6E8
0uowdo4h9DW3U49Ev7Ez6M0I0tXgvuyxsPwrkmRk84JJkyjOliEaZUNp12vgFBCW
3cnGfKHvMt4MPFusAM23MgavK7WOV+iTtn97irU6QSALBSfPU8BSi1H3FesyF/eF
VbihPdrI6pd7NrRlcYx7kJW8ptyuEdLbLbmCh8/NRfNOcagOQhzlB2I39yuMEoHu
Gv/WVQBq6Iv/ujLFpCTBBkPNPVagPNbvSMpUvH/DhJ+uFGqLwr80OqhZ2J2GCvVS
grr6uAWbYEJ/E5uhkA2PGhUetowKLHtjGUSjHLt5wwCOi+eu8Q5aIyZIhnHw7L7I
BwpcsRIZQTWM8jGNnTLrmmYGiTi8hHrNREPcfFAO8/hLx3FFN2TzO5LRHD/DwlIS
Z5N/GaYmW6brcCEoVMCrDtydmxSc7n5RS8rJla/BpH0k+ts2a8ZYriaZifIjItFR
/POiSUQzw+ovk+ICHYrZO4gDQPB/WKJuhE3t9RCv4WTwz5XY9otkN6a6rwFkhsf4
sJYevVryn8h3lyktNpUlNCiZR7ssYmIuF0lnqQFZDKETTtb2i6n670hDrkVSdgc7
XqFMWkjOeh+xo9KkQjRkFXqFPZlcvEI88FpLwe5i9/hmly5an0GVWllvU2sY4SIx
6FwMjAbC3mzHbCyA6JqOAYkaYHOyAGypD0cmWArn2iY05HUnOVFYI/ZPtNCMjb3k
TqaZ2I1wWmBl/tLG2vDr0dgPcfEwprX57ouXvywDwdiX2TXAKnF4vV5qLxQclCS6
ZDI2/J2ANVSn0c7KkKNiH5dOb/2WsQr4b3Vo30Hg1G9+Fhv0Qr7ct2wn4YRy3LW9
WwYMY5U6z4hHcqXCGRtNVKbd7ZgJTQVHsQuMk+5qWtYL1HjFDkuvmOOExxQR+N4j
et9orsfjM2eIb4ODtHA3oP8ogonan7vpzkwAVwSSDvUEM8neeNmLZH72BduTl4uP
946qpEixRbWce3RCmlUTc1s3IOHO1Ols+ayLeC7Q9qUnR+VrKkJRx6Duc8jRpvGp
3BQaHjAG3sKfiCftscB7fXDPXxDHCHewJhRphXPDvEnhX4SbSOrXVd4cbVLABPV5
Y0ZATeYvT/gxo3uNCqBX1d6kYQQgpZ8Q3KZbn0WN3MaYPFwpR5YUiNgPQy7/2E7X
zhseMQcnlW/VggPPbX3TusbUqG7yTN9znqGlZLj/fK3gnbBJmwlgIT75GtDSuXPw
Joa8czprmNBw/20HnEHK/Kyiib9zGlOluLhiUhGEkre9XGA2yYYRgudBkiT7nsbv
dz2RgOr48ArogOdIyH1aZytyMWk4fFuNEtcgg76BSkEcETesuUh6CzT2ru0wC/bR
GXazZdwN1oftkXLE+uiKbgkqM4HA6zK/pXituLjqxUg8KMXM6ABw/9RTBFWdfXsB
po3KWgEIBKLtc1sESkSezlQY0WuJOSI43XLwnku+lawh8IvlpruVbHUn3MCXN+KF
xEWKLYm3Lv7VoHdeTJcouMnqy6B53TNzBnRc1pNIIDcKd6vmDd3aW5Z+9T/aXNzV
o6Dm8+j5x4nC/TjlYByAwnVInu/41P95Hb5mTJNYzZG104bLhUXMYayNq8F9zHfR
l4lbH+Jpi3HjU1qrtTQvmie19Fd/H5GQxfvu+0ZdgTZeITRWSMWu+KIBKIhyd8Aj
mMShpttOBFqP8MCKzSZDtU7tYeD1+hixi7WTgjrmU2NtUomNN6qJfYh6Ny+lOSdo
JGQdo6gNUf4vVkkoQlzZkScdAsFZhqRDAUbQPzjSr7gzRbsIoCrZ6NDVepxZob92
4h54R9/xuy69XVv4+wEEQWJD+4jftPL9gRE8S8RVLzd0TCgTDpinGsHj0iHCOeJ7
cAv8h5nENyFl0nHD4GmjDijl/i4L6JkBU7Mzq5/TdqffaBdDhkOk8J6URvxICQs9
Pzq/QEI0b3zKBS3NACeGY/TrBNoSM5flio5ehQ44A+CYAYdqK4B3e24xCukjkTb4
7GfIgsQddcTFvk1/ZoiQTQJH5c+lkQNGzPzC9n+wUVmpinuaxuO7ZzHq3eGUPVbI
lEcFRnpYAPUWaDBmBBL3zneea/y7cBoz3Ji+7B8u0qSJW+yrPBav94pt6tbDiNp+
Wk+cX5UHN+P8ocqTUxuYgWMkjm5mSFeh321PNheMCt4mosscL1SnnTNZulE/v80H
v707m0Ehl7Fhjv9dr9wwgl5uoMZkRWgmbmAr26Er6PI7IQ37fMhG0SecQxwWmwza
Lxhn9XcWbH7IH0IMdPsEpQcVeqInhivHnhaX6xjbX2hujysQsWmYDX9NxfoqQhRe
lx0e/7jJtVUG954Qpbpejg8BxLS2hVR5q+SS6aVErh9dYPPmXtxVeY97cPov6lxT
ZdvC64180zKRMGvbIXYAcMvQeM0JzwEgJ/gA4ZuJ8nekSNyF2PLxFWA0tibOAY8m
fzHzgqrLhjdwiYssDxKBVMYrCMBniyxaBRW5lfmqvK5UmY7raSyy+mCHwrr+Niz/
UPbyuriB15cqTO6yVDRXARXR9mTOTynJM5T9gQDExmcIIBTbm+03UBjeZ5ERqcSK
zAy0oPB+c9QEXFnINKcWwUGfakw6TKuAT2d8r9X3v4UD22BAHOm6B0h+jm9QywLd
XchefJFKKvbc98cWrZBa0YXcyGpvBQqi143alWATfak3dcm30+wRZXCPVw3C6R1i
dxUa5PipOBOFgXO5zEGWQsZaT2JkJDdFSyVHg/XsxNZQ2GEKa2QE0TbWffvgBcgO
L7bKI5jNh0Lb80roDXIPBo88KAi6dSQ9rTJDWnJgK7QIeZ591/NzuzUhjqiDluCx
NS87eK7acais+6kHvvMYGIb06K23M38ci0YSvCJ1wGN38ywM45UfOPzEBP0PXnPU
75ifjWAjSSwDWerB9V/xPXkG9+1bi1bJGzGO6EPqFNg21TBbDvIVwlEdNhK8dLiH
MSPfPkwGcXhNeVR0Ux1YrfYw4r5ygkbif+1QqLNytI4IFP4Q7kzLmTVdODUMmrAM
Agq0clS0vC39HGF/YZcWUol/X+tpgjUDXpDoiBWkTkXaL6b6NSGKOTXcXuJ+Hacz
QUp6gb3U9zPxZzNeGFizU4dru4e6BcIijXGbgI4Kz8uDgYGdgt4LtnKq0+fILt++
rrTBnHtR1bHHhfvzH3WESq6TlpFP6k1eOjgmk6GMPdoFf8ikG76Ad1Spd7TuJ9lV
hlrbBgknK2vJokpO3AAEQTsWiFkRmSXFD7X56W9yu5vvuCmqfRY/OrNUp2XaXOTc
eb46oH5N8I5yjEvDkZjhf2Izl+LErNviK/UWo4O1eFfWXOJOI8PycrEnpMcon48b
MM+JrXpuOzxMBoTTbKAC63L5M/kBRMxxW1KkP4zRBirgIm37cFiXVYKuriyZu5Rt
BI2Y168P5z005H3EFB0AP+lyT08WboRcYDqcZZhB0Dw817VUF4SthdBXJfZY5MJ6
muAEsZR5bVNP2CNDvSKRT69cC2RNFqsgsm5Yq206+3BrSn/wAMQTKUinwPNkVTpy
KWVDEAkfaXpdBBJHJECICIhYszgLGmF/2fgevyFUfBONcO7hQv3GeNRecxFumwNK
MqtWaKD5KPmyGh7OUDxeAwC2VZaU/Plqf0SfGF8e9mV9Hl0CWLAc19fF85UShtjN
eKYtS7+wybJ7dmA1EHt0pugF3zlxnYnec0K/keDJ71029ReUYC9vmuByyE7ODHZi
WPLb/K6xDvgcZ9zfx5jzB3mwRiuru3bKAoQjwN8NmoweNB+6ycdk6n4cWwp8Zf4r
lClgMXbP3nD/fkpsiJ2bxqjMhB4eGg5tXBaQdbkIL6enE+Jq3OqNc90CB3Et7mzz
j3Hmx/+Nn7zAg0CpPm1xmJ4EbzzYnLAqPMVoXPskt5bvEaUbfUx9rQEaT0eC8Lba
puhPihUmBppaTeLELao4/xkn7V/Uvi4WVBic12kJoK+gzSv2iTeqMJ4KQYqRZqmj
tgQVjR65oUh+1SK8NIktT1mzRJ2UcphKDatMRttVlBBFLMTLpjUey7EQ+UFgZwtW
k3y/6kvjsZKcYe/uqgIedRTOcsjDb51VgutYa/Sf9Kft0FYO+UeEbw6p1y/nWFNM
kzw6pPsqPzN80EVrIpg8//W7PNF0u1CFph7GaHrhxdYgt5b64Dxlp2lhjhIdzv2S
mFlVLpyql8B6KuSUh+fH/y0tSJ2o4PzaKt2Id9xzXruu39WfMGep5l96L4T4gE8d
pqjRsVtFnJoA3iT+zFwlJwt17nnWQv3ReozR7aH3yIM8a9uzR/oLl1vGWdDdCUff
x1YfVaiMHAiuul94MrFCtL6Lwe8l/yLY9wQxBB5P9lf1v6qfNYxizAZZl7mDTfIP
0dT2oVlAia/Q5nHzLcuKSsgH1ta41PcZoaE1qEuA0L5tLR2kKEFnsLx/jyPYXtcb
XAXBPhzHtpZhSzvlVilcK2gJILYu4+0X+zjWYY/1zr6hMGUsYoo5h2RIuPm05aD4
Qp3Wa8fWShEEhAWh8uU5KjLUBskNg8lkXrAMy0k/pX/H/LWt19F9YQS39Cd5UCfu
HqtaSiroCHkWslLhO5xShoxHhnwtwHOqeR6qW5+geHEHrY85ZyBiAGbzRt1zR6SJ
Zzj7ga4f7t/LJQEmJL5+WCTcB0ZI32GVALDS4HarVfJn5bl1QjQLAvTZiDFXegCG
pYmQjznpxRIp1+aA2eOIE1PP9kzRnMeCukf76QW9ZhilKF32BKFJ5QE08zrxyJTp
F7XtbVsYYspeElV56m7QcFVnM/LlMaOsnbGP2/3pm4sp9iDCbibEvHY2kCmNa5rI
p2lfagoTcT+7JrTpUa/+9r4ss8GbbaUXQLtcA48jYC4g4QO4Iu0dVZ+RlR6pwG0o
HsDgWnv/3RwOh+Zo5C24qwEyVABNkNKHuiIbPx0P+LwKfACJx+R2XAAMaeHTDSJN
QR/kNaatTE4WxOwL+mOPRrpZ4Ul0rI1QS1bjGVM6xViXop1hpqPY0NJuAs2CVbyA
JxLRJm6esouFO2thzahoB/Fkmes6nQCMmmfHnrEzkCO/ve/3lnrpHncXQVvD5XzG
Y3MiPwsvzVjIls0m4rYdAP/OdmWPF7T7Z98xD9OgQckRY0JbrBXSu1JMmwymHh9z
7jGexVhYweBf1lmYX1DPePI7yDky37rcxf6T0oSUC3Qwnmq3C7Ngm+VZfA8eNRgN
pxjxsLaNbBZI2K+PLyYhxX95tPo+npDPqEACxY7BZYbyJF7aylvqaKn3VrvARQXX
pYtQyAaWO2aPPdFYlrx/xdLDZOgny3LYykKO4r7mpWyCHuAm2FtJHtS4I2xzW7MV
A6dTAPQ61ye3kyrvXEps/4Je4Kx2FJmL4iTJNckcWf2P9WksFRa6EBPr+Bgm8gO9
Iw3koy5/8/82/sczHnFm6fyj+e8Wk2VnfshHXom5wuhUoUtSGJfHV1WwjxIBFDMh
iSsAJFhg2Mi06q33+++sfqAfAjpNtbRUf3h/4MSIka6Q8kSKhA8dAaxp5wla2WAb
poZ1RTrHqxXbju22IMNDDsmK2HjFyrImXXIrpg6/H+vVgMCxHWYgk2cbbsSUtJqR
4q3/aRDZIoHJUt2NvmCKoVnicM8O3xPJbv4OBYURlZ/SLm3cFwcrSP9KDFh7fH4q
I5aMqTQphP0VPUq7jgcEMHRp3R49tmz5+E+Ouu+MNsXsFy/w41tICVC2GhHjCjoF
MuxAg8kV+ivocmdgP5zieLRQQ0/ofaZ9uihEpPPZ2dGgIDAPbLYvKe15LiONsU3X
YuzMwJFOVuLJKJysm900nFKQhS80xQgyF6nweVTBB1wvnospnAoqRBTG5CTsB7e5
OYRTmOIW3l/DjBblCu45ttWpi3pX1D/0LB/imVA5HeKwiaajSBpiFUEsnWyAnpoe
Tj3l0aP6fJOGuAijsbqq8A1OdPwLkbwNYDGTT0/S591sDSKz1ViAMRwhd1B3gZta
u9shSGTe9wPZKkXzpswkgGQY+Mi5ImbmMQTEE/eYJDZ6i2UFml5oqwAoPYx37zRz
ZYgqMwS3uWwGvzzUstKtomsAM9Nn8Ku8r2Y7LPOI9u8EiwR9sMcLCneOuny7/5t7
LGMLoVu2HhBT+A7zmbdVLmPDhRbuod4OBJEyoT0Y8G961buoXxUoAaYOpaE5MYhY
gHDg5s3j5Au0whl5QagUgAjEsAKNAmGx6Ojh5pf68SH+/FkC70Bo+YdMfZb9xzM6
HIEDGm811sIvr5GUPiz8Zx6zblnSaDFEEmApTMVFO0wzcAtxrY6NtA++GH/1abSQ
8c4J/UaTfPtYXtXUR7MouryoXTcq2CrM7OG7CqgSygHbb/M+NZpiG1w3nEcWKKhm
rnAcy/SSd7fA/KPpjo3VkF3N43b3nmngxvYXGN5IlJHH7CUMr5DRegq7dRorW0VN
ahIRmEZNGlMDyBMDr+D5sfXpkoIQ4Ms1xGkdLcUvAQo1ykhvYiKgKs3goDm6ijHq
b1OI1VIVnTEFVv9acDBiODwhFdewDL5QNK3jrGW8UxOJrtcqh+XGpbBIBomZEnI3
qVuOaWfjYGoHNbVVGKhhtPhTC+/H7aiUhWfZYk7iENqHAM7zfMVOmwEKWk0DEtIs
ed36tb9FaUuPliOrDpEtCnXNJEFBNv6pLZzFp8OJ413MWWMim6ZCZ2yPwm5QSm6J
42dhK+ZdB4rox81G+wu7sLiWfgFex54iWsmYm9Hs/uAq0X5HGulfwY7Tp8tlK3FC
YogHGbL4RmI63AUA0tZdfe3s3B50lyu0ueuQONz5zUouFiHgedj2Ijya+eGNWoK6
39VxRjczXq/rmVD1wovogjMMpIca7LQtcy1sc6xc0Fln+C9/B01omBGvdERIzyyF
vdh+Y656M8wsV3kSP15VGBZRffDeNGjpCwnJoGfjWUGLXaAHHsHRi1QbbIfR1HqX
eJlWcfTg/V1CkGvGDxwWfbulxVGtCmno8SzzWsYvOdrwBOnLM3S1Z7arsbGpKKWI
sftXIIHrpR3bMW1deBJBngHfglLX51buz0dkZ9a6VMXAQqnC84012jaHyuGMFqz8
vYd724BARN43pKepQf7+o1/FbHFOABwqUD+R68GP6HLUellYiCoJ2ZzgDz8bsg0C
mAklyxYWqAIvWBJ0X9kH7d3JxBGvBsKih6/bS5neskXMYtNKwKktpC3sno2/2uZu
JWfDq8vd93ZMFw1fCIa5YE6jrWRdTOsxaz9QDOVeIMqO9Nb5Ebyr7CwPRXuTNJ3A
4vHZGoDQe/xO2M6KGmg4I0IiXO3DACKhqTHQlVfSz8j7XibdBOd3+PPGj01r0kHl
HTjq/5T8aeScCeQ5fQGnz2k3ViC+DTi1YbqWJ8cs3G4bj7sK16UnbHLUjqU6pnsK
ZRaQ4x2p4yCJ+WGFyGqobciZRAIGYempAniG3y+WIdrnsNSHxj64ftw5HVF4WaKh
B5vdawFtEXWnSrjMcUgsW6ngV9yWsiv8kHtHddgxbUrwvdwfL68azfJ1TPCdSK98
YB04EpA89LXkC2oP1maIzb5IVd02dgEZvbHm9TdRPNhU8yIBiQ7hS106yYVQ6mCE
z+vlx6w2yUVj3anw40suiUGmKNo1tyACjqwas9K0N3E3sBBcJGINfko05gEA9ipE
GzyLfIQkz7rHLTp3GBLGeTANWs1YQKcoGYXq4UhLnaCbXweJc95UN7cbd+v4FcXe
ASoQmigvr7i2qNxaBhYH1eWPeFEOepMHSuKi3Au8gZoK80RmHSlJ026gCNwuE3ko
oLbhKpDFA4GfGbUNXYSCRELdu/YQlDbRCwnMRN3IMPd0Nf163MephV+N5tjYfu/f
PQV7x+ncDz4JkdKCL9dlgE5OKyJENpTUfg9XyJN0STVXx6C1Nvw2EOmgAGM3nbjh
ViA9tUl0/daQQDbFn4QakjdYvjd/+z/IPDLbdO+o1Bg8ggayvnYhWQq+rqS1lbLD
a1EGB2OJPg/WssDXHa/tMc8Y8+/uq3VYZ73GzdoRFoufRjbr1N/6cQVN2ZqAjE+W
Qo1pASsmL8GI2l8Gja1t5ZoGlcwRoughViu9uOJuIhz4RqpIrJjjI0kMa8yh/M/p
6anTkVrRd5SBlsZRHEWurVEU9uj6ilx1Erckan5M5xq/+qjIT+GKSsE1kQBtDRNY
PQhUrS4U3XVvegHAV5tE54CTE8S/DTj3Vzw/c9dlp9R2i0E/jhTnmUj47y8dN0/h
OtQ8eMJHr4zjFlYd68JgU6yo73G/HPdctVRiEaVX/8lVhIkq+mpPS/JOoVczOmeS
L+M0rksEUVy+gFG2szDxnLl8kvB1wVDRqCLXj+L0X+1XvIZ9SKhfLN5C6vRzw1Js
5pev+bcbHhUges4KzIQoY/DVooWGRJH4mw0jWzF7DbRtiK2OXQfv9lXBaz3vaGt1
n/1Pvr5WEKNIgHOKa1jVLkaugAWAeDYITOK6yU6un1dr7Uv1AHOujwp22uaNkJ3H
rFpYParBqcZ+dDAdp4RJKI9+jfGVE92RdbEdEx/JeQIf8uoM33yQshLSscPiwNRG
4TRnK3Ol95QOLOuzpUX495kTMMJduf7MTkml6OY4pDv73h4mzsP3tBHOCSYiYMwR
72Qg2UxPHwyOpZ7sJTWvPCCSja4c6yWgWDLbUUmuIVOYOKlCIUGTQ7uYzkPpVZat
w/Jae+THyOoF9NKogR1tCNTEHLqtIwL72fgOagmnnm91FrEBeq+Sz5iNc0P6Uqru
aP4cr4eKhR7IP92fYJVbt87qEPBjdo/qrxRqNKCAgR0DCdfvioyjxUfm+5ZX3haz
PbxUa/bYDnRcqVxFo7uZlinx4dtz2WBv7iRugzJ17JNAosG9XA0aIHonfpROKHbD
MYx6JkgrViD0QtYmkJR9oPJPDfowsxgrmbgtDC6E7jA+bhwXZxNCCBL3WpbQKSyA
iOruiCVvWkHvqS6zfxwfcTn/IKcwOYnoJvbowMwmhvod5XKiX21boA8BFJ4nERjK
NKkjyQFtMQbqTsdbGmxUwLYgzmMuvT/8JSKcxFkeFCV+/Av30OzNHU5Oy/2Bf4LE
eBMinzIUXFrC4V5+qzsPvE1XxYPtkt0PcY9rddpeSCv+7lu1aYstWHBLY7UhMHpR
ofQg9aBuzBk8/7xWfn1JZTHF2S0EK7/hgWNp4ZNC24nb3WhW295/W6q1KJoW/U2f
HkXX6Gils1vhBbrLCAuyjS5tXVhaAc22qggHyHGGa7Z34LQoHiU+F4jIRFRhibs9
xjgz4HAooFxh9MCe+ezqZzqX5IRaCfrMpM7VC+jIbLDkBE+rTkivtAHmzNp0NWIp
StDRWbH6kw1o3TIKacCnHjSmY3gLrH77ADxPxgPvgFqoklSCo3/R1iuU8ICY8Uer
n3SMdugLk3z+WZUfRfDDUCSh0JeSFcDqqV03krMiQ2VvYt1iNUNWw4/0ZOG03up9
ls5Is12nZPuMhchF6YUu2cWtv7xFFJyODnOr9wwCjfhhBHo2yqQOklOPu69f09hu
DyxEFvvrX+erUqzQGBxECrLwzB4NUth1XqiZEFNQf5HWTVmnnGaroC5ZFH9HEtcf
wjI3r5/zSl5jJf+CQs01F3/+3XlsIACQMi/lZBY3ivU+5uDYfMHe+kPqUzrPxTgQ
SkiM2I9LYpmbeaF3mTKZ9/rAPEVDNyiX2jscadYS15T6y17Hhv3m+g67Dc+X87mt
2DxYSJpcia1abqbYAg4aUerNQ1T3DMbff0iYTwHVN/e84hfZKZf+BHXRdy7otwOf
d9PvlizO3WN3of/JMMzFAyJxXRKmMMHBxjH7RWKr6h8QvKCnV3ReH+Ig+4oQkn7n
o4mm4eB5+Cp8jO9MclSogREbWcS7XmHvcNOSzPxhW48nplIyONYY8mwCT7Zefjlq
+stwA5VeErQasdevI+HVA7bfbIKdt0HM4VumF1F0sY/FazCavRRhF8oyqRaZg3SP
uDeGOXuLv83BYFIQ4MvFzppOcpvEFMue6qlzJWmJmWwvPULt0n1PyxXBMJSlEjnu
1h/wTSlpu9oMErdfd5wI/35ee1MM/yFOt/sc2Aqbegg7YNMujlwAbsP73N3uT6kY
2kL0BUfMh+ECE16+QdE8aiVoQV1WbGv1lmNY5pxGtkIBoV2/qozyzxNV5ujBKqPh
xCPtJ7tVYBednSgkt3E9mLMRrPyXzRhz6DgqUMLBZdgbTKNz7KAF2Q2VZrvN2me0
qT81v3W9YuAqEjs8eqZyCfP/xkrXI8y82vV3vXTOpIUWmlH4xmelI3Rj4iF85l9F
NZSizpFa2D/dJ/Vtf9s2RkbILBmT3WfOiu7+P9PMIJVkouWUJ1UHGhb1HMDvPWGJ
JIAFcuMtRHrr0R+wV8xDIHJGwb9gC7tvdnRgzXBb6TeWrOBYLsCRtXcjPTdeljVb
UDGRNWn9LbB9PoR8f0H4kK0M3Q1F+eRP4SZvzE+AGUkzH/rlnkrF33i+FPDfNNr+
EYZZn5D5Zm2qZUly/hIRH9XWSyO/6ZKSeG/O6VK9KDfhuQNEPcGTUhQ087eQnm+x
dwHpmRB6OlBuZoX8EOMoJm0ncNKQVJuSPvYMTJ9W0qeqKT9lvkB1MqxgG8X9A10g
HKpFgQOqEkjV5q7m1p/Msp1ZWG7aV3fMlbU8UoSKqTKIzNb0MC2bC1B89pk44Fh5
DVzMut5/3ejOyiiWClBP/12zZN+g7xaCCmE5+Q5wbiG1Vz2CVvLHyGAjfk6PFZsA
cnr8Kg9rhPsr9GXKGQ80BHLWpZqND83F5PR5g6Z8yER+ivHhBNZ/aUHweT/pvW/Z
qr3aCX+ing6dU8vVJeOFewgEgzMjsoZXOAXlRoE99BxuA/RC/Mn5ItlAHQhMcqlw
lO/Qn6Xc6cqCCYpCOjWTMn2G11QYO8S2GSRO2KfJawSinJ3Zmo8x87cxvv1lqPJC
wqkiqOCM36jsI4hHSNjkAL05uzBnBVdNy+WHFH0yGq6KQr3IA1y1CqibiPqK/A6R
1RcDqVi3zx+gNg6PW1byCGTtoHUcfiLN7TX2k6Xkb/i7VbhI4cLr8GlZnKUGRdoZ
8ZC6otKazn7aku6vcfNMfRQX2CWxZPUW+88mLYX8r8vXPP0eZkc/s9YEGBqeMbx5
a4Gik22+pCEPHnRFOCcwHnIqyiUxQtlNxgD8AbQeSwWxEYkYZI+vVu+gxo6YLSlY
a86RDiTnlL/b2djcSOwndDrjYF66mQ+3VZtn8s6WyrK9+2zqDeLFgtDuBY2fhL96
nQUEHC/ItnnUeBO7gvTbdb5sep7nOxAiXSs1+Vu78WxDB5IzRIcv8cLgOVetLzPN
Dwx6DIJU+8qPf04CJeJHcSWawgwfdzTw7SEtxdafuKajdSQQq0BaPZ8e1LoA+98I
lM0htLiZDSTr54DFkx9rXc+3K4ku4+Yu/Dt9zv6p+VzonXR6GN1lU4hCXAJ7N0fo
zYn38JpK3B3SMkfYSMzye2o3CWSqJ/sfayLzxS6T6PkFOz+zP2Q5973XMPRk6IXO
I++TsD+eXxFW1TOwz9ZfmtJrTdXhJZAGnIH1R2i0EzaEx87fxuZylJ8U3IaSyvML
R8VqdUxV0nUoALCgCIDZRLLPBC7nGZypPZr8hU5y3wtsGkCQEI1I6isAal31EhMp
k7E/8g3Z+d7bUKIGtW0CkQafCqNe40YX8kaO8i8bZNSk8wHE0LbTL1sn7mHHao4V
uhJY9KQ9BBYnb/6u+wgGejFiWp8L3ZcRuknM9gFgdVxq0b9RkEvzyep4Vx3Tn1x8
pERXcfkiYRzZXmKsriZ5UvVLms3jHnthI+P+KgGt2AqpmMWM9dM3z58AWsmgMmQv
sxf6E4epM4kSiZ3IAkR+9I/VeoIG2rS6n0mFgRoJCj6cnffvhpJ6n4E7UqA5NP3W
wwQzmRf1XG7wPvgEdQ6KQUVcSPCwCPsVSvNR/BM0OGCVzKwDyGmo/sdmYDXFML2r
5WkSKflaR4pTj1mPPFmFNRrJo45Qyy4NC3Kf0WinCOVfhFkdrtL3gQ/WzJcBvsla
eeJgTz1sZdq4l7/vkHVbHjvoJRxmGo2FDrKXptL6aam4Bsneha84+3icT6O6O2zk
EvgBCDsqdIbSFESIq0xFTzjzmGUyiWMNwtliuJbXCgCcfJsF6HQZhMgg2oAsZ7yC
BHPSXhunPgIab+NutqT9/FMMyhAhMCIQYF+Z4UvQUGNFUn+g2+bH0b7hGVb9M3PF
tLJZun/jwaj0KKFZJlAaT4QIvXeJoYps2sSpRTrmW8cv1E7A8/PlMOGCqFyHeroz
9WOycnHO3yCDai7RukFt3PqMQPev+C2O9h4+nj1Yfc1VF/IWsHzwI5FBw77jEon3
j8leI5Cf3KpfyB7Qv921g9VXOPnczwmjPd8OOQp266AzzwmuwWw6vKiaxfK4fItB
Zx6+xTMqlq1WJlmghmlipliaaVfd8gcjXk/Xjc0a0a82zi9KRVa+zdJK3L6Ss5KI
q2p3nN0sJJfLc+EGO2N4ZZtQQEO/DsONK3yeW6/JMZtzCO9RxDI3TMDRK1J3yjTk
gBt5YQOHfuChNKO/a/AH/4bRj43xvOsmgh8cd0woGVUAf2OJgJ7EnPCV0qqYxm8n
12FlgfFeBHedMHPO4yOJ0wSGo6p1FWVXz9ZtK+680XaGjHB4/8ssp966qmsR/Ur0
eZxf3JevMRbuZuYqyaU7B5lTbC1FXHaz0bNmChDq3HKFFqR5tEcUlNfzfZfR0R9w
p0AMTanLsWqy3OTJ3krbr7s30GVY8qzr1hPetcONf4D0+styNP2ot4ZTm+GVFwKR
Tj+bE2i+gGcIQOoTCCsqnHAi1eFgmcNe+TlSoDfODq9D6Hj6q+Ts+Qjyl4qsgxjw
OWNegSiC9HCqqXbsM4lk71w423sxlKWxlqU4cm7sZzvUBkcTm/wip+J/JEM9+pso
Ju8axRWSwlCmMQUNeN5NORVYRCIcPhQ42OTAGERmsDfSVYXWVqnqfwISQQsQE8eI
FWTyW6Y1eruflHIZ87LesHd36SkaCOe3yH/EVImFiIv/nt/LZJFmdrdXTcG7Tx7L
STyMiKl442eMoN7CLQdGOxEfAJoFm4V3YpgP75y7W8GHRFQOeRd9aCgKYDFW0AcE
lyJoSsjnZZEIvQzmPN5UkT7uis/CaM8mYeV7XMVPK5ox3UjGi72qatzVIBCf7EFJ
r9FnMHXGI1+W6Y9zCKjnYct354p4wbQlArE+CDbxTyWZ9QVpLKVVOx4fuA1gWZXJ
T+ZKLWQkdHJRrEmiTEYOoSzzZPRjbxK29gIVkZtP2tstHZdg9/gvGHZ1p5XcbSDW
EeuGaS5Bq4mDyoaiOztBXphkPphLsi2TOCL30XPdsun7gJBRo9vMTFfKpVk4JyuD
9xeGHJepDwfLWMsDiwbE4WlXwIkXB4LmXznhTef8zJnujL9fSPlpI7x22dtZnEIo
/rI43wYL/MttQ1cEPuKEhaiD54pI0SLQolqjRcOc8LiflmhR1uifqlMbqr9gUaTZ
bHjGKFradtseQee+m55FPe6Mz//90jbFIlEf2T1ln5lvUU3DnhVqqiIicfxqfGLK
cbNAdB9aDtqIUrI4lR/LVpH8CVe40l+Pgjm63E28p6rOXiDMTcqcQaxxcH7AYNdE
vJr4HMebyNP6PEZYkt9gXNdI0UnKD4aEA7dwuHSPSADF1jAYeUROtmVaiHBU7qlo
KQXGu4l5CrIA3V6vlzpNhCophsAHDa6AYdBr3d4YZ2rNTqGsCOUCjJVyWjDeyb+y
cAWloW7eRLVbk+SGtgOTdFy/Ovv9j3jrGzhMyiV3V0F73RY1ibVqoZBYk09ixldn
Z/coK3hBfK1dQnra1jG46t1qU058yHPxwqCV+m+uPgEfVH0UK1cHHYmdeEO9BvAp
Ypb70O3jHhmRWP/s8rOOw6E5/EnsFXLpBmGyCnZQjFvfuOxLU6UuHpOzeImmKZik
yQ4JYOZXd82j7x97IPoHbO6vxz2uHi60TQARUH1OqB4hViOdS30rnhrnYQEad3LN
5dgmLiPHRUgnewH6LUx/nzzMZEQRsX2XfsorUDcxjIj9aZKDdhFj2kNBEaLNJThQ
NPVfWqCM2WUf3UZXLoh1kV/RFyqVhyt8YC798ZlEciYfbwmItt3iELHhCxOGKSPt
ZdAxbUwRkc8InXvIt7aASwAuO2Lk9EOeRU9CHBPWX0LoAkVKadXkbkMiHUhD0r3N
WkazWIV70yeV+CX0ZOs8DEkipY4mu2++fEuBZQvZ9x6VXQef/2pzO1w+C8fXpa33
wKNQc+KBb5SW81I5TiTc16Qs2pxaKkzbc8/uaiS/7zxlLTYiJYPAQZG/rY+CHx6/
a4fxpU6OhvSujM/M387x69Mx1+s6LZu8JaX8D4HuLHfxsnS4IbwrA9KyD96ThKsM
SxT3nP1l5/e5mtfkr81LhzXrg92/Q8gW6jiyTmyP7/yUxia6ajJMJHlyklWDZGNm
xz40AWgndvZWeM0seh7A6fhO3yqnaLWdnftmpTjad6RocWMbsV9kqNtEfFO3/iiD
JKSVqAVrD3jfXNoMydVtmh7F6zfzRfuhSbpn7+xwaR4tfAPVijDd1cq884TZW8Z6
wGK7S/9znAx3wYN01COuVIgziKKUGLIgTOCqIeWBflnrKFzJ9Pl0AJXi9+elQL/Z
9OwU9ksJAeYcfyGMQR8NR3LnKu54ASL1ICFLrf7Q6XoPL9j1OrHeeZ82IkJGaYoF
irj5h6/inDEJgaYx/gYF80TNfpfVkMRoNyVQ0QNywTTksPnYz7ar4DVdT2y+prKn
7Rp/xEcNaOUy0AxX6ii6bY9n6yPfMRioyGI41Ao2T9dyU6UoLTbP/O/GX+r0Ga1U
+hrFiaCnNwHUp35jMaFBDvx24qItnsrGyaR9ibBQvD8pfwmFLKD1UUaCiYpS3iw7
vUC8MRSzBpDP/hickVgbmzbu80TZ50FlclewWQFleF25Hq6+yljLhTKMHcJUiDuO
Wa8M63hK/40GrS7eCM12EyLmcHEaKIdV29qeGXmhKdwdWdpxyG5EBPH/VY2XEJ6I
api8PiYLka/bdEbxe7TkT+eGdO/mUgieIjRnQO4xK4kLGWr5wV9Ukh7d0SknaXOc
Cc5R7FYwIeeq5psrbjUVGT3493LKxDAqEioTbu992lbB9iXZJM6Lc1m2s8wbMxiE
XXoCSnb9t978rGex1oTv8BElxEzSJx7pjwWBXYsuJ7Yxlw2zL1Jao1nEmed8CwXk
usplDhezpdoOdDRyLc7nBZqnKs9CcZwrT82HUsJvSYL+m8UbpUSDjcFdWRex/paD
gtngsPoMEN7FXIc9SDnEQ7M1bnjNYsUbpNgFwBxPi7+qOYnBTqmBuQiZKkR2WX8I
SJqoWA4aZycVVyHPvDzA3TEzInPq23I/mOPo/kF/eKfY2oaJA4Ro//7+86sqTdK2
9Q51Z5qIv2y0JiDRkDVLqaygNaPE7yuialQIGBRAhz3eSW3F99KyHceIjLz34Dh/
PJe1F5fTY/vtdyyhzKJXcdGsbAvQKQRL27bdRPVlqepZijjBvApTOwPrykx0RHvc
HdondmfLLd1DZZUmw7bW0upc80N3ETODI/NFkyCoyn6vI5SgCH/1WlCHDufXVX56
ML6fFlUFsxMXnejvYKlf0vRLfBjiMo1I2QcoPT58OYrzk6TH71JDKZT5/g/4scu5
e5hgEXs4sEOeVXys2bPqyB4faWlnEJpLS7dMwFB5K41uFOD86ItOFrN+E/FBd/tS
tOduj1WlR91eUwQv+YQ0u5FF3/xmwhtE1WPd9g0hm0EdxVdc8y1leSt8ZMDIP+Ta
xLO9oUalbXGcA/9cVPdupbFooF9dPBSH7c7AewGAUEPc30OJiRc56FJEcP7Tfyfd
Bj4YQmH86rOG3grBqsuogTlMgfr4ekQ+RrUqpPJAWCHyRqLe4VdED/H/SQZHmRuB
cZ/Ydgyqs3RIq6OwtGgYoZ5bN9NLUFjgc8XlMYfUM9i2oYkTQ23EzaBMOJZypvnx
dBiMUqHD94Ycl28QZK0W/FmytXzcdMEGg4bgTARxDxUrCVOMcfgeIe+kTnGKModE
WiOjraL2YHkw9G9LvgOAjcunhFrm9vLeNQ9W/m61JM+FwpZds3T0SqSBbL0wAyD1
0cIGvcYlfi018q1W/qIRT+9Mmg3K9HwQ0aOxYGZfSbonSLv9MQ6gal3VOKQOu4oT
aV3ZjZUvdMDk+AQzPnrraXZBC1r+A7L5ShPK8CzUncjw9o3/tE4oNlnj0UVBvaqq
ZjYxpq6MH0WvXJTlqVFSUgDG4ECku0TqSs4XzbGxxr7M1z7JTdsCoG6jp37UcpNQ
DQ5YOy0m353xVuuNEP4G6XlFkQ7H0MWmgpfg2PMJS2tmwarMH7slaAXCiC8ylj82
p7lFmEgRGspaldv6LI/c4Yez7xsKtRL8e1lm4mC21mGv/k+s3S0YRv27QVXH9Btj
E/Zo7febmcjO09QTnedaW8a1i+7f27qNJUm7wWGqer1bO7sLo9S8OkJhDr7Pfhsq
J2Ww3zQtmp4x0zXpgFl1+JjmXLSWrKlBcI/xdXa4JjIFDdNcI5P2mvxVy9hISCyX
VPLwCYnNtp6Ln/DsUmTx6bMQWWsk5WGSubJYXyIH5/RlL0UIaDSWvQugbxJV/cIO
bM8T5Yy8lhXZp+nI6F1sLjD8y/CDsYJzw2J3pDjmKLzzKAVvhSeBlEzellAYtacp
LfUtALDIJhX0JvIrlq+YdW9jjMxteF0+53S2xef6bpJTZ8T3EleKYPJpkS5BfH63
Me8d9oklynhkyn/Bp5Et21NkPcO0FS1pUxFDj06IuQ8J482b3Xqx9lsiZL0hEdt/
IYs1JWYtuJJSHSSX2118vlU7QQHJTFD3tkvw1j2I4XtxUwRzW1iuWRK0q4yBNUrU
zEpd2lRgsnuiyRe/IiSevA348y/0hoxv9i3d151O8FwQbjHRAg8LFalYzMxWjH/x
KZKgkbZdxaYsQ6+QQzrYzMyaMWX1mo9L3Ut6WJv03i5GupCAS+bA6t+hCKZQcN7f
B3a9DVw/euQ5hnGPftod5xWE4DF4FbOjMK0PSWyXRvEN/wZJPB4oz+0OT/Am9Yxs
tDMeCs/2t3lpnha5jwFxDg/Tm5ysP1bXzehi63guksHftCDMsFOPPjypo6J25bPh
bCwBOIg0pzffVu+g4GpG8dYRXRx/pqd9nAlN09NxwRRPkuu4gF7SFn2114P+ungm
Sxz8ZZj85qbFO6uEgtwK/mGes7MSYh8gGt/7FZOinWRYQSfs9sCj7O3eAyc4UI+I
Xg59fqilfPKBPh0xkTAEDVuFGggkts2IXjOKjlCJMKvbP+WjOhPthHuZs18I1kQK
Z2oWF2UB4PP5jWdT7FVgh/xfOHPOJw6lU2RSG50S0gnbXmHbYXtQzsuUMzBwmkfH
a/gp7ILVsU+5He/KMwH9eFBFH1VguhwCH+or1D+qGLQ6vn54SNV/zdNjfdeuH1fT
0+P1ya3UGrfsOIM0uczSAphf47ogN0rS3AzDLlCUTKLMwbpKi+dFB+f4jJjQuN+U
xyzbVJ/mLM/KCyJ8mx4vkzwD8VzGYAU0gqPE3iYiI73sZpKb1awf8ddK29Z6JtQT
2pQF9k3f2GlD2hW/RBxeZ9KmTsy1UUj/ZNu8BZCy4egzcxcHaMKzetv2OBApcCaX
B/JE4DpfIH24OL+aKZjYhmG9ube73IVje+jywh6re4cj5ZBu9qFEDxHHyA21ACEN
64He4IFYe6OIE/U+40NLU0j/JCgcAQgt2jAgPoZp7Bufk8nk71eYXZ41bhUzw+XT
piDvl+vfFPODFl8fe+zYiq+QTOYZLQ3qMJEray83HcvvyfYcSaHXrJE7m8pvD890
eLG/lnxcOSVBM4SCfKgJgi2t2G3kzozDU1RkmEvqvk9bLfARa/OScImUJxEyw+NX
lYleQSS5u+3P7HKpI7aBJ+2Bcx2OH7PFaTkwCpraTtLPY+KCTH710JjD31GJGYtz
QiyMv24R6mBxD8nCuJrCnyWSCkVLksl8BNESQ11/iiWyKVXlIEvosqE47J41pNfA
EPWwWWolVMfhhenwmtYQFhPbQQX/d0SiM5e5pNd3YKuC4BAA57h5x0JHFYE3kdsK
QSOvlDB/jdHpklT0sIH2dUrJ626JgGFSdBbneoyWUOSkxNU4YJqEvDfGIcjNojTE
8+zTpuu//C621xQ1IXqn0rDrjerxb0NlYtATFZeEGhvnL8UqdJgsNR8IbZ6u2iNq
co1SY3mLeo5V4dq4qkJ+95aWRfbmTNp911I0dqQKEoQE+ksCy5WmLklL+cL/PAyc
0eFTtXXluFatMU3V2YBzr32FB7bDnGd1WFtHDd0s+m8BjjBjCN3uvF2eMDM98Xgy
dL1RO712BSBRUgW+ANKPGfkJu86mdhoDfO0Q2pihOWc=
`protect END_PROTECTED
