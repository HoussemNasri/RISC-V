`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61ez1aFXmBKJAeU2og2zqTs7oriQjAQj1+T1oXmJu1jNhIzowWD5piZhmj47Iu8i
Nb21H3n74Lk6685yQsqDXj1lIG3S9fQymd828+kCoGvfBAe5NapQi/H05rGAawX6
BUXBXyllF3kqo3nXFIVeVCR81Vsy0jEn+HJDMt1mp2ASCe8RkRhER+WAFFaBJ2eV
02qol9N3hL60zucSuUY2GA==
`protect END_PROTECTED
