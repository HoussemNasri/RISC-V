`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRoBDeDmva9MnIXDeiExWqMZXPXxUDEj0ohMv/4Jc5WCxestXcbQXkvaYkylkeIZ
yLcANzRPGQqih8OhUYsqcb9msVzTyslyb6nd3lcYG457LEeelAVu2a6nWt7rumed
BBDsqLXnk272lfCxnjwJL5sUtwCqoX5UXDZ2OzMoY5/IYDRKIfjj6ZOc0cfw5zCZ
vtcUlAgoNQsvko5l8eGdpTMJ80Ws2Jd3OwcQJoVKnfsaxKtQuJLH817bDJOQ79Gb
AeYcQV0aP/FmBjkFlVFY5BcKMEBcajBwqwNQIEhbO1yBIcE00pCmREUjC4W+lx40
wlliDjoI4rUrDVKEyZZoTlxiQNtNsdpOLtdvMHuKDyuY3PqLbpiAVRYcaID9xxZ6
ZObnsPgFVnSb52bx18/mnVYUgmwDsXFUVL8HQRAZPB4GxzN+DtgTIZLZXu1o6Gis
SxXdc1JWBzSxYk5vvc5r2JDDjmDkRegdo2SDUraUENuiKbXYqiY2aFT6GNimTX4Y
9ROLWumtrSzu2LnWQvadqh9tVuoH7DarGiQcSdt/So4wZhHgjxK5yLvvDMJ5/DD+
IGd/iAlhsNv62fLu+z6Tb+QNEED+HPXm+UwhEUqfcqhdv5ZMRXn52sUuDH6RjlnO
p1fJaZgDGmH9CcSteYfToZLUkfa4rOngj8p+3VvlSbNT1q0m1NNUcHIoj5f2rM0U
citpXAUXDi1QZ815XqAoMFOlwB6rg4N+zhvX4u42FHln/gTHI+h7qj8BtK07I4P+
xp6E1RmJFzMDC9k6OxQb8qpR8EO8BFbUNxvGMvTPwSWAaJeHuM7n01iZDE1+ynkL
uXGIBzXt+DyvfJ9Xi4urM8tMivK9IoyFdFlK+zgmp845JOYHOgvjIjahLhqFXB9B
2z75fnuIBRsuBQron9E89JCSgPrKDw5VV9qlKimy3nMrzx3wmpT0vprzoVIhlRVn
GU+stovfyMiTNrvHhF9jsAb1+TIQnuRjpTRPo7M6LfLagmICLtXhicp8wFVxbkmH
br6Dx5Denvgq2rHwBW3hmIT8jA2rfeoQsX04EJvtTU+sQVpr/WdZh0DBvZpYqyuA
NKbLgb4e84IatIAFfe9ouHXsvgItILnUYUS5cPsaawQSxFMwWFfMo7UrXyRoAX6E
M1iUNYD7JTPKeC8TAOVRRxy8TfZH5FgjadmhA6zG6yW2PO23Gzh128uG5zt5/8Jr
i5naCmjmNQziEuS9HECl8F+9UqDgz6/HTu7vCBdDoU3Uc3FTW5Rgtp6ShroLoUiR
v9Hqk48bMktav/4cbvdhfTg6fVwCW6cp3SC8sJYQvlAULpGlOYRcDFGmmDLPWuDh
NdOaFFjgrcwOsS08DyBCZwn+8mQF4HEEBkSjOcwqCBGBspfY69BrESM2Z1KQCwsR
zWVIgs9KecDq4z9GvnX2qj1OvWb69ZgFhivGd+KEk6Dov/2D6T676Z1iBks1/coi
Tp9jgacMnEHVMybpuC9Sznssp88AqOHHOSYtg6ieYuHKAIAtY+44V+x+p1p5AWr/
SI1LMrE4UqaK3L+p8DgM+7SXz29+q+PA7uP+t3dCDoo87lkIn8DVV18/e0W5PvCv
4B10rCwvQCngRRrrVPJHvEsH/XCWeKqXj79ZttirIUqJiAJwTlA7T3O/k1usAJCm
wt0lBko85mYLqmwYSSS3pRH4/Fak1yBxykywikzdWeObxUCtyctJPBQqL6KjR4OZ
JRGjpmkt0gTUa2yh7swa/YV8e/dRTNOEzNPF2t4k3iUznF+fS2MA9jiv57TlC2so
fs/B/5fnfbm3buSaRakhLmikgp2Bc1Vzxqw9GGGjH8rdRYnndKrka5qieb23mzMV
A66i6S6Lc2T1IxWoUOpXY+qTEyuHx08EcgtSd2FLsr/lc19jsiDkNiwY8be6rLbX
T20MBujZgMHA8BoQVO0xdqQZdQhD1iyblmpuj1uBOm6uvOqj+0LyFoHnUrM95oww
5tK/ayAxcSfIiVoVABbG3uYoHtx8QuNAtZE27TFPNfO3OqOz4XkERTr+5hvYPDdG
PYJaRFqqXaKreDFR0xej+nZt7dwVrKU1P8n0TOM8cto6I9q8/0dtUyWtWiKVwCcV
6D92vY22PiOTtfB1lJH3CUkZsRWbif5iX3QfROtaSo95vmrKbf8aj5yw3OpMSlWi
5JNy5p1ZvjMphuSFci9hkiV9vghRaFeh1PlpJQY1AxI=
`protect END_PROTECTED
