`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A4aq2eR4q3r4o2+yOFznWtaGCjsxeJHwH73HX2hQQP1cts7XLQBipg4apRc/eCyQ
uFhQype9Eb1uqsR/6c42MwI1sIk2HKJCwwoOQTbHfr4y/xVzGqQOdm3wbQIgyNfA
ta7cBt+rH+GBCL4ro4zZJsg1FQrGAUK4rzUIXftWDRrzWzOe8WgXijExMvKk7dk1
vGgG9/YMd5Iz31lPZkV7Yy6D7Mh4PzzY8k6gDf2fNtCmQ+TRZqvZnkgjlp1dMw0D
hF2P4AvyA8YwKYvIIpsPCFAXch+E7uPxTMyFJ35hbz5WctRlpvjU++cJJ9v7cWUF
1OlbQV6YNkHLQBKei47YhAJHeSjG4w1kcMcfoyq4iuTy8MumXLCh7oiqzC6CKnI4
`protect END_PROTECTED
