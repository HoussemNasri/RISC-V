`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GaVXP4WVl2Sg3j8/H7aF12fPfUlS78WeLjnhXayVgINUqQet3FKtFFEi6AYdh486
dTkLN7s/08dEhUMG2Tm9Y0a/DWUH3MnmD08yxkhXWQzF2fx+KUFqvlZV2pgQB5Qa
upwF2gqz9OpLwZE+BYGCazY+j/UTlw7abe6K9SWTXf2+OfnjS+/mUvHQHVwHda5b
`protect END_PROTECTED
