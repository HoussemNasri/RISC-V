`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjhZIwhPEJETjB9nDENqtkOZKGVm8tKNVddhh+940c1a4mroWj2Su3yz9zP9zDhv
n+wv9difMPnQlIqg2wijfQw2Q9H/sNyAzT+ZxBM0d/S2xq7ndqsCNDaxJ9i0+BF7
M/JnFl2JZ0GSRMYFT9Z/Ge9h84OJBios2oGsGHH3gN7lTCUlkz2EtzxZkZ5cQZt3
4DCPy9nrd26v2oeKpw20NYKtIfnHrDZdj8jx5SPQqlP2HQXwiIhJupg8QqlbyZow
KL6gnzuoo52EwnMt1UpH9jRJRwfKAicDxACmbQtcce8jwA6rhgti2p7msVr7Iku3
liYhLITRpocXbPY3Y/3adC2Kt4KLqwRT0VJjK6iclYGX1pfRY/wgQW0an82t+sJ4
QfpBs8pwBiJMhbYO7WGR5XZfx74tK1/AL7b0YvUdNCrLtRenW/OqwGKSHI0QJkAy
ImBGbomryjRgm3lSyBilTaDsSVN7/37RqpVegfPHIzHsii+RByJzr1UTJ0T50dXY
ImKPe9Xj4b8PjTDq196r5dB5GBh0VBy31LdinLcRYEr4Yy/bfxSw8UCqCYDqgJuD
6UJk2ETrPl+GAsbACzkJaT0nY390SOsWfwiHNSS4h2YTf7Gkj90qbzpAZiIyGYmW
I4dA5M9hTVgxuXIVKKofkk1L4sx5qVaO8RpVxVC3rm4jgCponLleUWtteCfYWdQw
WOag25JldywuamTEQZMJVT/1r1MxLviqMzEw5xFpg4yCP222BY9FnKhgCvb1chaE
F0DyNOEv/DuYt8zopjaViCtm2jKTYqKSBcqY9ZBx7iXQDLQDOL+X/j95nnQH8b38
QYCkzGNSZkzUQ/VZ9dphHPSEpuLkU4kSXLgZ/lpD+I3xu6vsq7VfcpSoZlDWToSe
uQmwOxOwUVcdj3TGrFofIh5rtAYHRk6u/KfHl8+52yyrO3fbdk/kIDXSnekTQ0ao
Xkgb3QI/VZ2gWrz54GYcC3W9pF1R0BFtIVKtdeWJydNncrO6uBN3S9BeRjr/cdpU
svUuEpD2Yqn6Kf1fHVTIqU9kQn0AVGUMLvrT4ZaQ0zqfeYpBbOT90sdLZysirlQr
stFhsIDPSOeUf1/l8KLbKF2sAyLwH1kjljgfzDxzMU7SSuUbWS5VtdzFz9b9WZ9L
JVGWjWb0Ihz70BVgt6mJ4U0ydqKvouyBCIf0NLebjv8GKtA8j7x/9v0IfCfH4ZR0
OaIq8O6g0NgRy2qlfYZj6sDQFO6nwJBANfNoi3+YOBRzmZex9iyZhAvBDb29SdXU
AeeLQTnrkAqfw1j7899na3tD7d1TOiqgmOmN8y4FMaaW+sW4y/iS2+ItaxVEdu7A
3Lmm+oftuA3k4Se8CnES4Ltge+A2WUW4HR3jNZ9TbNtB8VnMvRcr0yTZ41Ouw8Wh
s8NSrdAKqzM/pa1CsdcHttmDPzL+bTcf7HF7zbL4uuQmUDWy47+w4zniqj867IN0
eSKbkyUxByYlmW4I0m9IuCZwFg71A5C4veLjHn47JdAeWEr4Ypm82qpYA1N5XjyO
2Bl6UpgMtrmL0GJHQAGGGGqfwJiwcM7/3+xWn7rmarbLq1vSJjxOIv4Xl7FdeNZr
wN+Z8IJ7mfQshRnij1BTtfYNrdu3wb19ol3W10rEqarb6YopPbL6nWYzVCOv1dGd
NtSTTg7fIEm1G5sW3243aFblMl5r3Tj5amg9ei10YxSrBSD8uQS+F1Qq694pcgER
qcRauPa+DXyrICN+jlP88sutOVMhYw8qpL/dKGdiVeSWzqc6vEAITAhl0Mp8O+AI
ZryetANSPKVj8AgInqeAecX+vFRGnEP092aaXX1sL52bPbPbTBBPx9u75Nr2eGX/
FZBeeDUkcN07GvddrGUpf7FbHQwCvAUF9owYIAX/QdyyCr786eIGSIDTv48y/PTU
Jnrn3GoP3JaCxajShZbehbO46pC1NqXp9U6EIXfoovBqgm4lnZPvmY5bRsqPrlFt
MWvwWF5jmYZfpJt++x4fWkleNXghDrqxgt4sx7CHRKvS12fGJlxZaiUDMjlRM71j
FXk9g+satxpnm+joqtXIvjZzjHGA3NBx2MoIBnKubpIquIoZuhYv2dU1W3aEqanJ
CcOEzUumXbfl2XAv9dM00QQ5c6l1eapEgpitoebaGynNcJsojFfGoayzXiwn+yIE
BjsWMvuDYD4/YMwkqyBx3IQv2uNAIwPsjuZRPBX3TiZZlN9BhDtFYU4/6ktpE/0U
p+q+arto0c46sF7gM0RZ/f2W7Q5zKSM+HPZZGhvxkqpWTVDB33kO5vT3f0rd3xLP
LQLY4TsU1aNDPlzfhoHFrS2cW9fHFgHglaXBCKtHXWer5Ynl+swBiYLoDj6DTUEy
k956/5EDIkO73JlvWB3FLQ0dO5JEuaiH9yq0I6B+wDzGTZIx63oapvrwBhKVYfFF
lk0R3jqbkQJzQpHxLOC/kSK9+1GzfeTapOlhit10V/3FPW629XXOgZmepW2bCYPF
vYZQa5lhlJhCJX0MAiXZMwCWztTdVUWBp3Tg0Mh/YEPqYVWGpPIt/X0AQjixDoDb
nWnQIHNlO2N/XJF2+dSzp1JaPR5Q+o8klTRj+7mwLe39e695xP9dydVLGlqaNI5L
7cmULgkwaHznu63SeXD1Ex0yDvLcqSBoh4pM+ZZNvM2NlcyPaHaQFK2/xGQI55sA
5X/l6RbAeUOIbSDjAGdBTOLS9xUxUGaEcO7QWyYJQ20LYdd9u5ISer1nLAzkLJol
PoX71otWPuOm3s0Nj4EAjLtJ8kV37HkJdBpDFN5tk4145YV2Ir2EqirI4cSucJvo
2mrqyz9Som8G8F8xeQwoO6QAFQa2UAhMwmuzH/CW0lnfw8ttsZtfZnk4Kf/8XCm3
Mv7aN9yYjt+NtOmgwwiml4svEJL+52c6wAbEwVGMA7qsSZZxc5lSzM6uYQwBr1B2
p8YyrELvXZCru5GOhQYCToQDIR2TnnTMz/iGTTH58Emc0Hg+RDcNxYpbKTxoxh/J
huGe631Tlc5D+prpkpBzNY8oov69121eXy1cig0IssPPqR/4E27QDwThOK0onx0a
zdVuwFCGw4DA5zGnsOGGB4pMoV9RWF4ZnW7F24EZwr3WpaxC3MMP5SyMntemjbPl
F2uEOuDMoy9AKPugEc4cfZAUeGM7TYNtV/GPCbeVVyPuyj1guH+Rm/Iw9EOCCX1/
WAut9iOUp9avVDJ0Ksiyqe5w+0vpPqfOyQOj8/HzRoswgWNLPc8vPCtCdGQm8DQj
xsGx/rlIMUXj2clnGDYWEhW8R3bu4Bp2IZvT7I2DL5Ncc/DzlNGGJyMcc5HgQay/
P3MiCXIbGlvEEkf7xM2P08bqfCaqEajCM9KYVAkBroyu3hyKhphaCVb9W+DpWUWe
wQ/R1vN92ihRw+tky/vIgZPx7KBAL8W5Km4pLfUFNOLgZ6MEg5vZlAS4yw5nm7+N
okg9yq7+ZXR1l9Oe3opkjjjn6RufU96zr5FnAOFbKxJItvM+xNGvx/1EfllCAta7
9/K96UI2pEWVaF8yXhg/CzAe1ZLrttqibrLKUzvRLWgkBWaNyVbgWP2QG5+T82j2
aX34oD5uVK+k2WW3AmrUk2VCMO/bWbfBzN6yN0cCmFbQmqV6kBejfry2j0ng5WEC
9WnPlQDzxFdlw+hYk4lc4aZieGHAKn+NEC2F0xo7nrnWqNviwx9dl8XIuOJBYpOx
806j+pw4F9vKmRPlcKh57bYNOgNAN7jVkxqM5DDeKq44Nh10/CWdscmcJ2pvUMwc
eua9X//d7mPuNjb0XJgXLIJq7693QGr88s5XqsrqbKe/OG+dm829mw9WTzGAKBI0
xQq7lASzg7vmNZ0VoGYe+dBidtLJXOsME5xW3o+hZkOXDiAkOJTh3HMKAh6JFgvM
v3Ym90nokNDCCZQjiaq2b+mDDcLDzdHonpgpcG3snlicfIxlcL+ZpWrEliNDZmwf
uX5AK0CSClevSHO2C4nWbrtXBMIt+DfAyENu79yLBgRFaM8ZNqEmWZkM3yrqeeu1
PInyGgmRYLUUDNQo6FEH5A2wdWoP2i4M/8fiIikM1J/YAFRi2cZUeWMPDs92w0Lo
j7nNW3nLL5LaYqyee9zeYLuttaGmrorl+MFiVGKuq68QlikWiEsjT8OQJCAg5Wjm
R3HGAxzEC2esFFHsynOPtObaMYXUS1BxLV+1HTPJLHqqJMl4sdQ3uaYLShBPFQ1f
60XXd/ELp7cy1k9aqsuq1Qr0nJ6zjQQLKEsMVS68KvSAK9hUqNQghn51HFbVOu5N
mP4s1SNiETBtCmPL5rcHlQF886gLQEXiPc5LnnNa4m6P34MYTHZ2Oqm+YTj9kvB3
5OXGILR6lt6Adb+UlOLIWq8P3Piy/D5DE2CUv6xbf2/FmTgZi5fr644c6MzN1Kc6
B6mIU3Y2AKddPUE6FqKzPsyAkUM+Qz//ZufRlZVlxPaKM33JAptpDnZ+OLpMiR7z
OKlcnP09wM3D1teOnZg1cVcszKMHsl4ckBDx/hbwbbm2AQOCdkzzaBTfAXu8RtAH
KS29HzBrez34DONUf3ZnKeFxlTlDKvr4s7OucZsImBZ299hBelJ1dC/PUuVPdsSJ
mdTxAbKynX0s3Qb74h+UGLcy7ItIApyRPRHYh6oE7RU9VdjCWf3NoqEy9nI3UF3b
i0j09BVvDW2bvV7byqlsS/BY3MK06O0LT8Nsi35+WuRcqTTYlo6RnGqaJxJmnwh8
lttvtcOrrYSpS8vxCt2N2zXmpXRsrc1ZklRvFfCGfipfc23/n/3UsZ6e+QCft3Tl
hOMtOB5tmAQX9Q49G8MGzzQnOuUwdWHFkYrBCHGmqbGMPl6VjabC/qnW1T6vzVQx
8WHmoWY6W81e2zPsM+XlxHtK1Qc+jpZakRRLTDvyjtZvQPLB5N+sV6u6MuAc7Wkd
nsU+mi9frBJ2X10cyk83Ge+HUQ7enCg1LCNs0UCp3WDvgI9lPQc+mruBA0eSqQvL
Sw2HKT/0ZRvepeCjzfgpB/5etCPwUX0B8oxdqN/AigcR8RzZGQ7ettwEQGs0HRnT
zGQsf4WxDFFr6G6nXifElkSNqvI+gAK/cJNdC6h2kX664HlNuXh8IiY9anc3yDSe
rZT/i3pyuiI7DRpO+b72ZDEi0KQhM2It/xGPQfjtnpGWP31ee2pDB7yUOW7geT0Q
lEMf7THq7oU1e6SFjIXCi5BwfuxK/2Jht/AdFCH/AldhN3Xyhj0jKi8xDx/8Lql5
MLkDPaFMBP5JcPd7yM0ApFiYV3TXcJFNCMKMtN8zohZf9XCoQmrOWPMH/I3ewD4k
+cuELzL7LYTOP9H9NuKfST6aD3Peya2jBikdTIydZtA4qZeZYuFGcQ60dF1LhZVh
B8TVMEoDR2rMhSnToCVoSANTt0x7Iu7wH5eL5pdNLu9t0GMHzMRvd3U1fPnJ6X9L
u9lwbyaJZh32WIiPNsEiMVakrtuCHlkFGxXItifmTkuQl8xcyr8RKXdRSQgWnVP6
80vKDsnRZ2tkqVVuVeNaAt25XjBN3jVCQQMJwQx9Zn9EEvUmqFOLE3hYCyXwkR/a
jOHexVoz8k1e3pXHoNdj3gEQwkshroWkm4ZQyZc+vX+nuTpkeYtxt+zQd09iC4t8
51g8lE+19cHgl3z4iK9EBvr0kl1sYbfOY4Q9c4rAi4GFxasNmS1eqDjgvcrmh+a8
CT7bAlciEuaUs0nh5T6KaruFQ8rJSpoOGDJrqPPbYY3nmZuHX5Rn47FAs4mAOD2r
RRzkcRHHh3TUjC7R3wLpKGv5bNDlpbryPmc4nmhfrztKpef8fnruaj2kaqSsvpwh
EwEjzJ6WFKUKcPXhP0WF2bR96YX6b/az4YDSOGtFCwhG8bfVMaPkLet5skOoqB1e
ka8hLCsPQ/7SNf/PR5/iXXiBA65RwpFwojyU+zEF9cNznbnvWBaZV/hBXUYa4jgY
A9IuU50jOKdtLI386TQsjzMRY1RPY5Ez7GJelx1xlq0jxK72zQ4u0CP5LmQa9aff
sScCEs94FWIwJzwziEpl1YNQ/5C69gahsOmuhnKevks7Nt2ZKxF0+L4opmPPiCOT
8Nl3zlS0c+C8uL6t8O6E9zDoJ+vFC6zZpWT3DT11Q5yDpA+oAfsSckh3lyZVi8sO
cJwo5pZzZksVH8FF3SALqyi6zoDJwkrSOcHU170hLnBE5+sS7dvr53lqzJsEtK4c
nRN2wnCYJD1fKLNDZO4549cBRml0QaNMT8+OJQdTSi5mafA6yEqcBeEAe4XkVvW+
+ZGHBRrDKD6ad7gNknhNvk7bQr7fHBkRaFbDn7juScaokMvR/8U0TU+1FibWbNEU
Ijr3jj42cNoo2zwQreuFVSmti8+pu5V3MyfTAKIfD/yQr2Vg9j9kxhhWy1Yo+2He
//vE2oZT1rmgd8dOCiO8pf8zjWM/JlxiQfn1zj2LsA5MvR/V41t2+3O9sgja4ERk
cpfbVonUiaVqmfEE5NaLxQ4eOu3op7LKPWpnkgESrEHsG4vD/zM79OQ6+8USa8c5
3lBR/4jPu1ak/lb3LwvWkhYyPuxxK2eqdi/RBPr1niK+ewo7p34Bxksr5Ny0TbBO
rdy2zyWylqGmCoCtKVX1H8l9Xj8Wk2ilRGojETaBNDme8OrP1ULVQh+B5IRBnrjV
Re5UP7KqpnheHTZjlgEAObWcr/Z2+C1ZQmNSo2K/s/IhYSuza9YkbUOddd5hnaHo
RBork4viFmMuF1vifqKpWby/WgnubW20A9uOQGvF/pYgXX4TC6F9mYgqfRazWoC9
kfkBYWEaVNfKTcLKJleFpCpQCwLgojR9pJVWBQERPSeaE0YNNbt1kOpMZg/k4T32
7RhtVu/4a8CnF30dJMH64pGIOHDKRXkiuCfIXCetZKQ3W3SVUTidRLzC/rkbp1Uu
n9gVBjhnQ2YGL862L2+dS3WitzWqnyKVlVJh1xAmQL5fpqvtdtW7+/WmpUgk9PVh
KOo4zftvzssijJG99n43fcj0Km/yMMM9KKTkuGH50oZByFwH0K96RxU9K7v51QbI
+I9fLK2/c22AikFnLMHihgQjwmkUOAA6YmdHuFeILekQuEMpDQ7DzV7KTA9LX/6j
unksqt/dMXSfz/0fG0cqKgbABl8qkDJtm5q6+w6VzE16P4F1Leg8kKiDhKrN6R3r
tQb8Lh4uxY5rdJqj+irNmFUlOzI+4LQR4TrjH19wgPTd2ut8CkTgJmUZ+w/GLmWo
tHH1QcUjVCZRlmLCRSN8x76ejeCj/izv3pi/kdHkPhlEotrBTtNF5bFnjhHkbFJn
Livw0jOfbwkyXfizSasMMg==
`protect END_PROTECTED
