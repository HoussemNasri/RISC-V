`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y78SyK2njO2mbwQbhaY7uByrXlq5wLT0/vTbRsEdFfYcDpMQjYCYXxKhrjzXCJNx
axIH6JmkzMy4szoj7T2/1SResIozDJMWM1Ib8dEjaRpMrHZf5xmhsM0s2VpAM4rm
eLYEYwDUFtB4ZF54iGu5nJ2RD5ybu3t60UDD8Yfh1YXj7kYJ+FG2o8FMKLKOBnrI
h01PYvlxFUdklLd+c2b0K4fIk4qVS/BBGOzVpe2aLpgpQTezZ3H8Ls2SdLnncQjx
Tgb2+I8HUouRYwY//G8GhcviuE1yb22VyKK/SO+Di01qgbUwvTN+tc4yOOFoZGBy
lUymLCd/65bsVkOLmLkc5f94OksUXiuChqjsKWjz/65cw0jTdwrLmjMGObXGUCQj
uXdujGJMWUS3q0stwo7zgRS9oj7GO7aoxjpg7lgRrkuAtAoBhmCex1UheEQHmIUr
ftiimb+x903XoW5TBHn8Ml2MQQdJToM1x2Q4aFTmdngMU3NimYiMXhFvYUE9J7xk
VPnzs4UCANkcRg4YcWSif+zH2YNDzaDVsostdtp0NBoaJRONndzDlOaj735eD7Hy
a1joK+3tLeYsAJyLLB4Azdn3d/iuRmMOjBtFjs0SQbEenW6Hi9BAZOrkPY3rfRwA
Crs+KEUh96GnqZZVdk52nqdeH2UV6MZqVqWRT77r1dyD+NDUCZ2pCpcSIZgz4sgr
RLZoSlclRoVw90BJI1Dw4LSQKBW/S7PLzObKkgOE4aREiDNyc4AW8hQTpO2ct344
kEwDNCl86BiTDCHREZErTurqLT+CvVqwIEyitGVibv9Kf+AdwR8Fww40hYaw9o03
w6SeEn375cILa/Salc7WPVOtqs6Qhi/RdMehO9pqwOdNIpoYAGiWlPEo3nJcsQns
j/o8oqag63CiiCo9qkysCaznIDzxXed/t6WFjFweUjI7qVBFOHIeamhT5l6xaaZE
sLQivAWsWwWvvM5GgVIHAEmZUodH8Ttpx9HkGRrfMunx1dtMA76QbBdkityX7QT8
e8oBJGq8dtGoKUMNsaMiy/PrJmQsNYAvpoNP4/08k9MTwDWoVAgzYBwISTdPj6qW
HhqAFrSv8+/wHjU+GKK9D4HY1JOT+EaIyiwjdUEYbqjdtAflVoMByfY/ZWMUsv7Y
UXryzaRF4JthMs0YL0v40eq/gg0t16ZOcvgwyyvj/IIeq12C13XXW9GGtM1+zyzS
QUZtUB7OKj8v0LX3dLP8+zEZp2zEyKCTdBSmSUX/xFlgSryQuY0RUjEHrA41zDsj
LJAPCTjfGSWlm8mmeOSDgNaF7eYOpVQGOQXVfs2TYX8U4mr4B2WfLBODeNnnsL3t
RX6n4J/C0R6qjTKo57Vx1OzP+Tqq8RLjZenjVpB/e5eJQ9rOWDAjO7GBBVGY8vAN
Ftb+hiDoMsXDcbrORQswZXUHfAdrrgosUD3sTcwJlap91DRVjDQjZ4ZpgroslLoi
G5mFxIFWh7hLY3Fke7bs4cIn3RSvTo3IDJweVERu8LLjVlNTZrS+UFO9LTVwNte4
UVJv1bjkMTSL/9BBRx+T5h6DJfK4ffBGPKDLmZe++OUtRbu1fJzazN0uK3zl+M2J
m1LTl6Dq7YVInuxi9+GBh0FJG/RvUTIXxrHMXdRJ9YkyGhW5uBzncmVIEL392ca4
9LgabxFfiUT3JvmnVW1fRBQ9ZvvmvNmP1/l5cG/f375mZL114aWfwOrT8mwdZQhd
oIyCT9UlMyvzGh2vbZ9e/wgvIBn3eqOa9JwFOy7OjOzHg2WwXigggNOTQesfqTqz
QlWKy3/8Umc89pxXwD3I/UW2MI1xywEpB6eFSE38qEMHLoxnIUXePKB1yc+32sDb
H3tsIutEpO0jBUinqAybSk/wnG9SnMJXXy0KupNHTuZ5I92Ce62j1TFoiHDNf9WB
DzVAHijOoi7M1ktZerNnN5NRbEuhNmZV8dcSW7r1L0U6fgGIh7qvIEM8/TZ9kw+t
CmP8elsj7ddgdBfl5lxP/2ZaXdfjRzRR6/KWmQZJSvmV482igUEHWo1dhWMqQ/ef
mJvK8y5ylgRdS+3ieOeXgYIhRcsgkrTA5GDg/IYTrJwkRdQwxMOh0dh3AcM1U7RD
EHpJGACUELxUm6Tt2gA8L11F/kCGsbvxb0tZVfWGlWZMDcEwK0yIyfdOqm8qaQhK
d7areve6NBBx4YZKpXItl6CbV6IYL3r8jloPReuIq3LOgX3QH84tq+Hmn+GPxnK4
/SoFx4+DPp/sMUJkDMf4kISMt1IuiLPX15cCuzHM0v6/Tvq1RYBvEI9Dq1pS1rsA
XpYx3vex8LaYOERknZz1e42dmWCmIGDKcylSbnwFYT+4wc4PBWATS7HBA0izvAuq
xGfgwU9ZrZ6XVjHnKyS7sGsp6Qt7lYL5+xQ+IQlqcP2Gs+ORG6o0OrUZ8hE4rcxU
raX1xAARIz7kf1WjP0eBeL3iKpdRBapnuXlkpoJbhluNG0O8Oz4IygAdb0pljWqM
WC3qAnhc/gec1ctsaanCkljX+l5NFXtIVECwoGpD+QX2u7mJIkkeVcS2HEynU/m8
WHfflxBAlj6AUW0Kxbg8sfF7V0M+otpxVr0rzuG6ZEipogYTy6ZsQubXVee2uGnv
H4QxPgtSSlOSrcTl3Kr/xogcQPZUh0y+OJLOzqHbJ8Zqm+5ESKZ+Q3+JYx34FH6A
g6kReBDJzyJcrwl33xiSAGWfcLIKo3a0kAlVejZMSwQniKsatFHat8YE8ruz0Ccm
wtS7pSnBzRtBi94VmY+/vt0EFZBfGGPgf6QKf/KE6/vU3KiRDAGVQWH/xAZxaCR6
Isixc1FSueYM2iFsYCz8kEVz1C2ZlAVNK7NnoZFI6xIH5g30hQDwdnBalkMGHzy5
3WERv8MOB4efDBjmv52NF9mBTuIjdUXLEFrynlzAgrSHDJFXKn2+Y+UNSN0jj8q4
DmmZ6JAHUlR13e1CWIIAav9EMIluur6pSrETRa4BJ5WO1G7qBPrz9SMCFvKxpESZ
zufeOEt43imBvyf6OB0deAg+6BePMTyj+u4vtUUObgOo1gMpujEuMu+/VVA/7V18
5TICyOFLhESkO6E1SfmswBipHLDgO3spNidKjgHRED9hF8/vqFpKlIM+TiEXvYWO
8lfeJBDEzupUaClx1m5pWZpfWVbFP05QiERBEMRsYBw0IfiEYh7zTHA87y9XQNZ9
7Usn+N+Fqg8/pwNyUAXx3cmEa0HJLD7ZOsxk4CTQzV/y21aWpmrJJY+79qvLhzVh
sH/54f+gcgG5kzQeGVe7Y7CW23n8+uHu3l4btmdRnFy0tWbNZkPBJ3ZwN/CMIwia
ZHuTrbH4dxWPYjfUHz5coOYVYaLnBD/M1PrVXWzvnrKjXsEQ2DZRwCa2Yqg8N+BJ
Vp+G8YI1/dCPaqb9+j5B3P60VLzFrc/Z45Z7LHgTHIEgYa3REzGBF5bcrGcDoUv1
JtPy4LwRcNAgBj/G8//dFUOJGGu5z/4PXn+DMAo2jKj3YTM8AVHxMRLXPNbzFN80
UuKD677w6rPuU4QfYdt7gyDlDpZrMVxKv5HJZMqLIrBTP5LqszN7hhiKujA3a+W/
dS45Wjc9N1hstga5BbhwbtbwSbyFYdpCWFxtO7ldn9AMQdDJhM6yktmxfIUKTlJf
Ng6tWRvWDP2DnBSWGvvvngZjAt2gdo3HB5F5hG5wM0YVncBERl6ZjrgXiB1VJKOo
JgBbsRY8bg5rUyKoteXBnQ==
`protect END_PROTECTED
