`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6v4XAAloMnibW42raNjExfNRt2mZzgTHmXosBDfU9VDIXUoaPKWOBn+gx5uGZXcd
MrlXwO2ZKdOoLwsRcvvsSWnneVwd4q2lO4u46odZsQyXw57zH/CRUypdUGFZL11z
dSMLBYEl3cxmHIKRIzAkbTZ9WmkNbH2Uagva/NmAUEjYt38zo6BKhxCs9HdWABjs
kvdrXA5h5/P642C7927noCDv/PinSYDFc+rrfm9DLxendVuOsrLH1lqIYv8cKax5
Cv6Z8n/4PRnkmWXkh8dKNMZ87rTeT71mMhC0rOtL59AhQp+pKRsxPvwPv/VErUqe
DKhnnvM4hPiMhrEDaCjszU1YQ3pKw+wCPNI1MRvaLdKBvWjRB3oE7i5C85UfBEhD
i/3Y5a3F21VAA3tKG1Sz/157T8oeXPKohcFd2j9hFEhUqmecYfuSswSF9HSmDJnZ
Ge/QG8uGj6r2ytl311qj2Q2a0CC0P0tfQYe9IQaSyV8C49wkLquHjaPxiLalyrZY
rMky+W5XfaPBVBD300zcXTJfto17NqFRlHgwFw9TeDI9yP6bSqLDyhvhToSBvZ5d
dT4BPFol3gc1qh2T+S+DU0sx6U/gJe0hL8WA+px+nyThI2JUZLDsjdNQ+1P5rkKE
T9CNrznij9gmuwCu2eQQ6UlfKZOzuHdXRXWfLhR0lkrEIgIVv+2FBB8ZxsnWp7UZ
7RHcU4rc09t1LDIrwhegQoHYlewO6NSOvzAw8OR2H3BCgJ4Mzluq3QZugCYogMZP
tod/mvhLnalZlHCzYATAYlc4dnRm4SPP+AHEIvUGv5rchjXtK4U6ycrDvr8vvExv
aSURwBs9gHB+cfjus0lSdWEd9X40xNz53ybRWf6bXUt6yB9n7sSEhtpss9rT816J
tD3Epron6tdFPqxyFQvz8A2ynwhlDO87ajK05sq9Bm3jQxzVeowQP4xbMFJIPNp+
HvlEd83T0LBlvFGuH9LuhK52ygsSl2VLvuDsFWOQke1wkP0CaW6V9xhrARl0V4Ak
Etimuu+tLMYzb1ZDkoO0/ypGeqlqMRSgqdvvLMQtR+Pnu/VrRc9FJ/QcHYR7J9rT
paDhBQ5YGEgst/XljzaCuupaDJSvIu9UmxZjZpHO3DkjVA5oDlMk2kAJ68UAdRhp
KM96tZmBUecYDCCLF2nFqczj6HTR6XZmvHS/rUD46sORdeJ+OxMatanUDUpDgbci
pvtO9l+om8+ycx2L4COCU/XSrHdaMel5AkHLk51yMRAWnp9vqTqg11nxGLyZYU6Y
/2jTOGaWWw/W58YbL1L3uWTXja797LsJvuObuRkfuM9xsvKSRls6uIUnX/5vOGGg
YTFTBG9t4TTWxymRe4jukxFQcOwLTpZojziD80isArevh9PpGeYUB0RPMsTJ9SPR
YF48APVf9dMpb1L9ac0isDy/UPX551X41qvgJO76MrKvRVIqusG76+MH/H80CGNR
`protect END_PROTECTED
