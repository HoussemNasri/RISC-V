`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vbayJCdPXwrLYrmShCRqX0JvJZv3di6E0whiPCO8m6qwnkpfiwVkTFmwsTuwc5YC
h+TgUsnyFaXFptxtH/dOKnKjPANSAKFFEx8NiGEItPzYVXimy4MWlFPLh9YTrA3q
2jgWpTQIVVLjKK+csMiSio7CqcjjH65J+GkNEc3qoZTDVv/H3DQUSr2jXG3orHQc
GXHG+2P73JSgkX5y6HuXLFe2FzsHsBatkMQIebTXbL0f66FxfqR521nFBNH8rTwj
SBpq2RML/ykpbrbcqTDJwp1yqQj7RBKnAYmWHEUMpO/FTerXdluWEH3qkmYe63J+
JQy09eLkuXt0hU+Wbse6woZ5lRlllQH5KQSwIviyDJpyJDgVZa18OSUyR+rF4vMO
hkJZK5Wnpwu+u3AAFwG981h3g75vsau5u8qR59RBjSSG3sM2hk+WSbUAyz76VQCD
BXdjYw6KVS92dwmSh3Z2ruBN9Vs1pr/dmPkjOvuboVGZVlytjYpGl6CgPttO5Y/g
mKk4K2H6+eo+4nTFXwNGrWhFeWVjiPCml1EKu1gdenBglk4Yrp90KuoSvhpgI06p
URfahsNL7f0VJqBvsiHkzvdbmg+S07sploUTPW5su/vG4oNTshRuy7LGPwFNY0ww
H1IsEYPiWpjDBinP5jGYiYXVm73hWBJtGUr2rO9CUM2EKvDE9Jtvry/6kS7264PN
EGvwhN9myp+B8ikNVRFZ1l2AU7pkStThNP6CdDnNGv+WZAz4TRCf3P+/9sfPACPi
2pbwExzwNwiVAXwCOc7K5z6KXezAmTNLeVrbjTfy1pxaX9xrwq3RDIiE0SyppSI4
8UB/74DAZIoYak5YMaBcT+7Blhip9Yv73TEfljDT4b5S9kuILVaooW/o+YgsHm6V
4P/AtSZ3XcatZm/A+SEkbdOsSHy15P1pKgNzeD4jDQEUZ+ejBd936PIYdN2rG+RA
j8FWliXl3V3fwBDjEHh32f7aGMHGkX65HV6VHiQVTIhBHWNsL1qrlwcdCtQV48m2
Fmmdsa0CW4dKM5VZii+XjrfPB9XohImphBatYBrMrp2BzawRWYH+4kWnCOHNhADW
ijuaAxmS58BCwW3hvQlRbLmh4YWNP/zz+EVNJbCmjUgV2FmRId+PeazWszIavcfM
jtj44sS2CfAlLDfKPAS8EShHJuF6DdOsd6b0MuXKJUyEGuQOgzZ//igUBG93nKTV
UXBeH/Tgh0YNImrgb3GUSaocu0JCbzC7yL6nHWShvhltQAi+JdYj06ZaQxt7BQgL
IsylhWw0OPHZ11t5T+Hz5x6thtN9PsV6J7XzI5sKUSADtRladsC2VpvcdTptqYjk
4ahusfGim/eIhU7JeNDX4Ne3cKzG08d3zsb+FP8zr2+gzF/SUcQK1oeIVWPbcnL7
dtvFMq5Ns/criUs1Ol7LuqR2682VrUeHPNiF598YHoDkePraR1gfJmRQ/6Zqeyo3
v74hgkUarRSRQqV1UCpbD/kluooc4ka0okHFOVv9LB/s169id3jPaWfowoRZLxFN
CMUAwZGAEQ0rHR6KJt5KviEIr8f4QAynzU8jhnEVIdeNe3IqVK2aItbafVHZEAbw
PdhTsKWYtN6rRXp8KrHo9vxXNAYpg1sSHU8Pn7xxvoYR+lQ0b06R6ydhgnCTbxHP
zrldiuZS+N2Ck4DeYS6dtLSONl1+JOKWfKFEPQ+HlGi0gsBcRdolmRWJr0Gi58Ds
g2ctdtlY3nRt1QDpKZm1z9xddrQbE1L2hXvBbyh08dhTpGKlcCUE7ZZHyh0gmgMy
aItP1OUaPgeFVt+bKgxycg==
`protect END_PROTECTED
