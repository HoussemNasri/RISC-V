`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4tNgwUgroVzI8grzVlHcQL6ZB0/4B8L39Tx53pugzxjPUdLPgl5yEwCjuqjV8byx
A3z8VBvqv5R0I30v3dufaiAIatmS3eMjhkfn+UuS0Ndjh46v0YfMdxqSeEvLR2UW
/tWRJ7b7FcuLf/5oVMVmH0oR7pl3uHOK7MLU0oaeI4mxOrQ7EgJR+fjnv7hh9It1
lyU3yTvtCbiLNfH9996l58vrqD9+AWhLP7M8kLVftznnxIOldh4iMG1mRuifMzTY
9RvFTFgZxkN/zObyJFYySlcNGS0K00MEu+MA9WMMCRdX5fOYGdLfREdTCSiSeVM2
61QNc/e0c5i6jH3NgveLk+PsA+qBS7ZZI300KgsGL2MSSkGmWnrT30+3Qo7094RI
K3JS+OXQfcgYVzg17TvqinsNhjJoJGX0m+C8KesKeBgwGYqtXiO8zIEsRvsVTGXN
rzJwDbhQk7LDc9DTInw8i7U4CENdGdo4pe3L2sr++7lvbMfOeBhpisp/EdTQ8aQ/
9yWB15onWSyiZsf8aMKHt3xGkfogGKPrE9/JOmBubPgrGmMWMv2eV30ss+yMOAZi
GQDONfEa6TvE5o6LJF6RC/xnmfLM9a0jSiF10XZ2pUiAcjlFeBTm79s7gvU5WKcM
HwS4S0ZQNvz9WOLiATgjk304cYeLfg8Oqbqh3pUu/pLOejNnRPW8bXvNSq4Avwe3
uAM2CRuK5U16Ix+6+WOEFO8mKm3d5I/Q0UgAjAg+j2H14TM0Uit46VYhHWbyeB6x
m6UrNwtwRLxLZyPWFg64o+xv34Xo2eeE6xzi5pSA7rhQpA4RP3Sg3jMisyFdBY+O
VjWyVUUJ69UF30mdltcsV4CmuBh5t39JR1SgAx09l0feCMijy8bVqeLyqZzCF+Rz
NuaLkTWtSFEsj/l0fTBXkRXdpwuzy2s1WlOEUJXKFzQqRkppUVQFwRA7Zb48eey8
wDwL/RrNWPLpQF8HLF+yeMg1XFU96hCgrqmLMfQfK5xszWq1wqyhvkvOKzI6GEim
m/nDpCEmZDxbgHMI7g4QqW4v6vCtzPWIdPYu1gj59jfv7JpW/oEo27AR1FDenF9w
bwD2rRUhlIILAI/KjfolSjsoMH2lEdTR50YEW0TFEjR4Z3Df0dCkOoouupnOp/FY
RNXczcHqIoUxUrblDkuo8O6ZEoV1PjJb61a26I53ZcSaX9mptCa2kUJlZWbvBFjf
Rxixv3G2t5Sr8cnmUkhjwM6fVhKr1WlGw9JJ3PNFHvCgK0mbMSWaW2XQje5dB5/c
InrJP116x9pvgpeXUgcZx4TJli/MgRlk9HvCq24DJ7cpbIYuhrk/zhvfWelgle8P
bSQB3cQEb8hIJcT6vq09HQheb7VPmNZXXyqg9wKmAwo18xGE3WYiR+lmEvZOZ8OC
+7heE0vf4IzihInFbY/+m9AXDsBqbv9+e+58nBlGP55l/vtlLIcIKh85cJJ8MQT5
GPb7inpJEBEEpKTi7BmAyvjbEharDxOFBMD7t17lLBKSswg6DuVnFKCk+D2D8Gtv
nnMK7VA3iQLDtcaeyX6sB17S3FiBCdTwe6UN8+MnbHy5wRu9nqkQ/obZu/3PdBY5
CTq6Jq4/KqNQfeg0hMbDNuVYsizBl269ici+x75H4PKSeSeqKxszhH35AvH7R9DN
K63pGUyZDD0/8eV4KCTPRy9+2A7n2QZaTTz6GU246t/9X6L7OyYuO8gsJXUeaKEl
bohTPgVi6v7R68m9fKY9OFHMUFL3rEY5/hNXapWvE3QHvbWSYEbnRzeNf9T2QryY
Ws7mbScnTTI08TDOMxke6HXvmnYd6OQzrnGm4qgGROdJbC4FvfiiZNohDQsg+Xpg
4+cS1MVqhlX+Aw2qmmcOQX/Kzq8Wa+qdcPGDVgAtG91+wnK4lMVwNdv95d+RBde+
HH3aOUqey4m4a4jqVoxv3J2i5ZmTwroHRL2qKdt9n2Aw03jfLjnjyNfy4AKx72ry
3MypuOuKUOzyYJ5S0lQ2gW2RknqBqLLCZmlaFSAT188HA/KkP7+PP3Uj5mb1LqLf
DqMJtS8v7tRWX8zTEnL7lwxL1CWs5KjJYmdDlvp+PdF5zOt+kRGiSltz1qabNU1I
0N1BiQpTX8vzUmfJfmEboM1xVHOvY4/bum7b6BHlb25HJxXpRSXTJjrTFjxRvWWz
NT8v1uQlN46tz484gm3N4tv3SZM/XAP2iupvc39amHmHklQSzy3z4n3QNUfDSwpR
ijPvfcj1UCP0+yi8pIJ/7TBs5yhmN75gDfrD1EOApsr4Zi6/uEPUPbnGSPXylMEu
WdrIKl1Tr3LIjGXQXPNAap3alTcbzHSmtzNfAnXhs4l+ad+Vzfd8nwlx9uTd9nz7
a61hJ5gphTfYqEBvzq+rNaGVZlgSA7IZ27hWsBvsZ6UgV2pNkhsz962GCG4OAP7R
OfeF01HiBTROM2sI2HRgJ7Dem05MyGvioO9vD7mUZbu2eqKVtZkzxEAPQXtpghy2
BrU81ICboES/TKnNLI6Iiu4zlK9bNPMx0AftZznXjzMS+lahLJ5TS/isL6cQGz/g
dz5QnGD39iMUi6ZSMW3ste46HmdSzp2BolYAEfPUECXU/3qgqwJMggIqASnb0EFr
/qMy3d70Bmg/e53Al6vmywnR5JVjchyxTUs1w1KdI0+Cthuoio7BZZ4XmLGHtTs8
270131vdiANGpQqXIHM2PcPxphKA5JLRSyESqZpOulveX184XHrRsSEFEkdNs4sG
8zlPUw218ALKsxCcFq+mycc2HOYf5Tuc9k0qt7CBJlXXIvG0CB0+i3WvSfmR6JqV
1SElGXyN7z8DqFNqPdhUgPrS/NEwOLgNTVDhJJsZRGiWoDL3eSWZroS9Yoqsfbsp
SjqYkVXsLe2aHKSC/0vnrPebxkWiVW2lkpdi+4MVssZYJ201nIbetCJUhDhW+MnJ
U22AUU7sAt+MJQH8kh9v1InXfG+ch4P1azizcD45UKZEYrccu0LvF9ftlld8I1oi
qnyMQ4Q/5wsVftMhZiO0uZxco0nMJQG7tNImrtHbpAXA1hlDUL5gi94MqKdXZQk1
AFBv9B7ofAoPrSdshCmvTqYGKPgKuYQWYLJ48jwJ2WPRhFVJ3sfE2TVue0vUbjYg
H6NEYNeAQchIx2cLNTPyPbCD/4sIqGWuT4R2/8bH13Y23ccxEAL7EeX2X3KFNmT1
Lt2+tXtCCm9NuxT/ADOpToRYWiLlYScZSz6vnhD/+IDRU0NTquflaX83rhnVMCaT
Cl/YiIWqodB7qa5jue059BBRQ1odLv5KmRxASUiFUXryf/FsvZ9P4DpyZE3XF396
QKDAbyXKQAZg6B6vsJip938SMnxuyoceAyAs29y7zTISAmZ35Apidv7nzduuD7k6
+wG+FNkwH+dpsCHA8Z3gQb0WIbVXVg1UGIxBNNJ36e8UEm0QlyBmpEAi3zUDeisr
rlaLgktIbth1i5Frldl6tBSfRi3ar5YoWEjUT3Spqlt6BPxvDuKPS4ALOIr510b5
+OKNUNZBA2PxSyBZWpTuRcKMT7IZbpLurh8aEmJQxAJZvLUjkwXQJXxmL8OAy9Im
jRgjMApYwZ+UXPNyjiS8c9Gd17SE3DTv+T5KVUGhZBV4fYckZFmW0+hi3P4/OX2z
JgxZW7lT4i1ibqT3gnq4IOA3LdDTJhKf62wuysziaO4A52Q2iuxUjGVub0Y2l5/a
fUn47nYLnNU79FYTKtQtAoUZBitf/UoYlFVLTaJA4d3CpaS7qCbX6rsI81JW4P8r
nIjINn9UD1M3wVVKXO/TvFm8JiuQoPCTle42RWj4xYLKYX5BEnOMAo2W9V9DT49z
WufA8+VuTHtYK5Pu+2lrQqbLrfVoN7AjpPt3aOJ1Y9Q+dFEgoKZvrBUfw2sk6OOv
nn1Hn4EAxOsOMaOHDQYKrJVl6VLyKoB2WlaIlOQR+x66Rt+eLpfH1xGj2WNzuD4w
PhOU5ADZxP44jo9EBRBD3Vdeg/yD4ARA8bOGZJzuaJWF+bUctDmHm+MHyUhaB52s
qXasYEOzxWg49imvReZR62clHWTvbJ0R9TyK09Q/mA8vOXrp4pZr3QIvMKlFmDei
IFSsLBQ5sPxEAqSB1X9RkF4UhnnvQmz52Ij9whRVkeRKppGg3ANmI36i6KVbRzFm
htbb/7Sy/3VdJxjn2XXxSkhSFLrIhidx6pJtxG960UC0wZ6VRkgotIxJ4NEmzB0q
q7civR2acfTRW9acm6snZXck7SgAsModIGsmiATK+m0TqUZB/5dWnL8+uvb/8aZ0
YNkNrEv/HUnW6BazxbuwXJ95hXh2eZdCIDAMCNn1wt86vmKvYR+TeeKNREep6U7g
qKryPy2a9Nw98w3rUFvyzT5wWW08YXgnJhSccB8JkbiFQ0T8DVSdSqCh5fYz5R6Q
vNLtHzKbHVIx4TD1JL/SXXgAPshpujh4fax5d2mR1RrwiqeRgaSUgUHKS+g3TFlH
eYktLL7r2DL36IAlpjt79QVFNKRh5QCeY6ZMgL51L4Eq9NhCwjcAHzc/PUSpkGb3
Fs0JL/1XaZ3yrEwn/c303YTHL9vxC1IFeAnBfq16ZsrXCaKqUM6iPWV9WPA3wy9E
ZERJdufjp1n7T8lsiwtGaungZO0LY/MLiW/4MSuxsNvH/dBbrHAaoUvvu573NKxh
sLl51c9SOCYNVpXyy7lCoP3SFLVq5i8ZRGk9bPuEwaMPkDzZrwVt+uJVit5mRHI2
wkPXpJbQNdc/147ocWQTkU2f367ipUZ39MswWyWyMvgihysHVzRezNtZW2pCmpsZ
hu67QktnhnoH+PoVocGyk33OnCb+Nb3RlDZ1lRvKrV6jWNx1vskuIoiwYJ5TF7jA
OLzr4UTL4VEhke67ZsQ+vNZdCmJCw77wrB6kCsRVXp5OP2MstDdhX1i5k1l1J1pG
4yfRi0nyQUwE5hPfz1xJCFsfyZoBRlQ6iFb6NDitV+bHdoJ26WTVJvx7mGaYI7Jn
08CxfifPpzPswcDVGKQE+TLwy1xePC51LCpkGVyBtSx0vr8r6Ej95o1H2HEw6Szt
RQcjIWEKCuXKx1NcY/E5l7Anb2XMLShJa7sk7rW476DpCGOMF7zK7xs0quN84TYx
8ZjEx3YODGyQ/HR4JlwpwM513Y/za+iqSmDARcGep9McfGK4FTsPyTEDUq5IXFd3
o33rlrn93vL8cF51bfMDqwCRWdojnzaKHoz6rUrBxancVu8mAHS22zzEA9v264NV
pWbPmVyGw1r54GEaU3mJ+9vsLzEUxL/PaaQ+3nE1F3MN2o+dk9DJfzxoV0vMGVfZ
vXlkVxJlTIVA/+pgkoUOXt19fkswx5en4lVXDgM25CUYOTbVmCXcrRQI40LT+gcb
qdRe+9Io4AbFV6rA0u+oZzxDT0TRZe57Y+PE6D/kQOo9/WCzHwITZQHhlzpvQTMD
7qc7CbAFbqvlvZP8HMFU3I8EmFH+qtGLZxbJSi2cy15d9E01nk1ms5b7DQLXRG69
mWeb9to1SXrS6PrkC97CVUvpf9Wcik1GJgHXZd8S8SPOp6cTORjtPAYNMG2U1znY
pE9DgLR1LvbgHjmR6TXiXoDUsRQkc/Gwbzh+tOZJVQG/u8GIAlUPXlgiHi2eDvEm
Giyr/lv0QOmPPdL3GqkNJS0JwoH12F1y9G4mUR7+BT4e/8T/TKkZYmuGJOzUgtZJ
q42ddR5NC/0kNZ+0MYlf9/bKbdCInC7MllpQf1kMeteF1TFhUSnswgSdpm8MEe9/
th3iD2rb4wGqh8x9+V4sy0Lwh+MZQh94+dV0QphPGYCWLgI8SuxMcn7K3oSEXeDu
qgVC2GpdIAAZqbALA3kivDseB9I3N6tYDwrBr0a3J5lmXWj3F3ZLuWkM9R4u+16M
GWNW4necqRJM+y07AadtoXfs8+FdxCpqU3Sq9JbatXLMaC5YiXYbet6SQLzwdpad
rU6QoFw6DAjShnj96dCL1ezhnBl43ChvCdjyDs72pqrKBj3uZygBkChRYCBho7AL
wmiZGB8cWxGnuuX1wGIUcVG21Rvk3+8t4RIjfONmaoXkGKM8IhrINgZhIu452cHQ
r8K4ySgTPWqamAp9jv9QFHQs0lgB+xizxFhEkv8ArYOLU+vqPtqD7fZn9szN6czP
UY7J8MsP4EpbWCZE0t3igVmNchGHkn0duyCueZdxGNmkWPpt3/+fZWXfS5FoXdib
iXnNAmvpqQOhd2AALxPzlgPYji2Dog/4QtkjZ3OCuWtNGjwlCNlgle0SKHA22yG7
baTs2O96zcAmyKIChNZAf5/ubN9YumpY5s0vvEeTXVHQjTNgTEVCktkcQ4UKoRfj
754+GJYA/OOFlEmHZzFuuo10ZgciI2XcelaQyShKp2W78m/EtYYXyROhP0PKQ4GS
jhFY8RxNC1j1H6fOxUz+908NEOZAbALVpW29nBDmCl8fMCcK2tR26d8b/7qt5yoV
/4mOX7nZlyHyYFfSxau73R5Id7DFySqM4tQsf9VN+ZDjwp8vgsJUoBPquGEHMxU/
1K+XZfS1M0n7Glndg164KR8xi+kDqBAV+lAWrhr/Tyl4+mztDK4eUE3CbAyBbVMJ
Bn9QuU13qmHcqugI2UZlPjb5/rVItxBk3XoTNYEfmvWs0UmBrr6nACb0wmKll/sb
xz3eUJoNskNRcWrVxT6epHvqeLktdYnJLkP4+3++GIPsH+48ZmGQzsOnEgzB2dLL
LjkvhX4p6xOrUnleDmSLhmTI5P0NBPjymtGTaAaRMCf40ewH3OQCiQTI9mFMIpLk
tbzxSbkillTgDr026t3RSxF0JPyg3UsEKebExGbvMsKAnwkrI+W8geLqP89vf7z9
jo0c9LYSNjznA3UMnn9uiXqszxVx/XTNArxq+FrIUS6O9oOYLDkAQVvR7plq9yzL
hASvKllfa9FdIzu549YBz6w0OP6gmE5bTZm0JSgqzr6z1NbUkHtmFInUbKQf65c9
A3/KejNG9SehVP35miz+6Z7goSt5DstDXZQY7V/GC8r504v16lHOkMIoyDUes31D
vVC+ydaRr3KwpHXjosNnFbLqDo2IWp0X3mBlJcGBX4eDnMzA/k6GtCWPIgsG3hxS
J1Ms7/ll62LlHH1IXqdomL76A2N1Gx4MduHDlh5baM9Sr0xdyKvwBaWJ7yiDl1Gj
S1lkzsehImIzwpERpbPTiwZib10lIe/JH+cRyLTm891MSuL/7RbisejthIAlY/PB
XrAPMiksNZKR6ITKdXPutRupuYrsekroqhWGX0klJpyY4LYVOZuHQP1ZpOBzajgp
V1mPhHkVfwKcsAmisTkUOp3pWjUg1B0eAhFOThGLSjYdieRxXpN1JyMddjx5oVD+
Ogahh+DUyanyu3m1XaUY1tsq88lg57fqlM4oXW4IrmTIaURaHbZdlBS6T2kAVgta
Km1HjPt4FM94y92iHhHMrAVy+dkr3MhC9tkvAdS4eURGgO7LsnJ48E1wpWVmZDA/
G7njJGl/z1v0qvGJP2Wy2joZxZixPUtHqrDBVBGjVtNelIwgxjF9/XRqhS3RUPi7
aP/9p9/HmCwDVY7zp23nblyx4p5QyrvU8dbEQXwDXpzce6Gk8cktHgHBqRFhk773
Q25UWC2fHFoHGaXOLyFxIfdwpybCssC9ry7My5H2DngfhnrgQlms88uCh4OJMvIo
YB+F9LTYbvZTSkHyW1CmFutY39nA0lJq3taPumWgHVySqty/ZsXYJDLtiv3/9cWa
NvUlOkSnq5TZkxqTfByojv3tCmhnebIxmO67ynm9YHwarz+Z+riaxlH/3ehhIqOv
fINYfIfjGt2FRqWKxYyNCJJR4pEy4kbZ4BKkXj6b8p9Bms2NUBT2ar+bTUdv6CqY
BJT0vCb8pL8r0Al42k6XUoBtTt0ip9MHcZtasV2zVED2P/Xks0Zz8rxP5KRK3XA2
RHKvkAMg9MSol+qB39fsXMcSLyoh8nsnVMWRVz7G90IGQJ/QTAfP7yvmXzr1sEjB
QAwhojqUi28QnXdva8/WFgRwB2hcxJoVqjm1cQraCVeuuvqAU6PkOPPzo1N4Bh6/
hq0t4sCiU4qGng/zIaxAJlfaLQ4PX7voyvu+7l7pnQXQNvzar3nmosaM0ouhLP+g
mJ41MUaw4qukE+ZrVRnKgvthzjaeEPyyT2uHIwuuampzl9qqe9UF02HsvbHcj1dX
LKBhw+KJyj0ur18dPgNKMUa7BefCNp2QoXzbGX9aA2Nx5V24S8gIcr1kXUdF3dH1
58Hdu799UN5Eqf4gvGF9E8Yp4fPJjmYYRZwZDdPN9xr27ADgXdmBlevX8pxxe3Yh
nrl8MCukLX6G8h/mk9jNA9u1dpIHjcxitKJjMVyGZaXJjaxSvTvrW+FVgHny7aOC
lx0wkQgPWZxFi2wEKg3gpyBvTfv+1fNSMaHf9sCdBesQiUvKZRCtxjXg6hutMtMX
k67osS/omT5lRhIzRoU9eJ8p5iMhkJKoz/m99JQhypf5Uc0ySm4yx1BQZpBI42lr
uJnw3z6FYm5vNRl7PDfE+bD7SXjSxmmMSOivfx/mCcNDSCJFb3IhFo1POFh1F2/H
c/CLQu4vCDJ8u+nhjMk6Zszm00jZHfxTJORrIlgAQbMnwFACNBpX0o0EqHug7DVx
jeO5cHPL+M7xclJoMfxGEwnfw1X2FShRh15YFWCAgOevE1zomhoW/BDeSVZLWvkV
UTxEUJH6V1oR+aTvB3envugQfmTGcSFx4MtACRpxCyyc67iLIEhX9j86mbGn6zEx
HS0z/uATNJXpnHjEwAhY1oaTHpn+fyRaEaTgP8ufc68lqc1V3sW8Mberskmxt9g7
4+Y/aMEagvMmYbTtvsnmDg+3CJg6Wu5CUj6+IC1srhgHBB7DKxbhCqQVElBiRN+b
np7izKRZJr/2wG41qS+yFMYl+XMCsFIAcwTvJ6FqfKipfGeRJYvGXQx7zPofKEBH
/y4/HXZ4h2i8VNEOW3SK4AfCPLTmbgRr9iyGXNK45Zc/GkImaFI4qmpGyhK5E1bo
EhjDG7fpAIilHWzHEDlYnN7OHGXfuMlScvItDwkQhC2GAkwq7X44Hh7DrVm5YTpL
SbSRcKWIYj+xu+pjevEVrQAcDnhx7uhkRdd9pNm6Sp6nzh0P4DR9IZH+kl/m/7Hc
VzAgZPWtlP1ytPuGymctSm68LxLSzBoXnhZdqU4XRikAca9pJoxecT4uXN9GXKmY
PUApk3vwWuP9sVyGaBWMUsPejM3UGo8TEcmf677jCwzNZwInwtgC0XJb+zW+CgUq
dUTuxzLqKrt+JTeZx0ifp5wb1A68ShORjkFWIckGrMtXogcGw81h1srFg4v0BOm6
ERlW9LHOwON0NHEKiGG+m5huCqdPiqrlZ9GvaAjMr+Qds/YvxBtGbd0aRjtEqPfs
5wqXR4anW4bzDnOv38O6EMw6Nur3jzEhsSO06sh32fCkNO/kobAJ4pslIUiOFpxL
NrWzATt/nkL6cUuXAyZnsTrft1HEZ8DCOMf+sF5qipw0P7krykWJM48NGPouBjRq
iuP+ad5HTdvg+BusXGKMywlKWnaFu1Bur8sIsZATt0cOcjPMrthiBvNzPx0Fsq7a
cz6L4L/mwd8fg2oMemJdx8kD0NeFXVlLPSuSvcGbjLU8tU1r9CMyuP2zOjTSuAzz
tXEc/s6XVtrbVl/n/L7ItVmJAw67DYY5Bfb7rckaM/JA78VBmUwFd6D+koWgfvtl
cbI0CurFvjUQbONTgu2gcOjU+T28NY00bui/5YdC2py/wmqSnH/wrcRu3SDOOrf7
QI8v2NMUDYfnAPiq5r205oXhbZybfUpabvWv1t1A6wI6oqjaiOHef3J5cYwIxpUK
rReQtWlFlG/bZDKhxRslLEweIAiOqK/vMF9vORtdABrTIjxfcoGFnQgYixVXPZ/g
3Z3+IIHleQpIgTTxqFda+ZWQXQuwkf2rj99TKQnUsqcU+3iUFGhdkiPRjmzD1RU4
sqPmnsQkdGaazFa5jS5Jfj4cFASJfIt32ERxLVvkaEdAAOaJwIz+gGBiiGFkK97U
wETJssHzWEE4xO8MgEjk5qF5Hku36kTdqUszaHUBp8xf/ZYK7lwHC0PhsoPUDHd3
GBF1gbf+32zFLZsJy7Ly2y7ymj/R7hnQUJS7cnv+ac7n9DabcarmphpvfFy6UBMZ
P2kTPnBjOiynNRgvTTj76IzN6+LaO+3PQpseO4GHKsjLRVltzT64jL4F6lrj8IXz
e4rK69CpCJgKQXakYRVRpcG8ZF3LF7PgsCxqyixEmNzlZjVLWqge1mPXTZ4JZemW
8v5GL7xBCSMCVUgIMgv9Hr0SB40+Wu6tsy2WHtze9YMzphv3jEhGyE4wtqmdK0bK
7ITPRZFhkWgSZ8pUeR7wRLR/ARhb2NjA96Auwv3bcfaIxD/nHlnOwuS96UiqEjLo
OAcXBVCaTFdw0NxvnhN1ryGt/4MuAw3+EQU0muFXey0XOZNIBJyN2pOntFfhZ7xh
tGXwLwbHpxA+j3El0GGMSmOAt1AZ3P4xb7+ZeWisUeMrrj439/8l5IUAqX3rMbp/
4JzlLV//Y4rEx4s/SRw/T1LF6YoxCCap0jyiaNxXTXNW/gkQav12Wt5/aqEaIh1y
gp5mI1wxSUje8+bWCLuD4xuOn03VIlkQrGG/JpuJA4LByFmgBZo0kFrmrmq63xXW
1gtT+EehZCXMum9j5RfmifOKRHDFsgVaVr+cu2GS2rR8zIxL+Ywa9xnSX5j7VQtV
MzaR9dC6s67bp1Lxpfm0igEKDshOCcWfQRwrUTcoYCs0tRaLQlMa6MEV+//ofeCd
8AKmDUBbJK9vlifzG9xjI3G1SzHX6BLFmc4IYHFYlR/Vt7Hcjf4fzZXZeneG7W0J
lnSeQ/QHwIbPqpkffeT3cmnQF3o3lAv9KWXiRQ349qIbnCZ6z1FYKZ0P3kPrum+R
5FXYTE+d5PClVqoEYTC2SXYdObypgMKGO+enAwOeV8MFl+PxQeDWR721hh2a60uJ
XhNv3c7MLCWaCsqGbfiVp1+OBPGT3nMiqVFKmWzi5qfjSNvWkK8IejD5KJi1d3cV
Je63a18NfqGD0b2AdM+7F7+AYmhPMMPAA0DarXPck10jufjKV+nBeGh4XhdENB2O
qMKvEzCZGHVizfg5woXHP6fMQNEbk6ful6ELBf07jLH31y7bFwo3zts8BLKb2NWi
6lDv1kBEe2yjoFLZBUSHxNhABMyflS55WqsazmcoSzqVT3coLCOaTTB1OqnB2bNb
PUpcQ9KspXw+P2V/EYAssKMs+jI+YkXDG874bw2/gKId+z1h4xqO3g5KTN8xFI4W
Nt0XEjj3nwrXnZCJMFJmbYmbvrQXiA47es3wJYpP1hD7/Xmq6sCQ3gvUR4h0ulOs
+pu8X903jwWOdXypNMxRxF4jNTr+9wMeSYNZVeLtVfBx03fQmG0xvzcAj2Dj13uW
xz8TxsVYGMNrpq8SVoKM3Bvmufx6Oa/NDbotPxcFrwm/HUNKpyW+5XjeJApdrNBD
SzLjGPSzk89eWwHrNdwPbeEg1U3EaOZFTTmv+7M7BaZ3URoaa23fF7jXVwV01y39
bfmnGub+2K83QbFUYOjbCVZjUXUt5D/JJFSIfHhJ88Eo1xECTuTQDYm5py9bPSat
6Cj9SxSXO32oN5ej638i+TGf6zTGl0Dt0SijY0CpwFAodKDSx+RZUTSo76tVK77M
uuYNA8qqxZYOhiZHMqUoFL0zpX/ZBRzkuyi79JoWb9ajptEmHGbcLPvuw5qvAIrf
bYw60IwGPJAC3iARKKO4N3YdF+Jjxf/t05LLqi3lwj+TvQgbu9ANxJf9C1oQoXyP
+uLOjoWt3MQIj7g4QYxB+m6GCwy9qZUOqau6zoj7Eqsa3ijmeCOvzIOP3kIgdaBH
4rVyIa8mzfsNcgxkX1eOj8Ac9h0pU4NeOxdMkWD7ObI/wTx9vpZy0O8+PLmyL45/
OqVUwUgBg1mmKQlyMTtI3k5r1fej/4za0/aoUcSErnbHI8DcenWQ0i8Bz4XSxXRq
dnRsjXOP+4FAUX7rrR7zWhVvA2paLj8if40qWAnmZa/g0miejm09cguZIBfzGvuX
0xh2jRMCfnjdEhtrQ4uR/oWKIsiUCX3i1/wUhfcxnKBn/Xf0BJHSWlXAdkybj5fN
2mFMZmxhNsm8K+LEvUUYlV7BI3jSVfkE+2bISnHf8AJRD59Er1lvt98+dQnmwasx
Vp5c3366E5w+ysYZ510HEQnkSJkY8MyClyNu14NaH9VOXCsvqaPBlPJ2d8Dl/buq
5bZsjnCmjWMn5iqRDaV2AnKGaFXihnZkfNOvRKQjOTGEim9OEf62TDwMUqia8Y/6
A6BYF7ZfhlLV28Mg9y+0re1k3aedfllxt2BJsM3TKTVKQ7HHM+aIwhOSGh7KCUcX
EEwSrD6UM9TdX7EzYLstOBVKxLc/4xcaFzJ7T+w6lxYaInq1sjmKz9c1S/pZEJMZ
TfG2U6YZ7goKBbPgz0z6RNF3AV/BWdefFmHQH8XZbp7J4j3q6p4FTMIr/GsXtkpC
yFfQ1NT+FuVzursJuqOKJT4n/qFfkFk3w2VFsxxUU+oPBaWolGI+QwTTgKaHymSq
cypHaO9esuAPVHi6d4ER/Zn4ozA2kta+etB3/YJog1z8pA+4kO11A083TcyFtwS9
B2C6XPZOlcRPb46Sb4LQgE87NmsFbc0gkytfekhqa9cwW6/JA8BFC2ZhK/ylZxf+
KeKr7UNwRXBHd16RdGG6BIjRB5SreTaWndOKSww/yyHwd3xW8Y1epKLXZfEFYkMG
BUPieDbV4EMF87FM7i4bl+zi0fhytDpgkIW7NyTtBHfsA5/o5F9N3SygZZZIKHKa
WsBlKdqO9bvewMtU/63QjVWMIS4JxhRtsWsKRBGUXw0vsIUUa/rWaAPcx1n8vhxa
47oIlV9phbnfq3ZTunxQWuC0KObbMjKXQ6pf8kCtSynaCr/zA7DpYZNQ2/pJH1GW
pVdtG34+yV4ISzzQuWTKpSnacTeXkbUKXUTwCNDW/5h4ljQZWatJrGim6m1L7Kxf
VWzqnIBpm3z1RckuacgUtPcCTVU4qiWc0pGObxT7Sqm8rQ0Zc4/lFekhfJA8Ty6/
DtF586J7LtEQh+EXRaUJVrBrMAp/9POlFlV8t/aRbP4tEhH644BD9sB6JhvQercg
5IUPxD6pa99Q+V5mFkiyn9sJ5A9CnVluqErMp7QFL26tom0RiV3nCtdhOUPUxnc3
lwjg7itwnBrsRVgUyMwleaTGq/mR3tVp4QCBKeD7lMjFvbpG8I1e/1ippk6U4ebZ
+7H/UzLw4SUVtDii8hJz/mRzrQg78Ww7IKppaLn9VSV4BxHRdL7NNbhL/uLZOtSd
yCgnQyJjKAPgLLTylW8MZ56vTcHCaAWs+5yBI1DXsDl7YVK+3ANGB7AkLq0ERP8V
H+BWlaATYNQF029lTrArrtRCnOy6LO5ScjP7YYiH1xTVxbepJA55Kmwsc4smokMg
0pWMPzSrvusecoqZZAJF994kiIwM6IkBbwr20i3ndR2erwtGO0sBVJB5tuOI0p0z
w2f6jjgV7P5fz0UbpcJPbxsjue6lWkN0qzaz3gm+/ChOXm2D3a3iMT9PzlmHDdiA
LX66mdD3MmE5pYHfwEyrPjQzokEJRd0uWvodiTYspofW+JJ566VJs9xqSTbiqdwt
NkDwzI8lUNR3j0ncsRGM77ea9pSVo2lAbzm9+dF+5FO8iymYrYmewGWfrHox3mf0
X2xEaC5AkHa9xCeCi/klGSLgUtO/GZBXNSChbKlfo58Q9sszPGKEFJhOJA38ICqv
PaMko9FxL2YyMa6leJQvZBiH2+SYOAFR8EsMOG19plcj18pY2H9G7rXulydgrFZ9
33MHpNWdXPAt2tRp7JGPsQh3IPIa4dE9H/fWcA7/P5y9YueaJ74+5hPHX03nVK1t
3se3fhebBFdxFJp5Rasat/xNPrdIexyjl28/NAd1xMZpdL8Sr4Bo+r7he4LV5TrV
tx7UKCmilTiNXvDZv1JumBiAZ4lXV3m682uNLw9NWQSxn7uk422dEngac1y0wMI9
AdcTSZXEHrVT2zI5En4nV4+bKYT4gqwVL6w4nATqi+KvMft2TU9PFKzMfV4mCO1N
Hn3i9Je7WDs6zHwqwwdxY+t0I4FaUYq0DQFdqf9Tjws/DXnvsH0LS65Vj3A6r/ag
ebQCrPOOKWDcBeO/E/7oHuDY0NMDQ/UpChMHoH59TbwviOH5n8MqwTkY9vCqKYYw
zgsm3JHzUg81n9xRvzDun/fnhYLr/rTNh+RWORgsaNUmEVj998ihGLFtuSvUM+SP
1IXISyJJOVa30Kfh5WzQ57wIJb7Sw7m5Ub179CTx45t6vNL14O3LJv6KIwOxd5Fd
uQnsdO+Az24xlJmdUME+aNt0rO3cLgw5Hlw6Xh21LqAT8yjK2g+0bqzI8/fQa1+O
YK+xbX4KQ+NgbXmpzw4KMgdW16ccOP/m9XbcES7rSB8l/7TmxyMLNYbFP49lzCWz
8QErWgF7+ZOpBl5tHxKh5zh0QwC0xEeGfxaGIQEq/33cQDIyv1uJNBmoD5m7I76Y
ZKQf76RhDXoKWw/bPMbqZenkcTe3DQsFAB/C95FM2ByryvRuDz4zGRM9Jd/3zdAu
6i6dqZguz397q9J7m30ipdIsXd1Whqg/F8vu0Qh2QOUkr6CL3SVK4HefLwyPy1Gw
vdM1JQyNdgyRyxvei4AT1W2IoMGEtJ7kXfVISw57fbRwGag2nRkCcKUU8XLF7lk3
dHZEhvfzN+uPkNJyDw4LS40yHvaPLFgFxDLBN9QSr61eyq/fSh/9swtul5/RyBbp
QX+03nmJWDJ0q52dpM7/kEkIrTXD1urgCQkKYLKt9WcEB29RrhxuRC7Eqfm06yeM
1Xwm7t2PSVvrLbCU4rMa2YPIa3HLAAxpfCRHMZB5wOwdCAgIGVH6FEhKbYobrj8O
2fStQ3pDAMpB5dfL8qtkmCZK/GrWznbTHxVzI8zvnVR9aEmcpwrPuh88bDXQBRKr
XjZA1V/WLGj9YmBXLZrjIvuIOjaEypc3hUDu7SjiqzkR7Cqjh7xkR9nMA08Al5fn
FZZICenSgMny8y8ZTLwU8JEmjO2Jts/YONSFhrP5h+f50gBD5tXy8l4D1m9NyD0J
Ag4tp/KclU6N+0gaIwqJfBM8cvbqW7a+JIprYCSDRnY66S+e51ykuv9TVHEIgYD8
HLexXadX9vbptGV2anI7/NzWgOIRYkG/nLPZphgn4MsVUOeHcDh2zzNo7fLsHhNJ
75kU6gk1jr8gEZi2yROTfVSp03SOSdvlmln+CXUzEJCkW5VuMPjhNXPE3aTro1Ae
Id4NObYOH2KIO3553TyJ7iYSMuIcJIoes2igqLjTxKVQ2vH+0lzioJrQtpUEIdOK
CKWFh0oev+ehrCDVGwXtrgpPiid6J7u/cmZPV5yoZEOypMzuGlgIVOlyEj6miAhM
R/pbVx5Y4LQ3k4KdxE7la3EVxUvnZu9y5BqK7hwEjo/N9feLgkgkpEqiiGScN1kv
0JFE0hZkhGYb+SBYfhQbn5NwTwlq+jsFl1kC+Tj2jwxboYvAkgqM0axerUanTEYD
VvVD7kS3dZ9WyU04UfEBphQXELZiYTl5FtmopQMmUqFOHxZUBXpCBC9UImlipB03
CRgVI4KBbY1dW5g9l8aNOKmDgoLBAB+Gflafw++2uxpJ/7FvNrc/NqR7z59bEyGw
PJQ3yyJVLcRFi3ebwSEmALpv9vsEwdqurJgNLG1fjpmFt/hpXsxew5b5Fu5O9o0l
/8FVzP74uhm+xNZlc9728lccC8/c8ymJTxx0TVRpQRhVamqk+IiXoTI5zxgGm8KK
n9TNs5mCIwisMwNU9DYlyxwAdTOzhxqbr5QqkhRzvA/IoAfYB3Hl+9BecoCVOoBG
7wP/R79h3CXTgxqWjOpx9mjfxYYIW2l3BlPnoaOsVt011K5suIkqQUh8gTN8qVOS
9fh80LQ//bK1dPdv2K24gCfStwunnzXRPcWHRKczcJAqUSHRgLHTjfHJ1NfGwMsu
bo+iLm6qGLjOPRZXgc2jqV6KpC5p2ZjUitJGtuAT0BKeb4HEXmJoDKjZZ72F69NW
za6jJel86DR+tvN9Ko6GJ6Q/KufynOfQWITxOS+vytG9cFXsnfw2R4Kz1zT2ifBJ
/dgehKj7SMrmQTb58TWzDQHkDr7c/EeuegwihDhdkCwpXAkJ6u80A6UlNMJxmpW9
GFPDYI0l4kbBgjuv9iNshKuZxEm0VNOiaXiflk/cLQdvTJy3VsEWEyf6ElFBo++R
65zOxSWacKZFomJllqSEpyfds1A7fGaNYHbhhw8vANNIDrJUe43hX6MTEMOboQq5
vNKv2DoDK09iWqxWrWIhE6I50sS5wbTyh2oDGf2y4pW9Z/eklZ9bYntdQ5wiDaHV
Y231koVhzqwtgHb2LlN9ua/MEGcQPgamXBYfopHhcaLmqbikX9Kyxhz9/k7wIUoA
WK1+5Iw91hEvvOjHPqNV/mMkGRk9ylZf2G0fnTSkvHRtcTaxPDiUDwBGL+oXuCk0
nYFx2VKQxw6CglL2+XUz7pu8n1Y3b0LEdWM1TEg1jMInZbHleUkds5oZG2CmKT3l
o+drEjBFjlYY6cSH21aEZ9HtgHSwX8kdOn3EMhMYLWaWPXAXIDcBemvf5wQAnDIF
qpBQ1Osr1spLf47giCHYMNOsjj2CWa5RWPRZPLTSUS17buIgloqodgULWcAriYmG
ca8/AKEOpAIW4fH5RVzOjO61eBSWtW21coe46HxMNM9VwS2JljFRKYjvj9csz9AE
DDxkv/h51oC7PNPHejigAW+kxkoHd22nG2B45qK4BwalfBubWTt0xhMYsi795mEF
S7/t216AyEvHCdJ9b7IQpmyFnVHwtwo3ehff1r7mptJhWGw4VznufpvLBe6ptlmn
Lkch3Ahz/a4xPK3wXJ8+F/XLS4R5zgvAg/WfCiZLrFNsSomEL8bPvcllf+WoPz42
P5XPHmy2gmDJavIBwbBSXSvJIlmEicjJ2v5baYsR0kX3mH4cFanoFAwhYa55KhW6
aHnUjob7+xgSB6EexROZFz3fZs2rCijjonudTmBEh10DsW12qf7o3QgzpzBhyEpR
5E4KCDuMOBIRSByoh8qkkhqO1zIJf5Vr8GbN+uWxHPThV6nFwrf4mV7nXBoQl3Wh
9/mdSFYOPeofl2sCZSrmm48pX1b/QuZQ1++rJs3YMERb20RhqMhJZGtZqyotqfbE
JKxcOh59RehPLqtW/ht9GZVdVxlK1Wdup/1hjXnTOIazoNw5vp8dKQLERPL/ftBb
UdU8AufVFkI6mCe6fexEtTfwgVdj7+Y/m6ZV3Obe7AOaIUg7d0Y3hYcyvP1RXZ6w
UuTIGjIe85+tsFHTIyjHMVNmkSwwzTZUCY+beo7+wiHXc70D2bqipbHmqmJjHC8R
EAjFBXN63bAoie4shUR/0ft+FRj+QmiMpdtGwJKjhpc8pl1ul65wzvoHMwecSfOE
pNzqRGujOXrrcysayHeb611nr6ghfXL2ucE2ZxIEOx9p1+TkS8C+1lTOGCJY4gRp
lGAORZ6suM4Ww4plp6kxVP4Aw+s9nlKJ2Y7XfYyU83urnzB4JK9wZb348Bn7OGxy
PKG8DGhKxIIiQMdWZwiHVJ5YvA60vekG/zcynF6vzjBzpk83+4OxKiItO09znSzV
zgWI9L9gZIV06lYc5CZm7XOQ6e7MfPY5c/lGkujRDMbzF7+/hjodHpOSuMbQcdq8
yYZ3+35+EF8RoNylawtdePjXF8qhqvXfX+FDQR6GnBuSRDZxB4nYgnr8VOQAhQ0a
icV8f7zetSpfDg0gMXrI3qFteyBJ9/aKwlTT6HurEuSwKeYF76PErCEVR+0tscIi
IihPZorTyh3hUskWffvz3V7ShCbnmpWuI+cenSKgsVrMnMO0ACpcWfDGCAeDUdJQ
Mn2rPVmDU5RxmAaqf04cPtzpf3SNonSZmub7MOuYWBSqWY/Xj0RzzuhDLWXbOhbo
Mwx8DTfSYV+4MPKsDP2/ugpdi02kNS2dWt3ggrR19ZK6GdWYyaYpCx9/KZwHvifd
yBoHQSh4ielfTytOmzsG8QOaSs9VupCSetweNDjeliat8+odOrfwrFS6ZCocBrOy
fJPb791/PJMC29uWvJPvnuEAvRFtwsGUOItkOguv7GKQ/I3aXw/n+NTJt33ydHFC
7EVmaJx0caXVxXqcOiUj485X4OSrGPBtarYBjqRYtIcjjiHAYQS1CyMGc/5SIjnI
TWit/WTrQxtUac2myje69ytIZCFPsOB4Nf+0LJSjhdi3xNi32HD1yB2/BVwyml67
swHZ3dSIAulyhBhr97wewtvmxwUcNFk2ylkZgM8f1W17YYZeaoHdDrIwN+l37u44
NWxBMnH6vn8QufTbbJVbvSiTDHGB+tgF8wl7oC2jPzrJN0agCeWd/zX70n52PK4P
uXFkrVYhYmBHRnoNhc9C0ujBr6HeDS28PZcf2WKvGBPiRAmI2LsUZuY3kXg4fdIq
zsA7SXWJGIg8I7WqKw71nLcNuom+RZkLmTOHppdU26IVuyu1CkznURtjjNZ6JIuC
uaPrfNxntj1HjR10ovlLe3aqWiraj5mHTo8QNR2297VEJriwsazMR8jrfgxmo29K
lxly0g4rHr3Skt3I4wsmfoRbpaxImPbK17oTOraeb8Q6NQS6PZdtRCrnDmci06/9
22mI1jf4fX+EVr5J4FiCcZhHj/GtWdrVLEkdyXC5GqXtYapg5Bug2LeyFwcR0HaR
opZ9gdeS0cW9HWY9CIiTpvNAsHwfDhFft1C5KBcgWcqkUlkS3krD0igrbKhJudzd
5J4DpptumB834J4pWo2VYqtFsjaLgoTNMHz3ECctts/eb428nnseBLOOAdLiwaa0
vmDRO/KX5h56Ji5rDue9kN8Lvh4m+s9Of1ri41eKWif8R67ym4jAGYaawbfAOkGM
7KdxmMF4/zkxal9v/0vu8Xnc4hKwKYYt070TuKDn4ytzc+DiDVV8W5LMA0PBpcYY
g+v6P9w/Te6HAY1372MhSaq3EadSw+HiNoiWZ6whPskspqq+hUAdXEIUgVUyEYFG
AzYPhErcJhqn/zikLCoBMgmCtfVURI3XSlZZbmc9cT7VNBkrnPiGo+aAMmFNOh/x
HN0zx8dcqTBapaNH58m4xciv8AjTf1HYc2hjuTPmyoZHI08vga3DtsSPDcfmEaXs
vkNobsl41RQb6ZCcm0v/Mtzz2zXBLZtMFaHOrzaZuakKLTt+0P9qVOJpYApnIDrg
dtjuuNdjNzqgJ7qhs/CO++Yw79c9mn1EuX0WnpnL6z3F5Ln6JWvhxdUCxj+p/vsF
U/qe9p9MEtjE/LIOZCgwv8O+uUpCX88caEqkl2ThsK8jyWa0pG1fMHfFKwh5jyTN
EZx2bS02ZNAkwtSmGF2sU9CDuufoKhhp936nt/P+rL+VEgw1OT/U5ZcJRAHB5G8B
XhIKIqXIEAVoJbE8oS+v6zp/kkHFpIHnZlOCl1RS67e0OQl5FlbQ5VzW2ewx7g1s
eRnLt/MRx96bTyT4XRqs0YSPQm7X9CCMJTqxXlMwQbPaNWniljVm1XjdMBPL3rXT
P5w3R3c68IKcdEz/4ousFNEIKIr3i3Q/DNj+gxDgZJgdo45u+QoB0ecfl/Ord0sH
BpcfzX1ryqvQov+UjUWe0pN8w6Ue1zwg4ve0Qh+D5I1GfNrhEj/X3VXjVX1YB/T5
dPDk++Y0TK46HVg7+fcBfCt/dhpJAiTzi/eN4jeXD6qqRDTHHb6pMxpciTfN2fO5
NtLdQ1OBQ5J5jcbe3V5OqzsdddMsfYjPC5NDY6DVWW0v+mxcZ5S2px2kPnlrIt7u
jIHM2h1+v7tx5V8LIkdiZXJIQUZSvRsxuSjlYukm6HgBmnjJpXXaS6zM4Lpgioqu
qAMmvbR5OLeS2dUr2n4pxX9BtIPbQmOStffT7ms4WKeL5IDsybdJ1XaybiLBiSyC
3iVtRfSWqaWoIiPsEUpuahCdtSWifzZsJO2VDyNojJSGlm15mNNe1KKdp8IylLYW
XZwo3KEUSeGriyzJ6Vdv6gR7SiqC0npLXCSn/S/5ebIg1yPthG7t3S7e89krCvxt
ypWUgmL+UHXIZR5R27593KVaelIMEtkNfdbIwkAiEWekG5ISntf/Xqy1E2TQzJSY
IOXEGBGY/VYRGvpgLehXls6KfXENlBsT6LrrcUwNVhEhMxKLQtM5aIp67XMdKJsk
VqimBZFS1/xS4v20DmZYeI1S+mgc4T1TbaAzPsVJXFldZ5g3X88TWozu9u//bH7x
qsjDo9982HfKYKJBzyfkatBH8yVd0fD0acG3oii4SzqAMEKGtFmQSEPXGUFn2tXm
C1N/Xr/FmJbkkaL9LXCCgK6/W8/oPE0mJk30QprTh08XdJ6WeKjIP81gQKMXbVRZ
aJPx+rMpXLacWxnMslOJg+ed6WLZ4F2KFbIyqapWCcnBf3Np/HWZ/6m+i1z9gwti
Uybcc7R5SBSoYzAiTw8n1dauWWw+P+k3M6i5gl+3QqJpizTVGmbxv/DaU73zRjLs
NqCEMtQ2ngZRLEWcCLvwZrnE9jQv9QkHy2SDjlf1JbmaUcGZb6c4KpiIx/15zQzK
dgjxOYvWjaMdA8J32PTdzK7kPO0Aah5vMmDvsIH32l2q7wh2gjqG4TjCgeMcR0Hq
+xHu45m/0p4RxPojuq48uftMaL4Kc0RzpHk9Kxq8yOXVP6Of0N5sUn7Fe0O3qS2y
DfTOtklhpt+w5h12cncdY4rQmnOD+CIgSiT4ZGCAVXxE7g/oZHrJ+ms1fOuZKxmD
W/MZLhiudWMXU3ijFfX1rDLFZQm/Viqin2nw+MSwKR8WDTZTw31N0Vll2r5BaiJw
BaGc0CC6f0oTh7HS24AZ30wla681sTXMm2Rcc1WvhK/hX7r/d+dQ9zRBCb/XKUvw
fREzWF9f1gl4ood81B3uhUOuZrxGf6Pw8ZFcVDWp51gtqBBfUguR0c6BVpYjnwya
wJPXmwhsMxK9e4M6DCrvA6tuQca+EyttkYSZTMTk/i0h1RSx70hPQzQhh8EEyDmi
qLpCZI4T2uI09PZQjTBQkmOaL1+1m+4CZFawiHegMvDJEr7UMON5lZr0qROCi5nC
RyVKSWwJAHJ569CZ3kqkWiBmKJr0Z3Po4TrVFU7MlG1IO1p04AGGre2JNn+7SCLd
6PNdNK1f8GOB7YEGZ+YS8sOTQ3/WzTjScn3KVAE5R6dJnpizt68avePmdwHOBlZL
mMx3p8zwlpEtuiYlY29PNPPhitMTBK2czE872KBGr04n7rg8Ml4N0WB1dEiHK3Th
IXvw6OFVdgaUJnHeM//e1Btf9VCDpLP2jJTHEMaEK+JyGlgCp8RHQhc1/CKzw1C6
YsOSxnVHIAAfC9BrD0uStFoeVrleACfi8sMAIy9Knka3N2Ywqgm8aBeTkdJFfDPb
WjayznqbilKgQqc4jxBb/UfRYt9AYZtNakNeeqzUKAqSuf62YvaX7MMsY01ug1ju
85IO9+tlOWHfCbLtQReTGrun5yvU22HXtTMAXIrnF4Nj+uHRdc8Cgj/UNOsZ8wSB
1cn8lYiGOpJJIt8ecyKkzGTANCFlxP/JDm5HSAfe2SPhFtQe1qhDVOcq8S8wLUGr
iCgxf5GjD9KzAvCw0Z6ls74rTBc7LdAo53SYeK1xbexuPzw1M2fPWgfna4aYplyZ
VK8Rf8elkUDTllMVChCTqCnBqP5/kdllh5UygPfbin2gAc/YqTTNF3UoqQkRVLL8
aTkwkbTJE/c/nZ0gZIzvkjcEqH9k52sZG+vmGe3J2QXL0xT2sgzyDjH/0u/FbkHi
rOjD7aBJPPZ4rQCNfpAiroxOJUjENhEAmE3nTOf8VF99YG5PrUenZjilqt+r1nxk
rD038B6oDyHP8b3+bu3kg6ySTYNGg1oGlzhqAteJ1ur34OfOQDR283/sExStgDnb
v5rRQmHkriBmkEC21k5/++nT6VQTGQrusxhb9ALH32FXG7appF1Nh+8Y7ShLpQpk
G7cYWmtvZ4gUrPPW7dCQDCHop07n0RX4slyQifPGUTyt467HJrJkpGW1Bag4AyiK
oYyRG6ViZl3b1eLyY/H/Y2N8KfVDXig04LMiHQTRAdJbuf7ZaYrEAKBICXrNJ5pT
taUDRZydTTFYq/Jl5KQdKBn5Tn8lzxmI3SIglhdcuQzKOlZMXxHM1Nk5hiueUDJI
TRYNMRp6Mqz3RNXlm97hW+Ip9KKlrPA5w4rkTAUsr+jA6mnpoGretkn46J9HtsEj
rNIAvlDQYNqNtx9caoqTQSL+PrOX7E3Qme6KVoRUxMP1T8Ua+Ae/WjYXXlaCXXVG
VOO/kCEbnojQRx7BUGO+nbhzplbNIGujbNPB0mptmyEz/+qBt+o78HWBa+3OOy3A
/oidB9yPA6aru7LxvHKmm+n2xUIPP6gqc/WL2yCwZ5SMOrpJL0vEOboWHbB7f46b
sGWyokq9W7f82EjKl0ys0bbFESm5hw0pIfBB0JixWE5BHz+2n2L+y9pJ3MCCj8Qg
Q6VdN2297n2vyG79mXihjp7mbaTqI0TGeiHQKqXEQDdK7E9rBWUFVX9mJ05mG/aX
+6GWOYzwL0vqCKMtYK+rJA5Z7YixNZoCpE/yhiOLCTAe5ZfISkBaqzb0lDJLyu11
pr9la0gfTg/y1hsMTOInOi7xRoaeodyayH18OBUiIPzbamvNh39vDRjB9vN0kVDW
SMBuSwwwJtckI8jDp42f2aucBie8gg+mF6rzW4oFY8zeJQh/nFLQfOdtXasZkz+Y
IBvE3aTeyEuWHzwSjzk3/JfGPIIAIUYnpJJn1NbY2L0ThzOwZ8uYFu/XBMXCUoiL
OnPvOplsECYqCFE0S8c8UdIkPPbBYE7ygekw3Q6/YqIFugHRjKNsmb4NOsvEi3/R
f5RiC/7ueTGDIvDluZiBlrCfsWemfgZ2kkkusfSV944Sxtc4qItET8LVYbMEj0f8
VbZcqhzAx8tSv/woTnmyLi+Q7xAT9MxBP3QVbkvzTGA+TLZpV8xWRTsIRBi1Bx+Y
ZcmRwEIB+VE5vzhwhsKuLZEfRqH5csmkUelZim3uv/nav7JIoBAhzPZE1jUxg+fC
vd+FAyEq5y6OFnOmsxS5Zmd6Og0ZED1vEDk6FQfDAe+DZdgQxrOJ4cV8U0MF9DRw
jHsT0bFyI6ELgqqWErncIV2q/pInpFcU9SNdYcRMSv/S+xRPJNg5NBj8wMSthIwt
WbXepkdjuChMq1mvxZ7pTONRElbCHomWpG16586XjDQH2deVZsl8cvYz2gSG1Qq2
uzi5TwDKoePBQiyqFgxk/y6TmusB8AFFmQIDtoTAUpF8P5NmT1KkUNrvJR4y65ui
W7P1BzZ5HcfuW1Lx3f+UT3ER17CD2KO9NaiEI/bGrTVyu1Z4J9o2B2UeQal5IkKR
iOiCfTcrampZa8vJCOcZzmLSYc4i5h5uCv0J+wOhdFnXJRFMVSbb5VlNoUAi4kDM
tp59Pc0EI97cOUX38qUE71a02tFXZTsawQsqJUqS+XT9aSw8ZJujGNIL6tWvjf8V
9aWERDRU8upM14E1Dvs8Sfaqx0sR29yZ4QeBl2Kcz2ffHTiCSYtyz02+yjlSXc01
WYspxCiDUj/RlHMIJm39jShZ1h04tLs75uLTMCF45eNE8cNZif1ubvSm0bu87RRp
U9NJsa8tXQbV7eYtEszWdzTV1kM+kmaYt4lm9Xg6oc0jieuTzWQ4Y02T5+5MW0I8
JnsfjGaLVgSWVM862xLBDXZNbEqn+6iUxPt2ulph2Qr1pGHRGY+waKD/6B85DqhB
5qrxukU2chnl9asC62TgLbGuYpsTpCWbN99eLwxENnLVQPYVTpCacS+7NTObA8Sh
l1B8UysvJJY/m0uBqBGkAbgrwedCQIT4xraZ/xYG3Dx+gtDIAW1CpmLloMWjxlDy
XTaWfaycqLRadPWFkRi+pjWUEsX4VvuepyViNK9lFLvNEu37LT7oonen9ctgJmeQ
Qkev6rOPOZUFte0tcZKjPPu9ilJggGIEeSH4VQ9nAlh3sD+0R/0FkjreqiZ2o/Fe
e09QXfoY/dNJeUcVCfVsCs3pxrTh9zvww8ljISg9PCPWUJpmg1lUzDER+QSikA6+
MEwRiUQ9MQm4Qy7KfQ0vZGK3WGwVT9pnhBXVpXD90ZZ5/JQJQA8s2IHZysjZRc2w
7+VGyEqpf4SznjgtIiOq+9ju9mSvYbfiKWP/CUCe+imXx4f/KP1jlTS+kVPErfp7
xNdMppn9F63+qx1G8OqOOCzlkehgwHt6iHk/GZEVr4BGNxmVZH64eUdfebNNx+Ez
CJvQwrfW5ysMv4ipUnpKul6CJAlyphh4vateXK6a7xPqXQyeYaMR6rhyw6Ww6URf
Tu4wR1Y5b4CM80eAuf8fwD6VO5g0FoeiLBCM5drbNZefo1482bs0zvEKB9gN5RVV
3wfYm899ZuNpZk2mcrTN7Vv85he4QeOoKsum8IE24rm0THkAUBYvZfdkM1YVMiob
/rTIJMQpJmi1hAVfVvSoaenvPAbneuxaynaedrEVLax4P0CCPbLFByZBXFe1UO1a
vPwPGC4B7m+kp272EUr5U+sDVTe5amkwHvW0teqsfERN7CYBbkZBTxzcLh0WdEB2
vfQkrLPIav6RpaOTYfmBobcEhg3nIcm5Kh4Avn3M3aL0PoO8mrCzRMOfLoPdZYXy
WxlUor8OP236uWKHsLWv7viPOT4kqVajTauLuJvVHkdh8tBsNTSjNh3v1pMfYJt/
/UyEztnuhUhau3hLl+97Pf2fcOD3GwYNwUJRQ+hd3NOD0tUSRfU40C37s43FnFeP
PEO7z+pKMsewIiVtBAg4qhNeijeEbg/j5+XFAirzeIx/XleALeAVgW+ozOGIPZ2u
NMfF4pDNBW7ahfsPYXHjWgwEOQ6PrOl+NYh4Xj4UeFrm0MsFnO2cxA4icgTcDZXm
IEQTgiK+WBzv98Znf8qzpoSH3Dok/wB0GlIObp1hsDr5OaQjl83UV3cYY549/p/G
UvsiByJmp4i9l1EBcbDObL8CL/Y4kdRWzqq3g6IWqQX3Os6ykqq8pCz8zMKbE+iI
rCRl2dVkn9tOiUKWSUduPwvetB6HoMASR/E1TzQ5qEYk1IfDZtKnObVGbvoRUN/9
bFOYHtAza0D7z+p0pi9ibeNngO+tAcBv7M7FXQ8mx9beIOp3ZVtxooxD5PizSsQw
cJpWV7LTMadIDRxO1YF8liWdeTLLc39gPG0dDBR4Ic647+43uw7P+vfNnjxx+ZcV
VJSfjweMEoPycCDaz9q2M8o+koB7KhI2APS52tarO/usIVWE0F1mRS/7alQMibZs
xi08ayRY+v0V0powgOTTgeO9Oafd/8BPV8eK4DkuyGD33bpeJPbr3m66jhWHXZhN
LCF4sOT+tVaFwf2nzpjm+MqoGZ5qaTxD1s5FDCdcJVcxdb3vBS9VDJzCHvWDIghx
z3au0pZmWJj3eQO6VoMeQ3X2ght2C0SWy2537ZZ+qFhXgyk0sXZ2fkK31E5QBjIy
t406Ziwd27eegUWyH6HoBTUjTdGg5WQ1PCBdJDTRGbfQYqdbkNZtdOenruBi20pN
3B83gWMJB1LA6XQ8B9k980WZnAUDNlhvShKW67nW9SAj1SxVwTGn+X03vfUlIZ9r
/kTd/yP55yaJad3zNozZZNhD0OMcRPLybDGd0zuszizK/cr7NOSXUZc5+yTRGrY7
MIDPD94BSvjFE9MyofMZDToGaPIBmF0xjwvUquK54rG/lWM3Obl5lo3aB352NXM2
B0AFl3xKj/QUss/h1quFp8zojoU8hOFn5/WrqEijGwr9f9WxxE7U46rEJGXw2+Z3
2T/n7IndB6zUxem/RV0CXq6QoIrviq8VvWaXfNaNzUzmeTr/6pYNqsYW8vNRX3wx
dGFUdjQ0GDxLyu727hnv7qELRoT+X2u+dt/Rrm5m0v/aeZBBqp9nyZ9Asyhki1i9
zaaSc/jrzhNkSS6WWv1wSVg9FUTMYGLSk7zZpYDgHUzEDrDFnQRInxxO//jBZiuE
rd7QhTmycoDDdnsF7PacQ0goRncDYqE6yIN6HBVqEu6A1xDBZhHkEPGFsDofTKDY
7X2X3a7nzPBIiEhCjYpovBQqYita5hBhB7hawgSxSOSy7nhOvwPg0ys/9y+DuTAV
SW3LSTfw8J7Pvdq2KW+bCNPiHDRXwkI1AzDKO/Uk8rBIyXmkg2bOGRyFtIYEC0Ja
9eotQHZcxX3pflBhj4Ibz9ISTzr6PNdqWf/Pc9T59gMdi/TCgIRvLd/tzVQFyNP+
1CkQKty3xrBYDb/LX5AETkGGPVqHhwyVlbRf+ygg6SkvROlr9cv7LpFow22wG7Gn
njkYFbJyQ0/CuMsF4augfoNkbJVC9J03foviuxt0oT12EB2XAoEVkMIqbPRmx9xy
L1fLzk4lR2YKSBW7y4OWWqn2SSqwsmWTfpTyJ+vQYwLU4LOe6RWUOzt/+8B+p2Yt
fofSuCTdcrSOSY16BE8WsfuzEUBgbFnwMNP8KuhRlkiHgbqRyFRlYaX4xv4h+tz3
OfI/X49Yv6xu4/sX8tKcjdBY9KBoPP55sXpp6CSTdZbDD6TQyLbcRJnRYAJg7Xju
YX3vhEfJZNdiY8ZXJgqqBpF2fwStXQ0wuY+JHgsGssGM7hK2E7u+Od8npiU2hP8f
QX7q8e8SQvrTylO+9mRRsZTEGdRrKmdWKQZQ0QzPHLyL63WKs0R1qR0cgWfvY0PO
TeZ2ngKjNOs7VAYngiMg7TrBbyOrFebbEso3nHysV65KS95I00AYBrIyYsTSz6Xi
taHb3LVwits7pzfActFweipKzPC1RRA04C7mDPXXaVCFGchDTvzZ4S5qMmR3bpy+
lGOplMiuQgGUCwOxbAItvtqowFUiqPA2AUbUfye0jTsSveOOOLQQ10EEKR03k/9e
J5iOqg34SKhhRGAKaYIefkTMVxLkMgLEs9Vi8VZB1M5F9k5oX/hY3du3+3TiFtJt
246LjTuPRhf4Dl3rHYgfE4/1amoWOxcKJAjGCU+AKsNmJzB2uU22nS/mX/2TmpEF
c0ljZWCxaBOo5IsRdSFxNMiAeLCNi5izQncfsFouZ4oNw9iHrcM7LG3lG+wyqKAC
/6VxW+8r+7IWzjMYfUtYsqDh2qLNeAeTuSDNiUMsv3diTnm0kFshTUQV/wOIcAgb
eaL669YJsypiRi8zAyCTZvtT7BzYnaskqknDlGIbY9JlbkCsldew+5kBo+JJ9tRW
VjyFvf+QMGQxs1ntQczxHcGWvJnF4TGwp1h/5AScFqgIcp3ObGq0p9+VoCTfb+a1
WPagHVAVsVHNFrVM4xl516dNG/5x2d9HwN66B92mWpSMUnptAPYymVGkK7xPhVRi
YqYiHXStBcfXx69xaUjyhFVp1AdHZdDCcpoLa5pwmcUKt/JVtFIJY9FT5ocB4nyl
sEV3cA7yMahRGAaewKhl/yjFjFWD/hLDs128KuKm0MmiLmVk4G9XKS83bQYomo9x
ckbfpW+Uz2YOYIvXsWckCvokrpgusodlXV2ScN5BQvmHUKRQwgL1tjXit2aElXg0
7reiaYfisur/NeWss5L+VDmyesMJdw0uUgmi6xIQkC7NVZab0iAtHG5rRMRR7H0f
NtVSYLezNbk+9/6N4PIWeR+ud6oMmJIdl57wl2Z9Lt+Fc5iuP0u9j3on4Rw0lhOX
59bImR4v05kLWA7AnQvl9TBdRh1oC+sCviQrbSY2u2GcVxf2NBeUiiy0kiCmDwAD
ZiWkTu2X4Wr0EBnpHfMwBYD/ALgEEMfBy/h0LuZql4FYGU5D2tnhKDPCFWHlo91b
xSyILAbAjkBfbRk77jQYxJ6eZVDA7eFbx5Uz23lGBCT/y7B7KqGvHETXUuP5Ir/z
gh8R64pIPl/dOvJe/stGzgjaIDElIombIFfNmxJby+3bblY+gzk+j+tCdrzZrZ5k
t21ZjhRSVKw4SsOfCqZ6+9/dQY03v8zg9RsT5wDyQdAmSUxiQTpOVTyw0eFczVIi
NJCkdQHHTUMPMGdsbErBxBoza/eKKxMDoweXQwpGucmAlGYF6r0vn31cjaf63HcK
5rAbL5d5l91QmXWgld8q6anqCzCKlqH1RC/V87YEpul1hGIFm9iYyrXrvc/zl84z
z7p4vCQoyXkd5jmwQnvtDG0NsqNGAAkB2jWECuUzgHMXF6ZAY8CJsjN4RIar0Db7
lR+xOAMncU4XlaYFBlqL6C8zlTds4ButWt93J2Ca0tRQpk23moWOnuv1lEFuck5I
KTz2lcH2Xlox4UnAA3coPXI9Wzccke9a8o/nZsxeTWMWVxcZVJDvBSbHubLAhxd5
trsWHFpfS8nqbg7mcxelRJscyeMEnYIKlk9JZtjglOgUrbb6KBt19wW9t/zI+Pp6
y9BI1XslBXVMzpBnLc9QUt0ggajaA+ZuSaYnLyPCqC9KUxCvMfIgpZ29Dx4OeQbq
qG7s5DH2pCxH6tzolx/qVNwfLfc2VO3GqYZ06R33cXYBYEQHi0/5Pnls0D8ena+X
2SKoU7GDrJganYUNzy9nd/V3dRu24+ko4YCAA+4MihRyumeiptVa7jrMFGVqvW7c
GEn5uOp3EyzSmN7DPWoYy70wWVB2j3h30gOGp6pwvU2p/7/LHEOKDC3n139GJmcM
UBFs4zm1wF/mqEgjEZJ4BJdiGxZjxaV+mZYHoBP5LyaEMlcYmoJeojMtudGFU8UT
XVrzxA5WJVPrp0emd6upTdDdxJ3ol7SVmaIJxhCFKgju0Knt157+P13+DDdjuzy/
unFA8S6/S+6ELu7E3gPsE8yPbpgg7ClTuekxe10659Fg+l5QEZ7NaPolcKk3IRna
6Y2/XUACxR75nqSebAMjrBOvpZ0LP5x8+W7h1eaBDC1RlmLQpPSi28bCH5P8BpgA
PqzlmOp2PwmHhkvqh3dPZ3/Wern31QqbBSdSArIKpuF13RCUOy23PGOMTP8QiOFs
sRsdfYSpSAdsijxUG/Pk5p9o1sMehcrcw8LkI5Ympiz/6NNHEGDxtGRzvtDHgvEV
i7DLkXSnEEuzE4EkBP+Yjmn46LFQBq7zyoP3KlUM8JnjoztmNQ2rbYM2NHvxvk8d
429AcXxjDohCyVQTtqAVKscn+Na2v7rl5tLiScYtw3BmrDUeMvqsmwz+1SNO0mBK
GVyWgwvMj5qnce/6UjIVAxjXPqEPTdD6E7eP2345LLwiGJOm7f5PHY76wQSeFhtO
VpKEqAvzLSp7HW/JD6qJH1vj1FV8l7fcUURQ5C8IXOdg2HIte4Z5cW/l/Gyb9RZR
zgGSVjjeTzILBEHMXQkUaj3g3ftn5e9/A0aw0pXUTKIPWCUJ8WqXMHP1m9JFDbYp
p2TpX07SSeGSm3vsm//N1bJsgyXKI4sP6/aSBOOh2Z1ilDjAkbu745hAMRE3OPPI
csVBgOlxtlfVxLo7HDbUs4M11Wi40yoYeUr1Mh6IvRJUfafpVOc2FK6CmfUeBBWs
JzEboOzn/vf55t6zKvqINoUoycH4szSnhpqd+Yf4iC1SMvGlnEtNVzLcDclLtqZH
8LSzwU8SPLoC19yCrHrCBFRaqNNXZohhMMSTQrCrgYEJ/GTfKDshi6cH6hrzAHqo
lhPAtlTRHPUpDiYNPwVCPjbU4oDCe4b/g0XJFuppTwgK6SwC6zZS2129b122dGoG
dScC4IlPvyXJcTYdny53GsPm5cmiUvh68Xv2+6g+eDt4eIi+I7jgxut2wxv2U+vx
3Dx/bOCKnYpIB2oGJeF9blSvDQLaSDvxLpCJp2+lJFZxlX5CRP9fz0r9ljxp9ZlB
mHH3SL1/9/lN1DTOpJDCJPTfXXj/iYSCcvI/XS3/k//N2gRKd7PJM4CvO5VLmxy+
9JgH26hplbNxI0Hc5XC5nS5Ui5+7MJrED/GJ6ConRfv94L8xEpT7grmrgXEOLjkk
eFMdQYDRTLnu4BCysXOb/vbYukSNMsk88P7xtYAlSmlELv61IPkIQU8NVgCm2J6F
MOflUBXN8Fwp1y6Hius2nkkOltFld9YO65CCCzcjYBU4rXYKwqTAtDqd21KmoBJg
mSHJbogeo6uJzchKiFBOJbG7Ohu5fHXMOtRQckvdbUXVyIu0haNhhkiqo7ZWTImj
XB+LeRajBOrwvD1y/SmX0+ydO9dH+KVWap+/ozsCpGH+BzIofCdRFSehzKlaQnEV
pnQczWX1/pakIDTZPTG2f5kogQht0+77oUqpSGiNPNhP6sObFxNrL3MMFZQzPDXp
oltaRYYhKVvnUSqzUgC488oNbgyc2kwWgL6OaB1sT6kGyeJnabeZxUgTEUghyL+P
/TO9bmJYFmYizKhw8qGWLvHOUUVP4tOQIZ7PYFJvgPgn13kM64Eysi28HFmomM+/
cxafZ327uya9ZRdP0Xsz0fX4J5wxLjZazMPxk3otiWZw7BNH8edj2tuE+YCgmoD7
U0v3QV7LTP8jWN0foW3B/gzXI8Pep+ZO6nsEtoGTzWX+nMKdyF0zYdUkx8TrWadF
kDP/jKcCDB+xjaBh05+8inDj1rn+h9SUi5iibhWbiBAedyF6mXrNvoqvy5GJ42v/
W/sGSvTxvInSnVCYp6QhoBzC/FeBcKS2XdL05/75gDwb2+fP/s3RGMvgMKwtVD/O
mpKi9dAI2pwLYIdnOYBKJFTpBFWHe5XwVYuIZKdfiFAgf1svEi4l5kmkfkNe6cxF
xaUuCsYnmXhVn7r+Domrnjrq/nsHJkdGrV6JaPE/M/sv0Lx4faSv0NkEMSw5hLGA
yJVDvPd4QbUvDQC8KE90+3RKtSfr+6Osf2f+Sax2itonAPTwTw+gbfbOWkxVeDW8
Mmjxx2BF2JxxcYbwfpD7LfMZ1BrABETWNcfy94U28ts1puuWu1rAH5jmekIFf0+f
lOB68KOkffJDknOzong1Abc/sSSg2cUxxdjuxj/2W1aohC6fgQBX94Vf7nL0HU/i
T1/HaXXi1rQxczPPT/ZZvkk/YaykpHzY/xdJkDF/+DQB+JFegXqdDH/EO4GXiZgn
+S4/+o4NZHuxJ7fJaU8Gpx/g/DAPPzWHL6mFIVNyExIzqSKR+LijpevY8aTp/4f4
Mzl08GYUzze78+YdW3SaB8gHdB7GoEtrW6iOQVoTSDaCxgp6GtSiR+o7ZnpyqkOK
1hCpTgYOKpk7zSDUfgBnEcz4BJcsIGCKmt4U6xSLRmS20yWszVC0bs/fwgIrsToJ
LOPD2FRkzfVVA629/xg/G/EwKVBS/wS/+SRyoQBFOn/MJpBReDs7bJ/g9nQxmcJX
7rSsw2z1ogwhO/eA8lrkCLBMJv+dFZwPaR+YZH+CMgXkuAUsIuGbZr12kb3I2Epp
f5Dv9vpSR3Fid87w84azyAfZb80T9c0cF5r1fwIJn39ASf0QYNiQgXz/4wJ56mmd
7Q8qetWkqauL7U0bj9vflVUa39RaEQmkg+Yu/SPF745TlEBIh9Fzqo0+z4RaTvGA
qibEAQ+x5lDEFb1znvKxoCNKbRk3UlJmkL4OvYgmZus6VOlRnz+54TPCE9JNSrN4
QZaTcv01rlsIAGoRcMgJIfqx8xbGgrTiJ5Uz/iACofbYGX5A0F5mboTIELkPJ40o
DarOiYCJz/LuArhA9NNxy6+YowAqvsBZFM8TlXSP4BVxAFFtlR7M1Nxqy+12LgR+
+1arW2fSNJ0fdR7DuZ4FSJTxaDej5MiecMm3vCnY8qUXVYCIhLI6SJfx9lfjCILU
HwSgoUza+kMAc6f0TKdQ59pGiHLIpgmradZopDnYNQlGWKdFwkPwVs+qwUHxugvS
q/liM3gvBciO79vuVucwqazMGSGY3CgAHIVHwYnjdEvpU0yOA/8ceHrgWL4UPg8K
PCrJ4ivy1VT3ZnbJCU+S8BzdziEB3u0070XXFVF0q6PPx5OR5lecZn6L5FkFpVxy
AEow9OMWniU3ePy5dQV2ymUEVeWdfZUB2vID2cOU8Y2fNiCQs/NotUwormxcCSNb
wnHaI+M9PIVO1qCC2PwjUPoc4ykewGfZ55B070E5jJ4Dak4aTrpe7p1d4qX6JS8g
Ffh614hpox92bkTOLBjWYbNwdHrUlCru/M//85r2eotq5LmCk+i0Q+HXPFB3B/OJ
P7RPuQRn9PfkxfcyTJFNElg/EE0TmqTpSQb3h5fuB5dU15rUa33hKOERhrZz8lx9
ycWCgSE1v3GuPcOsmslN8qZlt2U7Rpr3Q6CrZQw6UCJOP24mqPblUdjQWjtiW9Te
YOnqidWdotyenYrlz0lXjpQMtY8a03Hhh4xBE25lP9acV0RE6W/u6Dw7UNmyWWPN
i9muUnIwYyvawwhzQvFPtu9EMLWZO68gFmZIDA0l+ifEJ6eHDFn0jOQiqJ/jhHeB
Zmn3hm7912rRyp2yYa9Aal02qurMZoDkejkFMK9D+qd56q2TPZ3YVgulwePONte9
IYWOakG1BWP3EAV8TG/gX5P3iH86W6ueRWYuAcQmXEEXZk+2rYXAl/HLNO02m3VQ
QE67mhNbii2gm5TqhWcD1s1+ujt8yvY2P0zkrz8MWfBODqhf4dQyxyZfhJKhGVUo
4EknNL+pxexnJApHh0JKQqC3cCfOAWBVG5prs/iGdHcKHPWvwhJDOawhEugA8ugb
rLC/86Td1q/Bs6kUg6IbuY+ffHz6/FC0bFVyift/FfkLfG91iHRvnWSbsB03cfub
jwZCxZlY6JS9G9eDz4UwlftZDc2IQVm1OTTOhQGqATF4DCPYkLYTUBMvUagsEETu
72DmL9oY2jQ+i8kNfmOJRUEE4YG/wUwf1sJUD82VDX+9BE6fiwt8OtgahYMWrsh6
vnnPcpamIsgeqWYWVsh2FWZRU0CLJhbeVMFVP1wTkZ9yXzXezKyvagNj4Mb0xGYq
qZ0Gj/ribUscsOxzmgRsQGTGED6EoZQ+mn1PGVg+lTjexwUl6pKmqbUYsBtpwdFV
xQ2QjU22ZMS/2szzcuPbJUyXxPEersK5WMMxyjAUrHcoL9KrcUkw53GjNdk9xQ8N
WVND7XVOElpErRA6ZEH8k+pabu0bC1bV0rzcCKN9xVLpfcQgf4+57gKmfHshpThr
M/2Z+olsnD0VkRbP+8D8IX1YTKWBRBeJBCrzyy1c11tcuGXd0vkvuX/EwAkL1XW8
HPg1fIPIKj2g3Ll5KN56EWfEg30L4QBR7WNzvtkpUtFKvJBu4qVBpT54edLp08Ve
vz5sRbgx58iGscNvm6+Y27V64KAwUzUTfvYnpBA/Y2Cxkgn1EquOrZGqeOPlFOe9
n1dX9y0zVlrxD6NxcFBI5AnFoRHCoNo+wF1TXjPLLHr4686gXnLdVIPtFZgKhf2v
ChTWIKsiI0IzgXP+FP/9kMj12dH1w4OCBs3C0fTtRvBm0ZuW68gpd0ymRv3sk3bf
EkD1oppsR5cqGm518Fi0jGAqmbpILonWu1EsNDqoQh+V8/olhFuQ/m4CB6nQ4WKT
+PgSgkixeKCNSrSuKs3SWSqLmi74qm6fwrTGNcUwWmNWqHHDarseADWvNJd6SY4A
FBBkmsbYNzEJjg2tbsrwV0VWENM6YuD5kCw4ImLrHrwpvCJbrL3jQrp4rdUnRAdS
24ufK8+FBkUxLV2HTZUdhg3p3dmstJJqRJQsbff4V7NqHmM0zWMHOoqBRJPEm7x+
uPrZH6D54HPoAganSjdeecZv3MHjoEGSI9yDFw6mxv367sIu28cRzKK4GiEffmz+
7TCt5xvCdYvS0ZOTcDiBNpUXUWzQtDutvWTggcj5Wqj3Z9mrDU/O9RV8WmZiMuKE
7yhAspZUZIkg9u/2JNFqtZYVCCja4ECM4onOQWhxrVdrLWR5wOn/r/v+3SoWDDBY
k9AeqaeWi7LO3xNXwrF4YCFYSDWPKfCQBuRQsJMkDFEevopCpmJtBslY6eWQVNXU
umLnkumL08saqakfRfFQLWd/H4bgz9qkBVUxclSNG2gT3x4fW1H3JhS/dYxms3IA
+66WAwhiCiicaY0uxv0guwgOAsT1/PsGJr/ZM569M8m5RJvmxwYfvUJtIdhqTo1A
FHPLlzDgYKme+UFiGc+Ga79h+pIulqwoo+Ev4YcGKnOgtz1er3tW4z3V2r6mX8ZE
r5XHRQ5lM5fwmynqfxCHH71ozNQnvNEXj0Q8xR2ZSXy57x0/Mdz1uO9xFLit8Hs2
oD7kqrkxSDKHU6a4HdHCrd6jCj/xF32etqEylLQDwbBrUJFpIZH3286vM9xNXnKK
0PPTdCEzd5+7be60mEpwRSjJu+8dNYtoFPVGZpsS/hrm76jBeqJRxaCKsJZlXc6b
+HRcyXbYZAfgblf76pJAekpzn/SeIfO7WBG+hGnpfiNlIW2psh0dZ/Y6gEgBTUhl
Cz/k9Dpb348F0yaXv2YgPkL8Ei7jE/koWVnU4vkIDRaW3+9khIMpvQFWhkM6CJht
k2KJO6mKoI/AevvPPzVbOEzRn1O3ZG3hm054oL3QtnjmYUBAoOPu/1Mp+PGq2fa+
ulKvswtSf+8DRaxOSrOXlaK7vwPnRYj0ILPcHkj1kfKE2NK1A62iTbhEiGkcwBBg
+1qmNUbj9WE91dMT+YDad7dofLbG61DVdW9dKK4unr0kqx6c9QD4i0EqHrETYRja
jxgwkJmIT3DuCoeI0EekW3LIxB+Vq8982qqLImqw28wDO1kHuecTGDR3nQAbRouO
zYhbOb6BGvVom8CtgKJFz8xYLtOITnA5lQuVuSLHZQOnTgo6i7WYyick0jQXluAB
zZ3M1WD+JzzYXEGnaOg42FBuyK82x2niRIU5oHY4xPYIUxS5AAcsXJeyPS6xEzTt
2Hjusowwg/2IwQZE6nxCmcI3w+pxU1ycRi2sJoLdIIly40iCfJMBdCk8OJJ9fFom
U0Do5+EBqj+62Mek5xrrpkfHGNuEurHmQnJssr88ifQ6H9qdKaBsEVsPuc2s6Tbr
pBhws6FQrw4ugRFjdQwUpI5tfVVNZuekjgUEoEisW+uHd2c9lfZIn8HRjbq0STNi
dNeTsLqiG4CWGyxwzt/NBB9Qa9UYpF3nmdGCFGbBERu8u+v/fSMwAVLVN1xx0n7t
rLq2WH+bhez1+3pg6Q5rScHWM6837ErPaeI/mzRItZdRtbD5E9XkfzwZwaJCvDOU
lCusFYb2WwUQ49y9sYcU31NRioQboUNiKKXDXBr+936Ad04NqC1L5mnHF1ep6B/c
xb5gHG8MFz/eteIYrKrVtcBRwYIu38X0hIM02wRagsIUrnHKjGSynVPQmQhVjlxs
WY7NgHP+q7CLgBv/14ABDM2ovyXGbLmFufccc1EHTCFhcMrB1RYHNP4kby4/cUL4
wBkgUDInXQTl8Q9y4vQE0Qcf+uYaaiJCd589M2KPahECpCccZWbodqumDBaMiI4e
b/aMLFkqe/7Fx7bt6ZtCNljvRuuO0mStpgslnUqKra0U5qgz1TRWD6syZW1kODsI
VjXDpUXnJJQ9KFLZCWfHCXKvFCRgKJBMmzt7Aicr7uPBYJSy1thDHJExnJmmBr8+
kmwHwQ7Byue3nzpf8XIEvnKP2xBH0OgLDH7TbL8Oqe2uMwDevMelUBCiMAKKTqdw
9RSYAgqK0JOP/SS0x15H69y34apnZP/BH6Z+bT4awssWuD56V+X/taQ7RWB2AnyL
c6tcFVBu5EzZ66hSY11RFoBIZ8jQy2JHg9RBxIHZlpHphcEXA8X697iMwdUgSiGD
hRYiGlbwzJxmtQ7f1mcKD7J6wI7/El1swsnyLv9aKfiJ2GtKdNKNBOopX/3RRyGE
PNka46tpzhRhwQeW4Hzk3VCiFutnw0Sjcteqyrkk/11fViaKyihHJMTjm8XPC+vp
ZuZnP5ZVFM2oapL2zX5Gf1XxRHfus467s0rCmpGmuIbXtsMSz5TFotL4m17VibDk
npBYpZ4QHQS2nd/R+GFngdrkxMF8d3dZFJnF93urF5FvrrRIe0tTI/lAxljwJAsG
VCcvVcnCq8+Gdmhl5O2SWSPOz9/nFimKkL4S0wADJbJwujmd5V46dt+7CkeghPv3
iMuhecS3fxY8EGE+qK3yBeVmHInpXE+yNw0k/kQIIxbqCrStENXWJCyk+GiwTeR6
BvoCqQ9eD2ufUuhToaIoxY/S0pqBumZzjT7gp8LKYMCFTXm+2xzgcwBQB7XSjdxV
Y9eRtp8z0emQMK6tPXPN4F9aZrNyXCa27OmAL9cixxwCSWsUzkxs7kFSNO3JA03F
+2rEm8Kwm36aR3rYYqGTQuPJtzA/74FJG9FCOtxEkA1a9ZDJyGH5fzFNNc/+Dz01
0UQZ1q1akMaeWODr+pA+JhZln0OOlqECBrzUombn1vpmM5FfB1tNYoYj/UlLi7A+
b9Qng6vbQoUU9zEUfgNUhPyBZO0yapAbn6CSU45CK6auVwdyXir8O2CWkdmu9vmJ
czpW/jGZspx2X1LIEPLXSZjgG88dXKgeJVCX5456cNcbDascMZsuyy55syAAPPgR
al8621EGQs88ZxFLK3BR/M75g/5RutOhkdM8HTO/cpoJpDa1U4Yvd6G51Jrjx370
wzf4zg5pyPlHMT/vRP3jSLnubE7ZRvgnmLXneH0Nh+sekY3B9FjvehumxKVQM4GE
Qjz8s2GaTEPaC+tInyAKMExCiymD52+wFueoN+5xZcUcfNPjPQU1kUhfydmKkgE6
GpaJeh7sp3Ziqs0Bf+eQRZt7hhfrMV3oyiM9o1CrECDV5JIFTxrFnVAmjSzDm5oA
RIRYB412jOHGVe2p1RNgdqfam9RWdxu7iOrujfoCXGUFCLk5RBPzPr/dWjLI6drB
QgtbN4YlUVHlQ1GH7kP8c5Idkb2kktMe5av+rsIpG61Fz7DXKDamczdE9Bef+niH
qwEJJrIQmhag98L14CCv0THR0DR4Jmr3hxYTk5r1PW+KTgcqsr0oQoMX8wKdIsgV
yORY7YVZGBaIFEFxhAlQXP9sN6iGCoCMpLV+asWUTSJPymmEMCXG6DDyDl9EwyID
gAb3kVZq/68EGb7V3usUF9vl2yARlRiZGLm02S9VzjKG07o57Nv2oTRfwE66RGss
Pcb4ojn0Z9FOOk4YiYnwYtE0pgBSIc1EqCZFT0oq6wlHZS1ql0GMAXKTe78musYh
uI5VCMJhBMUrV4TOzOFAaJYxwLVKlrRBa4Pc+YrA8+guKBNCF3cGM2SryhV2On5q
uzbpaqF2fPuRQPnfbmyF+x+LhkjfN9oYL3XsGK/v08Ymid4aNPGRYn4jbP84tM0b
XRi8WKYczJhVc8/swqxQf8pcDy/CP+HUSNh5YNWpRV+5e3B4zCzBUDzEh/l6aVcx
PNhtSUcFRlmNrwPAl5POj4pjLSq1ZKVoXWz+bf6uO3rge57fhimYeMDpjTH65dbh
APtL64CjprNZROXf47SWUwfPM9RQKkS8KbZ2eFqDExJDJe7aGNIvPNB8Li2Hf8ev
Pin/it/VBaUukAREAUeIFm1AADJhfLlC9mdyb3M8/PLooL6m8jc+Zdgxi/l3sadO
qeJHvgI3hH14TYSIHryCFpdcHtLdC+aP6H24VIdzQornChprSrQX20gwNlyTWQFB
0nP49w7bT3yfL1R0cO+WCLOai8WFKws6f/Yer9OpHW5slDfKbDJGEvmAOUy+MNk0
pzVyacMFMA9aL3OovCrw47rSResMC5NWMzdF8p1ao89tSUl7Ne/y8H+l5jtVUmp/
BS+/FZQ/mRR5kOsZa7jXjA1vrrzWQXIzywNhnxptrRtYD9dV8h4djqqQ24AsMs8N
9OjrW4488HZeRzF5qfdSIC6uPk/1yo7dTHL5Z9EKCUd1OcdIonyor9HPPvCMY9/f
1MwP7oZcR7ot7lHgQCYoHjR7Jy7npkwUWiYEDTgVgowAnjoBdc8fBUVyoOiH2dcR
jVO0nhAnOFm1cKj1TdygG9SgOtMzzX/Vg9g8ddnVN7pw/kvK/FvLqUoiCMESoO64
J6ImhrcUlINNb26zKQnRtV+KZuKtFo15fdBptO4RsS9HSt/693a1Dfnt53GGAHrt
6HU+j//LZ2uznN1Ps8x8iQ5un/RYx5zQGrR3LcW/69t5EW/a+Y0DDS4g7aIHjMJD
fNkAyqIEEwboevIfwwoI3d8kNy4DvTc6rjYuPcL+VYZpXfNke+W7awYR6SMKRFJV
9y+EG1xzGoik3MEQQmwyV3OZuvVH1l1i3O3K55KzNS7rh1IOsGeJI3SDnmVEDRjf
m4DLD3E4LbDsW4ThMLjOfFd3jP4tVXd5d1mjGshhpVpHop+UPmIpFbf3Nikn3+Pa
6UMVEfPhtETzSjV4UaqgCaJRmLjvt/kqDeRImv1v7Q4OHO5vOlZO6g6c+UO3DUcZ
4KgtBroMnClE7wbsdSbnY6LeM4InJECpJZKZt3+/zbk+DMZIBHR3xMgDnNBazVZq
L5FM4wsfKaPtaQOAUyeNhcxnfcU0vv9rb+yk/Ntehk+311vRMrTvX1c8XXg+8ChH
UAa/JI2SfwYGNq6CZkXA3uMwPjYdA+T8RdL4ZIKTNE7tc17fpCSN1tZgyG1CwzyA
jJkSH9Xk9AhO5LILH+dANpfkLuBTVLxkD91TghGZL3D9/WDp0ZHpok0pzmkqLZ7S
f4n27TIXS/ABOWoWU8CsSEm6NQOktwtmKn8ddhjzy/0VP5mSEibv+1VZweb4S+xf
DAnbX6CUz/JSYNYKvVb4gWJy+fFmzCHrHVyXipBxh4Rwad/S3DFwOayP7sQGrmA/
jHGBBaH3rBPGN2mkT0t9L7p40XX91SuncM5k6ynMKDqY8f/YOX99ikzNDC5TgbJ4
ZRALm3+L3zCNqyztE2Z4JN6osN0GZRxbpN3tKCHQnGXVbtItXoqGrCy93av//RX8
LVUfi1ce1fHhSFdud9NthibofuaYg76HcS1TjVfR+mtnMErVoQIJnxXFOr795mrG
VzaADFZMH0pz+MmrI9XifGuz3e1eBUxTeDB9MImKtr4JbaFr7Ec8mimaDYzHopLa
+Qvsd44sRAow1NhAvQm80HzGqZvIPQ0JQT15Ieqkzk7mN49hmfApiDnHngS5VO9/
eCEUnkHtBJrDN7BlgnZVrKWjryl5od5pCAuWY8nzDVN9PZCSZ6xLra56Zmjy79Wo
J3YqkiGFg7/CNmDj/cLKuQVjXO3CSmk7wbixAsRSc0rPTCCTGcYIKJLEzOztd5yU
HcPBasIxMEU6TbtXAhclW/OB4nWHTZl4ToPAJg8AKSSPQ9NbtFwQMgleOiPAOwhm
GZj0R3HQUDJatL9W3ACCR7kJrpkOoXUM+4GKF0yBvEjuOcL7f6XN2yZurz2lN2sM
NYIIJdIKQwudsSyLLxT0lErzIvDWr/BM/U56MkGhvYSMbwKQj+ojv2d/3PEzsx4K
KMez/YSsaQn/WzB92LRkFApCpaIjB6D2xHCzZS7A443uxpHn3ETX5AW++XpUt4bT
`protect END_PROTECTED
