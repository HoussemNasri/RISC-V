`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDzrhWUdb6p6KsVOuy7TZhTCrXp4cAFUsFc5zlDt5zpz6srfjS/lJyqMn5LLMiyz
PeS1+GWZGGCHaZvHxWWX36gv3w84Pxtn/Q1gpd0sSlW4dLAX6hSl68hFNTuYqjdz
537E87ganzDtH8Ex5QwhveupeukZq48ToVsJqayF8rL0ZFpZ7dvHo1zzxUcJ73vD
tvBebTPYub4STcQbixELuABi/8B8uwoHURUl1QvAE4xCWWVtWnoG1BK3wAUo4clR
R7iGkKauXOdh6ysBVk28NWJMYe/bTO+1u9UdUbI4sFPqts0FmcmAzOa6g+1jqyTv
Un7EulKPwTqs7YB6UBAjaVCBCc17IfwpGtY5wH5ozYf25fVJdnRpQvinh3koofXR
zQ3IR4uGKcLG5ZR5WZnmOTVjPMKl4w0YGRLpRXTNyGZVTD1dxpP9qZUJ2Y7+RiIv
oOtIb6o5UC/67K9lBUkw/jEdOi8d+FnzL8DgejsyFpI903eT59vPuhPycNPmVbs9
bmmp/Q/Aqg5XhfOsGPGhdxhIoUFKGaMPM71Bl6vwMC0Ctxh/UeEOdjBND+sz1XwF
GBuNu+2GO9Ruvd+DnRouhUgaXyJ+0iu9hXxAHyB89Go+P7H3pqLUfmc6cGqKzAmy
PTgktn76dIZgDQe/6awuKvQduq0gDKsnCoXD5Hoef9sI45x314a2DDDAIJuh7gNW
R4vN9QS2ylK8ZwWueISxEF7EANC76SoXRtgaJbqjyK442iZIio+zfI24ZtXtOH2o
RE6FLSV/QQhoMM51ZGSXn4lHPHz4jRzbEMSM2iJcYPLCMXP35CluqZJqWSphJcZU
0DfwUIAGlokcyg+bKdpV4LEn4zU3U719+GuWmihwKCdUv/F/jmScoZsl9NNnIhw+
s+o8aAmfOhNfz7ojkwu06C/J7X0WLdEnfG4h+sIx2yaB319NCJ9/4n9+u58yrN8D
MVcIlm5RUIgM0SHx33XWLbVzAWwm9MdcVnvcAwskiSALBEB9JkbmZLXe13xAXnrZ
7qjiwqP7WF6ZpHW3u9kC3b45Td/JYdDPEO154JvGsGng5BsJDGYwhqEy17W0BdZz
TXM3Ktt1Z7FLxffRTvji1faD1ja5KX4XZsWy6cmPs69qEiXGWA58rl/+uv5Q7NEA
c6m/dmFSYI5Ac5nJN5qNyNqEVUFIRi1Zx2Ljf1uZss329bilPGPjoyEf/RI6vcWR
RwggZkJ2Bdsq70Rr+TAubEbiJFM76RbqjLlSCpRccGicmK0QD1TmmAmHERZXJ9z1
nyDgM54wU4e3qQPoEqAA199OPae7Wy+BnwIIsBn3iRQGTkb6yBEz/NjFtQ52gRMd
YEqNuQZdVPlKD4YXTEMMDiMTCJKoqoRyr4RxVEroC5NmkvZVCnvJUTq8oyu7Bbe+
kZ9KnXwn6ZRagRHZWa+tXf6oUttQyKQj2iefgsYcRrn8RZ1xNHv/8blawdGEPBNq
mtsEpvxVFN6wk85Jh5+wcFDteC3Pxn8LRkUvmu1VWYHYF57OtIFhU6GuEe0el8+7
cHzpgM3aJQ4s5Ok+FxfNiO7mEh2+/Of05kbEF7dCtT/nVrel83wmSfpcTlq1xJYJ
FlUf9qyzl6G7D1RWwevY4ejcLv01DpV4Hgs5THfPPLD8i6F8YIl6W3L5gfRBP/MV
PxIC126qRZC4JZ/nn2rbwF1i9Q62FOBCGjE8bIcLfovwqmCjlUpEJKkC5i//ZpdJ
wl7zLHhRf6zDmBspbqUEa5bFCM0QI+u6xY9VLl+4j9aGUAP9X0sbvudfPV+NgH84
DOQlma1PRlIqv2tW6Yvl2pgYKn8xsPT6xy4ImBd4g8G6iC8wD7oDsBQxumo9PZTv
g+KW8fZ8UTkyiTXhAOkn/4dTZ+lFzj1XSGePkMY/K/d2vVt457I7KSXG9sVYBHz6
GTFSmKhm2hjQi4a5nknTyy9BQLBtB5nHjEg55JuxG7egObQ3DZ72NLcDgyyeK9id
INuxbqHNv4uCWR6JuPdC3DL5Z1hUtQiMTz03OUVSKs87XBWs29Xj5yTR1V0q5RZa
pgVHSaZoJH3LgmwMS4pPaWYaSJ1IiNw2K8iHy5iHhPjZ7G36g6EUZTuF6EI5NhF2
E63glfhYQAWbOIb++S8AR36QQvy8/3mNM6QnX1WjAcqH2ly6LBnyAcB5aVWmmhMq
CMbyerDvkzLtmAhq2WUXjAbcpFvERvubRZk+v72Q9hjI0AMINU7F9mIcUg2ZNH7F
6UCHvNqlRwVUmRzMk93H0OTj5u2rU7qCv/IdJh7dEjn+wKHy71unZb8I6Y9hqx5d
CcQxIgJyGt4ORjowQUrQuu8QcEvJdAFDTIsBegYb5c4ENQlP6hXbDkKOJsXJYym7
CCp1EmP16FC3V/GKA8nteR/1b6sGm5ZfOEPGOLdRC9COfiLinGmX14+OboA21eaw
xxeFgsFQMOYBGlOLXzFAO/0wXUEg0+XgTSvnrpi88NywuH8HtLrY2dK7vpjcsB22
h6ZL7RZFVCx6V0xDjD0eDM7o2BC2HmaQ8JlDmDRmyJO6kyNtLNUb3xjaZbGoRVRX
7xaoAND8/mBWBq2voTurSa9egwKcI6/kUnsOjyzh8r4US+htY9IZAJDgP8lD0Y9M
OeUEQSAMwJ4pmqKf1QPvGLw7JaXrjdVfibe3i4V4eSnN406hfKGzIqfVofZbWDBM
KIJpc3I5QCD9QEAnPafvz56xsWZ2Nf6d6FqcGHc83SPlCHFRdszG9Wi3SP8/FMID
pJRXzAqx9JTquy/ZcBHLwqyjFJ/4HvRv7EoipxVdfKIb763LmLO5PJH+6IJi4PY2
3NeRAF0YaA7/qleWaTZOebT+fyW0oUJHrUIMHW4Gy83lEqaAcjvEx0NDl5lNBDJ8
RrYYmcyoBg/QqmfImjfEftjC4cHo720yUSf6btLPDwzweOiU313remWUdve+8/xK
cittit1eSlbmJ8OMV1T2cLtAHT/cq/0lGb3ppAYHd6PlFd1dcsnf0OqPJEnjmULU
L4GekE3w5pfkO25GeFoPNbDocBFmfWZSs9d4cwtHZp9aFFQ1qxrfLIiJsND0RiJq
9doFjTdyyrqeDN/PGoSLxXyHltnbkdgKAJ0mLhgB+ewvzlxzQt62xF5YqXFszoNe
Xw0kzEe8ZU8aSCd05nFVrb3D7PtJEelOqYEbIL7zEtALllCNpynYpJyHpOkD06bI
D9Uc3+x5/GgvUesmVNdW5ESms58wMAMjlhw+SkMUIpGIRrVlKdZMXyytQobRnfx8
K2f/osFUjSef/DvYHRYh79/GrBj5WX2QqOFvET3Ycu5qaI5Ve/xuDOEWxFv6gURb
r8sJuKMxg+TmdK20/8hcb96IH2w4+9zDRjk4tWcX7MKqBgIZa1EbP2VVhabbrOhI
WYbgovpbcD/KFYZJQ5CY+JixO02lL+eWdqDIJPYvfYCvisDPtKoPsUr0sXM8jLoI
YWSssjqS6jAlyZw2d+8esbkAkP7eMux9O0jj15gCrWui12UF29vJt8rYjIrJgI36
l23Iwuhv22c4+areTK8WQ2Azlq48n42QvgS+I1bSiLAG7lJWyfHr370+Ttw4q0d5
Yeaot7uHsXOc25wJ/FftRKgkahNIzYeMuEOpm4n13dgXLdVxndbrnG2512wb97/r
ux9A28ZsHytg+vNEuHFqpyRVSHf5Z68O8cn8x6vu/E0GEqbGyjTYBLY36ZcvsBxp
gmuyGDLR3CYUDwl2YawteDxxAG80od4e9xkAvZFkXyKPZlFUIv3sj8jSlf4KhDOy
6S3eb5ctIj+dPiyG+AvoE5lcYfSrGBwtPGn/pJ+SwDKg34vif4fRTizKGWj197mN
Ph6tXFx+JR1yUZl6RFAo7wSw85wWSG66EQnLMDtrkC4OyLvhIt7uxTlsCNM/4IQf
V6MomFj3jQaq5oglSsbnvi3JtjSjUcVo4jhn3qG5SDtt7BUGy0IUgxSgjMkIT5+k
6q7ur8TNEjoY2A8OXp7gA/qSElWiNa+Udo/jZHVcy0sreXpe0gVL+J6uyQjQwxhQ
JiOjldc6gM7Fb6DkWGa3YQxKemKE24f2rjeoVPGt+KDJuKxbH0P++HgKwahtVEui
zMFsgca1/fXdpqj8kH8emaOjh9SuSpXqwnKER3CSm7ecBtlHUWuq5db+tltSldkS
fWu2O7/QUXNBsVC6DjHPAKtqo8K9fBXWNbXM2DIKC4/+APi574TbpqQhHpktFVFZ
fe9qIxS9n+WbA+CEbVQWXoFQhntyc02IACIxP9fINg/9ocli9a9+7z5HVrgP/Hez
2jEDGxIhr5tj3jKqvb5OkGwbpboMgVMmHsmFY1jpfrg6oArAM0fM5Prvr0fkrdXb
Sh2ZgZakGvZsXBMyIZA1G6B3Oq+vJzxzZ0JCyEA61Agp+l0kPEvqLAf7jbWmZZ/n
fG3mMlDMldx5cKIzFuvnvNCTokD2Rvr1vnWRtuCya/kcP/+Bck6Mmc4pPeox2XAU
ewoG/n95FIQkzgChuIzwgS4U8o1tmw05OfskdB60sJjpND4tEyRyeBMGkqBvH1z1
oiYJMbuyC7zlgRp57Bjb4fzr0mZyjlo1K6UiWwOk7k9kBBnRc2ys4+mjn0lysOmB
OMkBUQDTtXRWddsYPrMQ26GPzJjyr/uXI4R/rzqVML8diDmGZgC5KZX2+CCy5v0W
Yy1CJTApJhMazlZSmDjkzj9lp9xeMKqY/Z7pWd6m9qhXgvRenheNVpjSUQRCsAKk
Q7C33mE7tteb9wyz9QGxpmEEyAt1AEinVedgsJl7d3JGvmM8cyhzllUAtz8TDk65
K4qXwRd1aZvWzHFO/OVXT7DhHkHsW1u67oVTBAwUNvVDYXhJIF7y51S5aNgKJ7v5
kr5DigZBb9OuxUB8vBX0TaVLFxG1Okupjij6pV1fjSzFowDWAbZFJ/Dh2jmR4RaG
fhSNAA3ujAQEVcqedK8ekDQf9G40c+b6OS5nzAc7yjl8SbitDvlgPKQ2CO6QJ9lW
jV8niCUM3TZUFerkQ4aONFmEsUH6o5TtWdkS0xn3VJ0WspFNHjtg4Np8/ONd8jx1
P/yvZrfkMPxci4jld9078Pfm4kIYpoY99kD4AEJxpnmHPo71G7KlHo0iDJur/zFi
kwKlXgHHlWAcz8t0hg6UoMRBEEc88DvsWYjHFZJTs5WFsfB//3vFhFhE1lPaKgBv
JPgWJ6JAPReYweiU8SDkgY4/fqKfTzcZd/MI+OtI2OUhOFEHi+nxXEsQUO7Hab34
bzopbBYRnyEzp/oUqJw4GOTk6vKQ9LqR7liW7WU1tph1C1ITKVHbdh1A75YEHuCs
yJwK9zz274yIW3dBPG5OA5lk6jWilgpsD2pTMU5E/xuptsq1+ZT4ArAEGeVfqOFA
QtMxyP+PYNT+S2BGfWM5wMbwc1iWNVRHXSA8qN6IDKfm+GKGOKD686pKy4KsV6X3
txMMalLBIG8g+4+uaPT9tVcp2eER5D8NditOwS+WboHHMUuFxaK4VZjw9XfTznOO
eVUHhP4lDIa3L57qLNWwqs5tMMNs3E2PLUsMP7Og/aUpt6fUIN+a5gDAAHzmm82w
YZ8JKEcMpnhyttkvqw4RSJ5/lLsUlMgmBONdMSYuah6RK612tvFIgTQH/yGO6SsG
znwHxPMx5MWRAD4mlqzNNkMoret3Q2fUae4QyKf0i9FNk0t6XUAJ1doRe4y4l2qM
N1oVac43nzsugx8U03QFCMT7IrQux0IXlwFKqGD/ljQ4PNxUPivwNFTM2n56nH7Q
UnBZySpPsL5aKPhZCOLcIaoQF3s0DY2O5jg7k/vg8zFdjP+HtVGN18sYd2md1Yq1
AH4lkkF5sAVtUWpzLzTLF9M09KiatDngzG9qkEBO41xF7D7A9kUMYP5LoQD/4B6n
HkgpGV34JOEf9CWzVivjnL8jIvULwJr7Gna+30Yf9ms+qQjjsMlHr7N+0T9qUy9M
L2dnDNNtNEtXvJy6wk9VkzQT3ZaByp+mFR1GnOtKixyEyoHKHzZJJAjLmDWsUxhn
L/nFwMsKU5xxhjotH/N9zFPuao6dDrTlRNuNDvnOVFr7J+Wm2/RN+p2EzQIU6X8B
382LDCAdi7JvmFqT/cb1dNkUgiMItwbYxrARwmxJ7E6B1SBY2J/0jrFkDVBjYByk
90XaI1AInRk8+PrZWTjlsFSEdcE4jBOa+mlPb42GaSy4Q6549Ejkf/YdkaSiL34z
RyHeCjrlJ19i2KpZGbhSpRzSCw797bNuRn4x9BKGJowND/0SJfyG2sETe47UCdqZ
HytTxjZC36kcl5Ly6txE9Au/40cnVB8UeTPOJS691Ah2OIbWjJ8pTjEu4zuocdNW
AEFM3KfGVFyUfN75gFeudv684T36nWJhzqZlqPMwQxWN9GvM7lkPY63Hy6+JizHs
97/f4jfqBLqCZMvdBfvPSCaUYwFR4FX97tZJYQ6R60bU+sit9yKWO6ey1xWa/4Ip
1ismiN3FkF18TCDKYaYAeNgMVGlwVq2kSQM/Dhb4MQNxIGVHk1DB8Uxy3mqHLvsf
AtEKL4M/wPGzP+e6nJGaDEiZXB3/SAIIe0Wp8Br5rqoWELhDXkD17YPiSvsIZy4t
+mI+oQtrnx9BZICI5PGOLXRqlRxusd5kH6oIoizmDlEf0hZBb2He2oeYMte2Fdxo
T56eq40OhJsq0JZZqfpuBC9cFX7nZf0GsX8Oa1ME+v1CUlOydNOmLCTPtzJA+nd/
KVUJnvm2un7VioiuZDYt2eiVRTSf0siLjVV0kp4jojtqEqsmdLF8hAI4Of46okTc
bB45ZC9tHD/FaPkDq+ouENNuuqoOV/V/a9cXLn1WMKwoEK0+XsJqrGHDZvZ6HLGK
Y/vCtK9VMPuXjAaaNF4g1ADlyuWKHyuQlwlGNmr4BZ0xvcrFLkwrEW71Hd0eTck3
G2NkqMNcWYW8URy7zKMmMgXZLXC/kHTPXf4BhNWLDHEkbe+IAOpcW4MO96tdx81t
tD6P0dN5CdlDFbMCA4HBSV0bSGhqC1qCL+L0NAfrq40rB1YwfqC9oT0sMMlzIfjc
7ogpasYPXwOWxINBCnrBv7A5K5Zkek1cK1duX8pBdzEb3owKZOMKcjQxEwMlGoTz
oFgzKtXT4rx1KV5S1lhYn9Axi2MNLrkvvU9c1iNhky/jVfqXec8Zkv+L1A6anHq7
o6UjQhcI+nVdIZBFqe5coTQ8rAMdGhirMZ41FiZkI1fSLRSjquYz3o89psfOEql3
8WKko8+2dTjxxSbev7VMb2BniLDHsQtcFS3HNkPeloW/8N0zoLVBfjE46A7186fV
3hbQpnqH2oOPHS/dQf56DT0ZkDWRBLzHn5EE9Eol4Y41dTZ1nrwWWVBptRQA//A4
+tFkzigKQpOvJmMLs5fV7f1P9wPLYjMHWaqgJ36eagxynBFDQ1WVHOo9wis9a9kK
N2cIeD/eCRITT8CA8gu1N02ddGkTk7833C1jxRhwIsPvwkgznuilSaAD0Iu+caM/
CisLURXcZes9TKDnUs6aLeJITvwQPB8jad7vk34kiF65IiEBoR4nmNI5obybp8KZ
U/vmOqPViR8/EfuQBs+5fu8FoH+gz3z4hh0Q/BqUcwdbb7XJwieYJ/xn+Avw/rbR
zdUeFBPqy2EJksQmamrSA4feYPxUCI03kLGDnesMwtogTmKgxr/F7wiTyjXMSW97
oLuKbyNboFn/zcu1LHxFxx/4/psFYq7bPr/VkzHYVk7P+OCl1rzKPHSQ7ae3L1bX
5QFDYNimvvN9YBDQB0JgiT374jES1YdFZNMXutFt3QvzxiOSeSGvyMY72xgiGQwn
Bj/ZcNaubbVkQ21Yi8cCa93U/CO5fPaoZbPDxBM9Z1aMR1ZmcWd2roHY8yBWDfFo
D3QaUR8yrrspg+BlKMYhri40GMhi56tB181mTnkkXTBQvr0mIJDx81moBrglj1Ix
1+7IJNl1hwUiL99Ikkx9tmUo6y616VPGSIU6BS3bauOYf85T20OcbriKKEfdmDvO
zpP7Y4xCsrZr4B7nNCSO1xXTZzYwqB8LOra1dCGa7YxZJMocAQew847VuNKifxps
xob0/K5SG0DLSG+PINJQBlYX3e1NDu7mQvrSioKqbtXolFf4J5+8NtcyCHrenKJH
UGlRpI7bHcZz/DBLNlY7Qj40djSise+ON/04dVVu8m4nACcNKSOb/mSjMiGP1aDM
2C41ZpX295z645cyA9/BOULHdGcUGcu7C5cGj8Rk/wib5vkszWkq4qHwNDkGPyL7
0CFUhE08LQJ6wx76d9U2rOyRY1oqHaoMuRBtSH79LIZQrFDJiOIlFV7+fjEciJ65
Yiw8y0hFETbaFZtz+CaE+xzcnUUj7kp26g9WIk8i/kSzFly54PI753+4SyuDCO/L
8Xlr4HtG7rQxmSCOIlW/OwR8v5v7r8Dp0rXHY2j6GCR22aYpe6JJRvqucFjSEhmV
HJGAhJ2E1QhLOxJq2Yqtv53PkP+cvAseKWwz23yJ8ozR3J1NmUKJzWUDdx02vwRt
7mD/L78nLdYcilAYcHxEROyU8sPlTyLynrhhW6cKJQ0p2LIDCG8kCH8gEbdkhVq7
adcvr3yyEhIJZ/NQpFHzFCSCCyObXnfy1CBrTH5a7Pz6Au0Rjn6WrbTb4qi1zHzM
04H1aWnXHd9+KNxorvqqHRTmHclNq9F4v+C1VNz397tUpLjk77cIG8HyAIGfYJcS
p1Zt13pGkUwEudHjTQHFE72a3HmU6RcuotddThLrQ488+GBohK0sFaf3qUfGXzaB
W6ZpuUkYgaXbHU0PhOCD89WQAu/rBuV3itp1hmz5oadSuJUgJWSfGVRI7VUCkD5K
vmDBY5jukZDh3lLk5jtYw1LFU0WLg+bZgZ9LkOWNnPCRz7TCqDBhBdb9KRDrGLDv
v+BHOsCXIbBCZbP32e+kg4j+xjZXrfWiZnc/6GttPm5eAebmQsvORs5nxU7WtpC2
kvD0w6Uiq0FI55y0KB2Z30oBwQ7RGIn3v9NlGJw2sov8Kx6eg7cw4Z4KgsSKUHc2
U9Y+4q1YO0p9c81XaWkihn4gui95mKZfnGbthU8HQ4YxnQjFIXnpPecmTCMqx8Fr
61/BM8rmP/oM2bameBoBNiy383DUYaEUjx2hJ39ayDUKAWcK03ZbGMoNDV54CApk
n7cyQNTOQEWgjV7Hd/ZyyYOgge5P8F/4wi7zQUgbxNqcsQuY4KAwfpy55svWmmpf
+pKgzcn0tbJok1Tqsm2M6p0QaXxck/XR5MZmS4BRkm+hEBTkxz2YhKBFcwcX55wd
2p4Q8mvm7v/xB39Dak/HfNbRwlCKtBesHNg79YwtYYSkZe36M7J0+Ho7jdb4OOn5
+QuX7+CNEVWjPesMwjOVAjrZIvDlFY/q4t25S+Ja4FJqXNX+O33ya2rRgFNZsOdN
5qIkSwjmFf/RfibE+yrywpx9y/yS9BThW0NgRqBGb6baRBGq5u9iHBt3h1nRY1T+
zyRV0D5AcS1M76UNkKo1TfrWJmvMRrQDS2Uft+We6rnenzeJZvlx1LKEnaGMQ/lO
9lCPHPjMrVBvMZbpwmUh4ghH9x0DWKt9qthBfECFbfaWicbH2RLweGlCrWh/1JKk
DIF5pRwewWIH41POB3UfSEjGXGyBfVO00cJrXMEfFRcpeQy0bgF4quG59+aAawBR
nrLnc9IbbK3rM5zlVtwDnm0tnbJgV55/R/hzlg+u1hUuxT+zVtM8oD88hh1xPOBE
nEcijTiCS+ykSSS6XSuilXgJgybIliLEzO7dlR+iIpuv/3PwnRYV5ZcpA0qfE7DP
8kDqrFK2jskzx76+GJlWpVOzTvM27pjzuddhiXGYn1aePXF90NbYdpOBeokqk202
1wlCR1IPtOLyUwH7JcB/UodjCTSfIok8dE1qWPZP9HoTJqRFzntPbM5enod4uQLR
G2grJfODzo9emViRH0BGKyWSMIjf258do7OEKZsesioeF7FHkdG2bV7uM6o2ZPKR
qZNau05w4dbOl9pWWuXSMKWckg92VdujoT+OBhCWU1rCUoeQuytH/TzBHoD32jdt
VFmxwDiax0P+ZiLBRqb+Q+x3GnZ8frcquiN30ef9lQ9PDc5PmfXzf4jJhMnVzCmb
e0Sb8SeH1QyS6FVujogzSLQMF7b6mGY30X/NSS3JZvXtOrlLGGrwcT//DKnaBbhr
6qoOLRbFY20YOayG26Ei602o+kWIY7As3IVntruPOaxKcS6KAh9guCvLmx4ttT43
vQ/zxTqNB3SFCbIZddNrxOt16sebLjPcaFKnoHYIKVzk5KpvHgaOC9EHuiavnUkc
XzCwG1PgV/mvjXqOTIwoh2pLsSAfHOYdxSh62lyklc4A1OVU9AMkAM//b4zrzDz6
FLXEDlr7RRpX/tEi6J3xDS+Gv0hHCry+ncaw3ih+udAmyIkUUtZVU6S4SmUCXBMn
iWxMc7fqIdn3jX8QsKEmyg8yttOMe7r05AqwwQaONiCIBIAg6GsTNfkUsur0Nzte
y7GtnAxRI6Wg4TtwtGw/dMlPJ4TMkhUsrYmx2/azSm46WKGVUel36pgJ40Gw1YeA
dwnErla5iiaYBt1txhdJuC/xajVg21gF1w8sxIsDj+TNgKbtHdlFjZqLsxZRwltA
+eq2d7mN+r7tirq/cHv2BbV0S5pGQBdLqS0v1foogKdDeXvpw6KcQrz0frM8AQPr
o8wAiU3KQ+vTQQiVcbzIXCuY/zExcY6Y3OJIXyXCq6v0IDl1KsQWqRJqwhA/OYu6
YqN81QNjyeBAAzeoEmKvJxE/T3pYXSmHGDG6y0lvwdrNZbL3ITb6wGsbV3O2kiGb
8nsIsnvCdOso+jL3mHjiy15i3PGguyfHkRlMbOY9CU8uDn4cjpNqcOi8tq1Qca/A
pNDylYk/CsUXLbN3Q3nrJAygbLgyY79rPvZTwL3382ZAXO62RqLEyqGDadw9B1/7
/kDk7UlfNTBrmr/2h3HClkoKZyCJDY8f/NDQJfiSC5bz8yn1rToxQ73s7FKItnhv
g2hVo6VBo0G3zka68cSUrCSVioFvvnyZTzArbKFh3R5s2co7thXmJ5d02vY4uvnM
7hip4YLUtgW3wuTO/Zn4X4AtjPuT6PFKbaNmzNabGCSsMn/DU8d2lYkzNfqPT+h7
T/tOBkYLLP5KLl/0Lh993yDITu7Y3ZAfI0EDgd1vNhlh8EjreyPw8S+V1+UlaWok
3hke7ngTb/+gkyNnX1dj6MbhbBOgtzi53QFr9Mj/fjRTfdlP6qEx6GyLJKk8xA8A
lntXAocOJsUm5BUr4GouiSusZkvEBJjG54FYMjyWoKx0SDht/Q6bAXZOYC6JwOeA
xchVqWanmJehQVxls6vX3TPgC6U52oga2A0i9AUEGjdnu62e6zizS2yoCZ+zcHYh
yastkHC+e+fQPhtD8JtUWcjyc4aSduSuSOhfHy4h3OSsrNc1iOGAWmfvjTSAm/zk
e+XSbp05QUEjughcD6GZWUkvGfDCYPRjg5uwX27RodSSAGiI2KcL4KQKi6HG7Mhg
tUR4XMAmlKnMVpMQ9oytFPPzJHyohxA5RLGfmi8eAzbL5HyE2sx75XKqfjnUsgra
BAt7/T6AaCuzeANNH13ShDCwDidbksGnRNMTj0awa9qy4bWbX2+dgHvtOf/xSav+
SAM0Ha3bTDDorQmuFYSFTahIiYaXpBPl52A2fe7WNxPe38J+I+J73aFais5xEywf
15bDh5n8WYSZEsQOHHVfAZAggr6eZByy0Jtcvf4mdMreJbhRNsT40C3dSSUkBq5J
hBy/eKluQ2Z7B2+iM44gzMXusU8E4JMgFr3i4xme/hKSl1ME6Iyyttq7Uy+foUdk
VmcDe2/mBCRxX6hLjMqAApvALXmFRSj//G0mTz6DcIeoWBGOt1ylQ2KxSmOldTqR
DQtRgMcYBk66dk7UT3IVxK+A+TR98WR9Z7EGZpr57sLPqjRWo4OkFmr/Zj/DYTfj
FNZxPnUkuHmV99quyo4Kjet67GKuRqrKD7AR5Y9WmiHPMA5z5Pwesb/ahda8eEM9
s3O+3jy2m+Rmguse+LYEVD/vPLebLpp7xk43oIe4exZQMFeTo+l/B5GXMUbkghTT
v7EJq//7/LIEYAyWXXkzDSgequ10MEUjm39Pm/53OheWyjGfWYdKyF97EyFzWJ3N
vCHBgiQ0YyL7ZB7nNRLa0VDNij985d05fiGySC9f7O8ZkCUq66dQx14pUeaGB+SI
y2E6OxIqTG8qOY3seYyr88Ga1r2V25pzO4MqTeYCz6P5GCS+Wb6KToT+i5+mpXfn
bXO7nrIQHryiNNkr/ZCx5uAZcvP6tTbklLhya0wXOPuqPgoToBuiAnfwW23547WZ
xp7VWXegPgMNCB4QAzapjE6lYSHbA2QTd+9AP2ELLXWEYexK4l4PW7muv828I4Jc
a+g8shJY7UUFujHD+bRCh784CFjzuiyCrL/h3JOsznqozOW2fNQqKSE2XM1kUvML
Tg5Rjp3rgbmfdFjCbvjHyMsP27IHLxyNQEDiAoGbXr9lh6pydg4yE4IlSSGbwoD9
Zw1W9qKaeH19LnCL9kL0CArzlH1unpycDu+D+wxqoJNoVrNt9Nu2KzFyDm+f+J5R
XLpRBhRWsUVBjiOjAQLlpPi9yDKozg7fUCJiungIOMq9GLBdDVzS85qAfOvYuqI0
W2YJTTo9qLkivKAlwYQDGdPISBqfsrXeFpxNHJ47YNpIwSkRv2wbQQO+L8Qxr4Ar
PbitZ4H/XiSArCjlFanSijbWDLIYEG0BEV1XiKZyLzgeKS6t96c6ctYVD3hZR8yO
VKWL25fKDoGwn7ZAUUEFmV4sh075t9CzYe+2Sod4wXyrl9fgdAGI17liDp388G6L
2CY2rAMRG4dFH1ooaCFYbpR4Ah7LYy5ODpokHxwSolzdz1rXBehq9LXQxgNEgWSj
P32vUgANujMBscbSH1hzTCBwPIcSy6iVvF0FjH+hSdtPQHWMI9UvP9QStK2IuC2e
Z2kdH562EM23KFDtbJfIViX04+OUwQ9A9i/8aPdSAOktemvRGZIbTJCyVFDEFXgL
SP1ZAsvInaKbLpjSGFe135JF4DvxhUMTpNYXLKk6BZj8AM//vokDkun8kTo9jXMK
8REfWEMqYb5MJAoOqYIOgirMr+P8xF1ZzRrCfSQQv5w3g3uxGzgCZ5OEkvyv0d1Z
3qYwB91trePPtSrXSFeLDuGWwdkbvEFLBjsKsF9OGbOicGntbKm/b6IHV62XoX5f
S8MMDUdsCYYmeclbdpio0TNmpN0dwy3DKHVywUspx3b/VrlU0n12/jjkYO9WypGV
Bf1yCyJ0offfBhK86fyF6brN3VJ4IgVTSTw0N6bNasPGapVOydsW73oNowkUmIV6
NGiLEZ1hxHqMkYEwUR93IEP6Khd+ivPWb02RVjQkdN0KgLKysUW0yPOnhhYY3Jiq
i6REB8BZgdv/YW37JJpBfLlYLtHN4WqvBaRLzoglyuWizp7QNMLoXsKY0ETZh1Bp
NtpMcf0l4+kmFFEBBdvo1S+3QaZHDKgb7FZ3tCcfvCwDJ8wgqukb4MqLGSWy9el+
ehpZQEhebiF83TVTB8Rnx8Ci02/JZ6yeE1snpyUSNrwIQEF4cHiGGYwHDqN4h9vg
c6Oss6BbyFQbJruwssIsPNnBwyqY2IAL39IB5S5EW2x6gtyM06afUqfnaf1NXxdo
czdreAnJGEIPkKazo3GA2D4PmcQIGyxj75k8HCh3GdA8bjkIcGQbhi0NUuQjRpdH
4D9D0nHovmGsTe1KRpfWsPrOCbJS9NRArTE/Mm20HDtuxntKAz2sVeuBJvDTkXOz
zgwH+bXl6tnkUxmzfqCxvz9fur83W4u85owyeIk+VeD5mc978azRlDG2e5OMFJe+
gtG4Hd80VyKSD3OlKsljf9ec8Chq/5vQ38iTZGIF/yGccZ8TJWAm0+LCC+ZKOo7U
NMyvEwCJDpFy0csPVcTXQgjHPopmRd56/Jh1+btbDTLGDhivX/xqqxoC1lTHEq+O
01/rBqMROIEF3XthBrhzUhWDrqoMp75s8nxEF8jcBVpOAaHk3xhGad3N0moFC6Ab
PwpH78+xR0XVcqDFezgU2mgY/CLk+3LD4SCCNKTz1lAukRJn/zhXTqPhNQi6D9l1
V3224N+D0XKeJUvzotiqTI200uMiWDZnZVIu8WNJtof38UymgXL1MUihQleMCXsZ
uUNVB3HgaRpL5CnY7F5I5HiEVjxwboTzKk+TyZegzco3U5sh7o8eqW3Kc+g6xB7R
RzJSqnPGVIqUHxZtwGfrFaPjrQ/JwBl/8+4/WilnPDiDrPz6WFhpzk2mebzcQ/ay
LbixgzmmaxGvddOTpFhM2fMa6AhIZf99kR4SRgK9dvjhaSi0lkWWff5zeKTpsQ8l
M54jl2BI5U6kdX0xhhMm4zMsGoG5x065KNsdj7sVPT8M8z1Y5CSH67pLIkXeaH+w
3las5qzDzQKYIkb9S+wvYTPEW4mM4zcPHec3aoNfee8v1x/kQfsMXNH//m+Yrxcc
SM3p+sORnsyg71FbGjSX7CXECVMm0oG6Lmatg+JeR9GZR9wMMin8eJ+hx+CFduea
0CSDmHZXFZbwSXSXpPexh44qfDqHdVaL2vuQOi+aHt8ivQoOqc/5eL7cnZW17eCH
9Da5j8H/RSPlKY4VUhakJwR4/nHD/53O7lLNqXd3oA0GCy3tjdRoBMNDj7Zm4fsy
CkoL8277um/XRnGwTM26UwCGTQRMvBHBH7Shf5zrNpS/ep1xraCzIAMAzJ5p/Qpf
jQpOPQGL9Bg6tLzxvDQ955FaCxK1Qf6rtsXypRfHiPvOL5HlrI12YMQGeqbNSv3B
bT5XKmuwa6ONPt+0KZsb8KM6LtThmpXCmvwd7YBKWRuKTDVt34XszkI2/YAxxNyt
m3HyLmkOovwzGyhantnN/LaX4L+Tmy8kkX1s3CRx8YWuI2f1U7SNyEyR84bYMIPB
YnGg9hf8YybbNwtNtJdovU3K9EQT4kPgW0YrL2tO31HHmp7pmfLQ8KyRBhi0RBNz
oSQQK9r0V1EC8DW60AN2koPADCwDFROKj/uHZC4xb9gbFusQHATcwyrw/fVIl2Tf
tO/S0Gbp763mtcOIeMTl4hJdAcFlASdIAfQ05MUYi36pUX5qsN4q2yeCk2ZCLRYy
wBP2qfAAPeLaZ8cEacL0feh/bahZ10R9n4oMMBHDiNsrt/6KdeUdL38ARsYkn0NJ
z+szNWml81wIA4vK4GYz8Dy1tAZ52+EKQ6xHO5Z/JBBboKGDI6NOAvGY3IcEwcvU
YA5lZ8lIdEK+OWV+z2xKBuMWV56QxOhTi95uwcSY2qbhIdPNOtnm63zE6aKSfwDJ
bxfO51XBv5DbEwrmqIDki2rVC/PflSeawZSwOZJSdn6i1Q3fKdClC27AaHRED6w5
hGQICuxVJuJl+ssxByfQsfJvyM+mVJWwcmNbz4hxacZz9QuG9mcQJ0ZFmVgLxPdX
hDkt4OixGEViSBjWaR5Cj8Q3xwu6epWkQDsha7TiuQiZfsJAaDEas9DHYLV3UnO0
ob7JG5jmReE3wlTHHuURQFypdeCM744idU+ommlki/FfQdZqoYFWkYqyYaeeqEMs
B9e/bmA+uxNJAXQo2VKvdnKR1CGtGH6FCJ3JqCiam7awWSrAlhGV/jaWrRlF7Gfo
iyrx/m2hz0zjA6CmsbGoytX3rkLgQLbYfJ9/XTt5TzV6Kyt8P6b6LNwZS+q7h4dc
7/RwpVz6UXcQQPsVDgh2jgh/3rXnxaCgGVRUbuptXI+Mimjdh8/t7tcNXF5YcOBz
GwF/erVyBz2GcpaA73PcUAA54Ggtkud9VQSQgcn3k62boInJg+zqcR20QBPz0EPx
Lu9qTAbg0H3Fwc34RzrWnV+DFqTODeYDzwqmRoq3O0YX1gDXS5oyVpP6/AJmJ2/T
W11b/u5Et5604DMcN8vSw05uBth+h23oZ4ZaMtKcReIDzdXrRCnJGjxDBkdVmDoX
jwK9AD+71II9LIkotfbWBgaYa1fIv/Q3WOkmx77erS8uLvnDIq7jn6QVlqateUR8
I8KSX/TM/w2CWiOWMqnw//oNWIZtyHZ2IJ2IqHaVkU8NWl3m7+Wjx/0VHlJcgFsM
6KBR+ugq0+kv5/nd00x0isrLo3rZWCLd1L9fQPqIjmNf5E053mhvzr5uTro7Rgjw
XGO1bWrjdDyx91955zSFT74qWvjKtNbtVzXa6qJpDDt0VigkCDAwm7M47LlTdaKV
tslxgYj1s27N9tLCpmnrSuXXAT3WsO33uh6SxE4yJ3/ntiBm1uIXA9MhzSysbIgL
HdidvhwQfOXhVGmynU44Iie78vRp8qsrrdV83+oU3gbPj0ha/WKyUrkAndFH6VgJ
eR7boXtg3iMhV3eDAubbWxQf6aQWPHYnyda15vzyk9ImPXi8OuVut/4Q20UINtb4
n1z0qKPoahnhWubHENe5HfUQMiipEXNI0HpwCcgrOS5lXZz7AFv7LBDnI6ZUF3ZE
WnhlrD2f8TNaz5XDodb3xp4Or7RKfxRFx3Xwm2fVAVZoOEJqabeFNxljBh0bs8/M
vuQ43dQ3daWJFj/rEeKuJBK33TnsQbEoBE62Txf1MVJfndFkTQnu6XsGJQW1iPxU
xZM1jBqR73Sc1E2Jd6/79Mgj++qZOd/FaL+lI2CQJwZ2ZlF3XICvM1dyQWC34SdO
zaOkqeBW6UvSyi7JoNPvLQFqBzN5xIv/Uf1KgBajp3wdGI3dLTfwUAfrs+GUk9DT
bcwqhhmrX5ykDWDC8UwssJKfmpwmO/RBiLRhTZmk2T2Kj2wGg4bjQwH1/r8P2vZj
0xg5nD7LBE0/mH9kazapy1F3LfCEDGC8lwXCKfR5Zi4Rx9EpXSBU2EoAWwVcQ8F5
H9J2WvklICb7eZ98UTNKNqhe94CW1O6uF8as4vMXYCCBwvnw9das6z6uC1IU8uSZ
mx1n/nhwHiViL8xKgvu1eMqLMqPOq7R97iezGVLhCtDn/+le+bO1rO7D0PaVazfe
x6haxQ7wJX8Ebdy9wpXwkpYYjQRYOucEPk7jYxbeHYxyxNBqQ5bcTS/Zwx6hG6DF
miIAF1TjCQdmeICbyvuIIq1i4ZDE70/Z95XQ6d4kTSqOmBFu5kynHLTNRZfZlAdv
Rn5PxLHxTN9upu0PGeJwublGaXUZCjy+3x3pfGsqEXzxAYM/VjKeouGR+xSc1fsK
o0xzf1eY7RTzn5vmZ8+FJx87ykAnt1hHnax3r/AQqSkS4sTlBIHicEGv/h5X3QFr
iw0SkliYjJdMTff3VXT/DeV7AzgPpYWvrJsQJHzkXR3ngXNnokYbRUCNBS9JnLTZ
JzD9nAA387ghauSGfO/Ks78xH0qhDzylzaX0cP68nLUX8cl0qcIqZ5kV7QlR9qcA
9ivJs2uPLD7yMkIoKRn/NwpvCHw5X4mJrfqakqCUZnupo1x/0j4WWvDdYoNR+c0h
FpTxYEqM+SDCSBHBC4Njx5OkUAOvRdVbcsZm9xEx8kF0kmEwoblKqVrI9num31bw
IiCXpsDLTebHtl5ChMTjk/lIWZFe3kkV2fRCliI3yOOEAAS+aZ7diWv8TnrRnLhk
LE90kL1F2fCmfe+gD3MGkDif81+PCAKPOypGHMIzdbvOX0E/uE6khCZrvtmiIrJs
ChZBpviM6SnFdzierfOD0czzkUrWO7Fk84broiFRgcZxgAeIdrWegThxvpRJuGyq
9JLpdY8l/MKLAzFQeqHfQPIL+QZLrVvIi8bChQbrRrZy/RD3lLQo6CJs/pgrCxrD
NV+Q+vhwCONmssrqhaOTkPpILk+1LXQC2RsHoj53DZYg7kPzlj3EsBUmmNLM/czK
mkwKVjy0izrtP7GxEoKpaC8czAwKe/g59LJlsc0fea01nhEjsqiGQMnucC2RVVg8
HZgkDQUiTw1XDcITEQlqca0DVBdv8lugaG/FloFcW+AzMSfT1mccxhqLKHV3NuLx
VECMiA5GgOD9a9hcYT+e0tK88M7drNOHtHQJTS3cTxtLaOig4BjZm8xKPgdVIXTR
JoG1mF8o2OO8ROLB1JTc8RI1CvB73KzUpN819Ds/NrYDJ79/Z8gJFY4Pn+LCO4E2
bY3QGleHEhe/KVmVUNgg8TBspWWBaklBR57LJXBQXJQ4z8ppAyhSrCcOixRHCKET
RwA03nOItPI5S0LgwmsoIhdPAdQeIry7A2zFKQH8k9TSxd7/HkLJZdDF/Lzr7x/r
ahqTBRlHyJk81dkfasCaRcObVQ5tENrSP/2G71mF4kD2TL4+p9dS5ikrwIKTi3rm
G40a/ErgOy45UBIIAoXbO0hu+M1u4vsN4sMxp1vLvFrJXDwwQxBIsQKFlTgrFAO3
/K20b7SXzkemUA77tvqKKCO0bR61+k1Dn2k9/m+Udid4l1A30izUxUUjd5s6eVGx
guhJKBKCu8ATnwoldueePttKAqvIW8uIloCF2uikPJZjfyhpwQwFOG4USacm72h8
i8HwWXDcXbO4SYHIFz0kZSN9IygIlywu2qQXOz2Zt1k2vHLxxtUsP2RXBZPMXZjg
HdpYFEt1JB4KJk2TXMWGI2VSo25Vp89DvmjRhAuJ2rQOuGaE5Aiht22JgQJq46t2
sXCpcsqJ9WIl5D4ckyZPTkbE23lzI/m2j/yTXnkGTe0tgx3y759bBFZg+gapK+kU
CoZyoBYF4KyGI+6udhKA+ci5v1Fh5UOF0cAVXjZcDpKF0+rosr1OmSlxVptyRy1R
IgVWowGjX0mIh4pHgLI2O9KD7Znyn6dT5flsVBZrrdMvemwGpmgmeGRAABpGVHG7
xr6bvGBxibHsUuuXYtEVB0krcR7WgGrCDJas0nhTm8lpUW+6KUVi2NGhhi27cfYU
BkBkO9WX5hsAyE/uqBKBWgPTNvOjn7kv1PdqgEM/ZkmjAUHNz4iRKR1Xx8iXc2ZQ
7Vv+MPECGrtEqACfhF8xtn5cyvjoke+DY2Qdd2747vMCW0kxT5QR79bHO80zCCtQ
bGOLjuuDLrRXkhfUnhLyczVxbOQf4CSDvnYU53N4vCQBakoI15d279QOzi2mLdzj
GYkywq/08MPelRihANpWlfsA2xxr2/hLGhzY4SxpEKytDf4DXp2kd4xtQbT7yOmw
aQHlg+bvHbWlkTnxbnORwwETMLnCH86Y3BtPKRYffEYRyd4D6fSPJIj6PdDfzVc1
YPdYU8tJ40Tw5OBELkMMfeBGIQZ9scGQAFLh5P9AEoOBGsu6oByi30I2DTaITifz
jPnt+nM+hDb3nWmFtfx+ZFZaMphdd+350dXl+9nnAUmEvYdFbxcchVEWGhem+GNw
V8unNRaNVpGYsLvynW8kb3+MgrlWF5m2QbevN01IwSKLnNBq5WVxpasvR8qeF7q9
7fLi3wcd0q97BM3fmznEbJvvymCDt6Ymt60OQraOu1INreLjjCiQTaBTdg6EBTX1
W4G6uPF1x6gG4q2tzi7PG1YSxKk3VDF3GVnXRJbu6q0vqi/XaV6+/ZkoKy8GjBxb
DBJzduM0QTOZniYaZM24hsZU9jSE2yJn3WkRxXB0PKD6RHvyV66fOuP92e0YqCGA
eijToMAKBR0jjrgJ9XAzDyqwOw0AyY4sZ8fMFyMBWZcMLMSnGmmL1ct285Ui2WmO
xtnTyjnWRQCkaB76tkg8h4Z9HANODX3Rh2yogzxLjErMDK2EUBf5qd6aruQpyMpV
u+QSZeSf85sE10k1SSwLCvVMvP1ZED6EitnXYF5dzpQXHfhrRuPxHjtLGTko8rhD
Q/E5y+8OP0Or9PCk+Svmw8KZkubTcJOa1qat7r8CUeg3ffpMjBAD5YYXTZFr23JF
GTVd095x/MBW/qFl1bew8Q/f/gzTv9EPcxxLswfZ/cMboBNbKVOkWUfcu/inxxp1
zsRIqrMJID9CxHI2xS+LY2WvrshoVo2a/3Ibm+QDLK4Cfx/Q06IoYU+R7YvHZBZ2
Z2jqCKe+wk1NLyc+nYMnNWMMQa/HIgM606CcTeZu1LyfiV9M/eb/kkZk3Sm99KvA
X5l1llyoMUqhyjhgAHL3ZvGHfUzoJmbaDPj5tfMFJLYsfEB8fcr/WNjaGyW2Z6RY
PhNv3mam309Dony+SWo3+ezQc/vXZLIbC11yrQl0ft4t+OADT98/rsA/Qqc44ZoR
VrquhuxLm61azflixjaQrbB4sIJo0Y5b9Ces8Rd9uAl3sJh8dBVkZvSc/DNFI4CE
UpPSFICgDW1w2Zw1S8DZgMKXeNezd8J6ZzXKAr0oLrlubmR6onbQ48FSCutsYZKu
wSZZ0TEsDh7IQMOdhEgC1Oe0SrgKXulfA9pj5HytdlfzxCQnWQ1IHr2uQpje+fES
QKFrsTlp42HQUD4RI049QUojoik3eerUeevySuF53dNU4PZv8U+F/9F7VbgYhT3e
S6I9o0WrN0jdbYzo1/735zoG8jRxqiisCjW/HsaD+55TrEEz90TW415FCTxSozlJ
3QRa2vdxKTniHyDJY8eS9kEpo2u6KNEf03PqGDDiyD1K6dY2VSydUVXxsIyEnY0t
XQKzuaDYraMUH8POsiocnK6bMyKlqQ9D4FY7nDw+7fygIz2IMRkVaFLTIBzyIS8w
ZCyluk7fClftBZ3hhR73nJ0wTxoe2hGkPsYwanJJyyRgBsqkIBf4sBATctLYB/jn
q8BHpaiNnMU90OUeX9KsFzvjmET6tZs5AbuyvfxsNZdhEOZ2aoAXrNDW0FXsge8k
sfFz977Ves/gSaabYWuHkBUvLzrGQo9XjIClAZtVNhCp8w5lbUgBUgk5u+lBqxDP
zU68jt4cPm0xuyutb58H7r9CBJ/D1m8a9FpOvuQES6QqrH5mX4GEE1DHl+pr38Sw
QRVbHykAK7J1x/0TgssERlRhjGnuMEnm4c1NakVne76t84hBjOGRIB2R1qGOc8Rn
jNovz83fjJxwb9L0Q387Oq2hTGFTtlMivP4DhisdvqjYb3mHZ0oBxXcJfCRgltxa
k9lvkq/i1gX9g8QKDkb2wy+dZF3eLvBWN3wF86dfCMSAhTfrrznBPpiW3lhIR+bc
0e3ZR9l7C1PKACeENObM99rnKViFMIcIe3R5fWhdXh6FxbDVow/vGVw/ITCDlG2T
xkAw8mmPzavAc74Tb1WyXbTiHj4GL3T1dFUQOpHk9MXqAjfOCgQkPSBqdnMNj426
JTFIUZUMD2UuYrjB8Vt/3C//M85oKhO8IcRSkzyUA/AudklpP2tYP9ag+X7JNFaO
lTf5Vmu4y7pvYGj574er7bo8kJunXorDgmu1wm7bWjV6vw7G5anWJNHWEfE6AHEx
GgxykKOdWdZjaj5hmm/NtVrmh07YdkBMKTdLIUqzqhRE0oxVgKWIu9uesQlRscZe
+WuPzYFRW0lpg37/XHF946z5vpHrgdP+YbJa7E6GMwcg3qegpbM4xDMkRwTN7A4e
RKy/XjWf13c3LB+eGatxiFbquTW76TWj4d7WyM+RSJntdDeja/B5PghGPlvw7NCT
BOAJla8lSTWV+SWEwAPQbVBTiT7Ga7T7jgCDZ5BK7qRS1HNjpsLKS68gCOVT0/32
LOMPC03yipRxqZpFmueSOVDRsnW9fE5WgtdlEYcqnle6dkYTrl5He5SHV30LV13E
HBFK1lMF6FaOnFAwbTyDBe2N/6oAFOmb3pKU2C80nZfMIXZt8yYERpBsl8dcLTCx
AakTuOmbFd2nTOa3r9Ttl+GIRy3mdzqpPoYgtXhy/GwyJ3wvbM7LgPpBON3ZOl4I
c+PVOYR6jqycG6+/91Lkx1RpEaksRYILAxmBdLKEWq3pj/E3bzcCt5BAvBtkgXe6
DYjYzCYYEzeMjqZK9NGmczz72bdvtzELMOzXCh6hvVQtS8pFVsHE9DETwrezNfwB
S3YlsT4rFx9nXTahG85taocBy+ycnKeIr9+RB+4lXtbYYrTcaLzIVh4/CF9cK9k1
2LTbDA0ujxwVonoByXE6QHRDxvY3w0SOp6cXqSqmQahtp1IO7o3U6TktCKqW6i04
mHYqoALSFavcVYdfcma3K5l3CvR9OLn5KZgdbpWRtpyQfCu0v5oyc4fRXzA6ML5/
v3hhZDWIc5kTDpo6Ty1GCmdlONNHMTudJ7XQPI2yxZr2ZXUuidg/WTamQu2omtWA
3I4fTiyeMKjuKqTi1GNZvRd47u6S7c8N+d4O/xtsMkohwLfhjK93J+bDLV6q1h+U
pD1mnKh2DG0NG5/ONv4E4I8HNpVFCkiXfVDHyJQCgwaISAxPHgVradQ+D5R2apui
BL6n1kf5ehhoX1qaaQHJ+tysYgJsTvdREWp4xAMhp2Q0htNyYoVUmwuoX6l7Sk01
OfZG4I/vykBJ3vZXA0Ar8aCtXoAh3eWaeKbRcNldzTGXqcfEd/L3ewx/9L6cm3YX
v1iAoeptZ7XvLA7kEjq9ZW7d2fHasdR93iZrfFPC87mkYMCG6HU3mG/REn1w7xws
MKm/PHLnDHWhHwTCZqNz7AgutH5fZURGZ9oSGp0CWra+X4TS8hRKDfQ3Qc8/1DIJ
BQv7npGTk8S4X2Do+Q9btyqnFxQBlHYhEPyZMPojcsggbrBtvVUD5PsvlHiWmLsu
9QmGrNoVhjpVFuRiKbTvAWLBgIJ0YXpVcOrbYAwrf18pMo/8AJTiVTnXIJvaggIl
ZCK27FXaI2jvbMPwlZtvKnCJ8DoBCG7vG3l84g9752pbY4Kuwbr/+Eo+rB0dd7Yc
DyZIuZx7r/fJSQoDKqamHTOOnVgK8Vf5RCbolsRJUxnIg4DKVfGDn72d+f9oA/7C
ZsFXwNckG+9Hwv+QO+DBuBQLgr7PrP+fYd93eKFykB6SpiM9e3aQPswczHLBsqsb
spmu72L5EeypjnNqsikM6pMkpstqRNLYpkaJXWn3fzTSVRpouqMo+Sh2+x3ep7bG
26u8Am6hgDDlSyNBCsXVZZLT1zjeJqo2mTtvMR5SyGYGQve/ePk/0AqWkQuenTfE
nEHXqpngRGlo8mIs76Rni6KQsJogvlgYRPCCRI9pUD5eRjzGrVp5J3hoFSUgpvZk
k0KoQfOR6M4zce+slm+PMhVGnEb4GZwj36ZlSTOO+MS346SdfhDzek2mSdpYIkZz
+gxPLZ1VkoZgPlFK3Yi4oOwrTT6YW9hg+E+1CBj7ta6AYPI4pkWdHxN5ec3IatzX
BUWBkxUsuiz2iZQTW+SrNjHvtpKCuHDFl9/EEp9USebl/JpmJA18GURs1lYRgEB1
JtyRG6DA3WbTsMz7NBq7BwJPRldO52xh/FRiazTOKaYRDn1+UYCuA3Ulw7fV3FnZ
bs1XJIeoXGZQCjs8yjjNcIrM6wBGl+Gd3SzjK29rEh3niULl5rwUDp7wQOuqWau2
YLDF144+EhuoSBq0jmXq983rxbq9/OX9jD7DKpqxx7s+KO4oMi0HNrnklBYM4BBd
euQCzcElyiyY8xtY0MGHRDPkSwEDM0PL15eCeV5UChSiKPYMTFoVRBc7EUp/vDB5
urT7gUFUsHynPAkyf/4Axhqt+Q6MhWls8WzgMCqP2Wk5OYiP9z+45I34/C4Vsz4m
ia9G+S2iiB97VNOXdq4GkYlVdRlRJ5rqqPC7PNr08FBy974aX2W7v7mEVTEaDz80
+RlDox9jFptZaCDoP3gscY43ADjIgpH0V0t3lgc63bEdwprwTqv4BaKkB4gK7RPd
V2c/QkN9+Odw3XP+WFlP2Xsgwcaxs5P0qXJgQX1jKY+02hWErArajkfsyUcYyKIa
4K4QH/EsnTFg/24a4LKAHvE5HPilixEERSCQlHsgNWjOKwi9N68amniY08N6nwYL
p0VsXhnkAgNpYK3pqUIJ9WvmeB6MzZ1P2K7np5QFRc7SNZy1P9qzq0CFEV2DkR+y
b2JKamBObWyH2hdXGS8iOantcJQeX9uAQwda0MSOmKRmkSaOOaN8nsI+knT1gmpR
obgb/hIfM9cofhN3r7Pqwa1XC9NDsNk1nHbURB2q/dvVJ7Eed7lqkORUoTtOzotH
dEzhGHBOSiUziqgslTgI4fl0kR0AqZj00PNv+QfcSQ4=
`protect END_PROTECTED
