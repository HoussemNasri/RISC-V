`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HvGY57EJP9CMLgXRLH5hGMRQbSeN6yyocLsP8D7qSr1keW6JaThAUkSJtT7LzjgC
FYAhwx9OXDDlQe6LGFBiUY0xCPXe8OPCLuIW1CqjWJh8/Idv7zM/5dcDvfEScPyZ
28Y/C2UnPjV9uh5NQxXCUTa0jG+FTi3jQbTTxA9gmnIm+xmUr872HDH/U0OMc42g
zmQlAafeK2PLKCHhZ+MYv/+ZyZhG91/tT60Yp7mPkAIBYRrGsHtHCuFJGm1SWNOt
UuvcOpp+bqaR+lVv0ONxiXGlxRl3WokDatBiYI+ByXdz7wD98iONFuDPYRYHhvij
EwRlTA6SYna1gSthPyq15dS2tFxhi7oMGgjT/pLo9Kp7N2EouLxAdzVRLs08fPkB
rDGIKTGmBK1NzI1dO5NOCKiw5tiTpXaKrijTUnPngTN+eDxoldKibq1MAM1Ju1PK
+IQyB2sDfVIUEG9Ou6Jyuu6Sin750LG1qMd7XzI8VwuCw/p7ipw0kuFmfKzxMydH
6oWM2iljElCI0tml+DST7ojIzpWUpfEPYApJ/Ej18aI8pT+m4jqWUL5oFgvADU1N
z9IDyN2XKdOhSSZYW+OO8Dj8ylClC0oJqovoYOeOBuWTQDrFhYmZBfiOLeQt+lLj
LlaZBg8cGES8ZGZiKQTPz6030QhxqBw2lowO8GU/WDxPIPHEVwIWQwfFLTfCvOEo
0WsaOlHtgaP2masOi8AOSRCdXcx+0g3YHQYQQyU6eRPYWwwPBzzcjUqxjzyDr+8l
FR0RT5v+hlhXQfrrfMWut4cX21C+wh1VTq4TfzgZXU4yvM2sj8Do0bqUGuH5Xwy7
gx/aP9lFf3lw6myUbkrfZtj/9qFWlIn5Ouz85SBg++7YvoKxFEzVIV6xaSXtO0L2
zxx0CgIdQAs8Cf6Wk/GrtK1VeSNlIrPaa3Lf5vfthsNId+eCSwADI/BIJ/ConNPK
i9acKN8r9vhuYNVQnM5h7iDfQ+MOkAQu0EOtW5qSeIyjYByVUcMgF1ocDUGhc0Xr
3U6BS+5btLNBnIKUzj+YkCdh7CXRqRek8yJSBjVo6AxlSwO6rsCHG2C8fxlR37oT
kCiNNv1j/NhLTqLZqygyBguxzXzYfxgl4i9xvSPjVGvlgK1n+Lor/RKcHSQYj2Ag
di5cKGJ8ZrSCblFD8EgX0vWGl8m7TDJcslI0TLBlHZSQExo1sTekhxALVi2GYb9n
gU+YBcHXpo2z1+Je/qmy1hHb5JUPNXgEKjxVAWtP2CAe/xJHj/j+x85U0fSMgoXi
isSMYTWwcROw+5X+ugx1eDy9yci9qMfrcsqIzx3vEYVsjvmgHfjLJVUjzE0Nrhkj
u3RuyVJTAceHY7mPUwFJiqNtTilajSbXuM6vxItEAU7/gp/VsemmkCKF8W6f196t
sUASWpMt84bqP1/toFbEzqowsw/3Qn0VwO2RJWgiBiTHvoWcaGz5WvQc5SFXNyBD
0s07PPsoeebyt80SfrTbs5ufXslj3qrmmXVP0waO+E5WIYwfYy1f82ihdtrW1tvh
CSnjT0jmYoY+jLphwB5Nb+43UjVG8TLrnfHMsylhTQXjJFutvHnGJ3VQno/YVaYD
f/eb9SYzg1muCdlNvWVQmSmvNXl95Q+BeEU1cs3lllCI29W/hhhaD/dnZZP4/PGB
MykNaQqI1ZH40dxJ8qZnAU761yr9Vto+IwiwNKFPLQilaEz0D0G0cuqL/BfGJcBC
hjFuGrij9H2//CbDVjp7s7m3WQf6ukXr3S+pekrY2HfuEiN3abnieGm6DQ4pKYYl
`protect END_PROTECTED
