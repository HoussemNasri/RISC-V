`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m8VyulK5/sxjSSstmib0ttsjiJ3lvE45z72PzmcH4H2u90z0Xgri9oQMqh4Wid6A
coVAmpBLKgC5R9XgpNWgRtzRW0HxxH6MdT4sQ6lnYx8En4LNDA3JVwJK6tYPGcuS
ZczQNu/FhyZtXB8ypT27Qgo1EYfrCLETFFBqNlxh7aAIFRDIACK20vWf54NFgIqv
F1NVGAuDVyBKm6uR04znhoY5g0yIwXBzv9YM+bCyJ8XnEG9dLcaSplxYUZQQILQJ
Wm2EgDvINLF91CCHMAsm22+rqGe3k43mJBOXxHxRmuMZML2fqVFqTNvsSCP9LJOZ
NwDwXOplKacKlquF5imj/WueTznwCGSudBEfSFfRNonSIE+tz+604J7jeZkB4YwT
neIcRe9LJn7zEsMfetuNNja87G1i7gyEqjdLG6iWrhyP0Ri568vrM3r6duI5OnSp
C8HQHdaHofH5A3Cn4TLgoEJnkfoMlLFFMrzhsNl/pqw8t+JzrSFppp+h/BptGSb1
P51vtKyZL1M7Nuork8I6QstaPk2N+42YX1p3cRfhUD6NW8YHuO8orZWZNprebAER
Ovq1hJKyD7d47NevvEk8Zx4w4BT7NqaMtCz6w5/JX5I5XVjb6GNygVP1MjKjt/6S
/ofGXgiBGi7L1Fb+F7feNpeCSgNt4j6EQEeD219UDIFw59DuWOSyXiFsyF8DU7y6
2yi8vzEzvbIF0kbiq06ggPxUGyC56pnJOwDWUSFUzHy3NpH/jmD3dFzEMCREPdWm
pg1dhYIVlzPMA7ZVs3dpQK1p/O1EnbMKL8yYHf6aSQqdvYXjR3Lipwjo0A+SQyVS
9oDKKUoa9ITd66liUcKgUhrgtyNsXBkb0lQ3F+D22qrAgebUA7KG6C6SQUzWrMSC
d7cORC3Fj+OOhLi03OdfgnGR2OCzMOJz3iWMdcfnK3gxwE2rQ0PtJQMeSCbjTUuK
us8iJAnSHxtWEwvCPkdghObAyHeQIUjIrQcRGdI9WTQY9MA/85X2IiSAdMrK4el6
IuXDuTfh+8m+oCPlhIR5pkrLJGNji7OOuIrcnQSBtDq1sXBZZ+B/8EPeLXatEh2x
AAkNhGPJ0wFJKGzLGQ8nrnoZYbV9L/y6QDued31hfWi46owxLX2Npq7ByaNBZIdY
QlY8XN2nGUkqE0O4kgDyHtwHxHtV8/LsgR559Jp+fps/7YG7mpLNyf/0fVr9JChl
vL5290lhXxxraAN1HntHKEJFdsylLoy1KAzpWWvqGdMlI4l2a2V154bE1b2SEgqQ
CK8hxSnEMcrkr7JYqxTMTguCv46ePSM2FASUrk+6J5OM4TI2LVFLOSZJXZnfupKA
rCAlgvElYl1mocemMtADiMi5pkTNmFUm2LH5WAUeAxWgeq0Xy7J07NFLnE3Uqx14
kcL04VnoafzWuHiGsf8Y2UnjazcADML6b4N7PVqN3goXMR+/ifaJQ9gZkkT1byfm
plLtxzCHa8GV4mC/G2dZl4LtDtaZsF5ovFHVLGFIsEOHKj87FE8nFA+0xOz44HC1
Qsrk5b88Zuf0QZXP6IDmLXDQmbPjKVJVVSW9yBNj3dSaWGeV2LsK8sh17Kw5WJH/
NVb2V9A/GgeyaYIN/mvxR4/SROgeFG/7IkCyhYMV6uBqsGvucT1ngtPyP7LuO3YC
H6JF0zhwGqxsm9JtRpOLIrsVW5Fd5UBj77eb5oLYBF/i3hxuQeUiAbx7d1fZf63+
v2tifhXoJIWRlhx3BcKU7wMFG2fqpJ2oQJ5Qgh6Q4S+c6lNn4np0Xd8Vd70JFpNU
tOXrLFx0GTLrgitm7tDSG2iOgSZP7x3dL20akAHKin0NOBPErsbIKLZuS5in6mAs
tkkz0AhKohCIYLA7eT14rbCba1Zpb6gmraFQTrePKtCKZ+yuIaZ1H9SXuzBSqXvE
c1vCTot+WYZRNvuf2iFHn6OxPLFD7hGNtnU7QqCLo3cY1KdCFnC5lY7J/CvBu8B2
jgV3FFbdy+YC1S9mNwSokvYNaLgMopRt3nhEaoritE8WKGING6HBVbG6XQIUUdFE
mTa+gmEFJ2W9K2xUb1amLGoe8BmwyMsn59V2XOW9tLHjkDbYEXQgpP/z5u95HK4w
P6okGkYkrRV0RnRNJGo5mYspqK7Sh7psZpofK1gNK4zg9qz+BZpVliTQxNZA4erE
/6LCQxM7qU2w3U1BeYiyHyoqaLgqk38BKlKIlmy5fZRK9ID+RbhdBON7piegnq2R
+I5yiN4LT2SkoBm1kpYkfPeCKgA9pi0VVR6EiqO3MY88ljt2ibMn48eRJgzQydXq
pFcwfWCH9x0zXBACoC8Biu5xpVwwgsoo0tuNZyPOyc7hZ33TkMnvmlllnv9xDTjU
JbKbGHps1pVmmc0Y+lvT5fUCyWKRTfqIOV7pxoSai8XkGtaJylpKPRPI9A2OF4Lr
oeuzoUXt9ZSqFIwt/JYwZEsrF4mYg7f9H2Hmpb2JxBaP3sHypHV5GIoyGGkySgiX
go30MdLYHef4jEvzGnDS/qWV3lbBUItolm7kfkEDkxMzTjSRA59l/N1TsMWLuDUX
SHr/h5Cz0xQxtaywR19RVmz4gz2Pt/bbpYMGyVl6XELXRbHqFyYtD1087xz602Et
pn5c0rfYCgJNQpyYHyu5colm20ncKe6ntCq+U9w4aBuTSR9dIOwRMA1qL93wKxm7
1JG41n8jqzSmNFVANkajSmBvGPMTYthI6HlHz13IXZMkPxjHjGN75oKz5uVbDYCl
YVGC3CWs4WPzjZJKBGfo6XJzlOyjXtSo2z50CYfqs+oGC80SSfwPAqz+q5P8u4w5
rDpSAgSxxc9VZzytcvm27jO9MPqPRK8ecx8aiAEPilsxFO/02BfY6OIgBuJcNEAg
cWsiWeg+l5mFsUFy3HGd9nL2+epeUsIy/AM/+zxDCTUk+PtvvxAApeccI+uCuq6y
xrSj1g0rluo08BiIr23Q2Kr1wc8RjGzvF4JFnLdUmjR2gEzRA8PYO8Bno9J4Ftpw
1c6K5RpnODDKHK36BQWBy1N5ZNDG9StgENui/XqnFaJ4LYmOaaBpJX1B0X6K1c2j
70FM/aD4MXe4wG5wj2KvEQgAnPCfQiJSs2MkYfUkkpEUp+hBCMoZ2QI00lFMfS35
YKVsJf9vy38vEB8p1sTe88wb4lXIWOeZnrFEZg04IytbEHXQnQxI9AgAfKX4Fb4+
fZL0eZSxdhMCTLTZWUiy6bA/pUL7MfRSCB4XphpBi97xEkOMhpZLAe32v9Uuw7ao
Uepwyt5of2XenZKhRDw17F4W6/2ZyypicHw4PIfTLaNX3JO4KrkpoP5IrPf2wBOd
OTxg/Ax/aeJHgZnD7e35f/D8mnvgTUF4/TkPaOIG9P79pSn+BCCnXB69wZcXGhQF
327iNkzFrgsn5R0Xdh9GpQDk/9My1lAaPOxeCMr2QGSttz4yHjg3bQOSgZUpnyUs
D1ZTTF1Ohj25tNNAIksHrMA8Gi6X6ByL6SN4ANs1BOA9lC9Fw6nUxhO6N1nByEBh
t5wUKmeGArNHnTb2BbnUET1VakKbs8V6z6It21UJH5bTAYS0v9uQ/bwoMS6ACDjQ
Jbf/3NqxVs1QyVMZMEWQR6TozgO5uJHHZEiRmISWmswHD0ibqCKAJEJISBlW7Te0
gSGDtVZN/IDZ2H9ulbN7QaKzgOyniEb56oTL/Ajnmv5575rkMg3OEsOR8xo64MVR
8nYLvGcnz8QHqldu9vXhPcyNGd9UjIwru2iCfV53KZKiMRsuVwUhOPbqrPD5Jv0Y
v5KMnDcoEj6P8mHchFjF1GgojQfQCUi6dHzmpQXaDVqQrmNHQYiBMnJB1/6InPvS
wgbaaJOLusjOBhR6PxQNacAw4d6sPYvNqCHCF4fmcoJR2ADN2US3yUFiAL0zAebS
rJWN+VKa9fyWQYPvCfRTfcp0YHOaQ3nICRN8kSu5zoetvT9L+3MEeKgGRi89BHmu
wapcWwlYJ7tx62rNoAmK2HqnVJDI9InjqMMoNesXruPRl+2cSjRMUwXDuh9MZmxH
3Lv1Hi19eBRqMSso3LkFXX8htuLGPJdw09D42GMIPSE3oPN1IbZlH07ShRsomNZG
9DkXXNkEAkJFF9lROZw36u1ArUXJBFVlaHynhTPUTN+GgKHNlUxIPp3opp6Pzjpm
k9QOWY3kwd/v/X8UlyBbaN40XfusA81216K+HO9dy1DnkhIX8iTsmHCtZvcGXd3r
Jh3MgX95DsdDzzEktKxq80+2UwPg0HFsNYFSrlsAi0L5nt2m7h5IfHEVsPG4/lzU
gXkwSIrGNlRXXaER4ZNIoC1I+u0SQscqW+rF5aejXrFBVG7/IXp2e2djrPGgqeHO
NQInxUkaUystIQIXNDMhDzmxXE5wtvQ3JV9roSkvJIBnTUFKCDUjntweD3sqRIOR
H5TWcnB38zkIVaZCJKkjZlH1932a4A0+phZBganvBJErUnAH45sjpU0r89XKUv7o
Yd2VPSmHha4ndypUbjI2YpCuWSM4d0qDQF+8NvSs+GnkqMI6gNv66te1RgdIXCZu
/H2oA3+xhGgn+V0Utx1kOIQAzPJzMjmQRp6zx55pJV+nkcwvqXySAK2iHtqmYdtr
Q+PEFrBxP8Tf5+B5RVXZfAuY/JhgOh8+FDN7wgwPln52IogAz8lsWc+MyqTCSBvf
oGii0cPR2A0+L+GpZ/pp1ElM9VsJRfgC9Bd+hEDNqDLEHLGGVdqEfnZqn8EU/ONH
jVU+UNCy3wh4h1lQkERX0IjpFxuwl05n1D3Nryezvkm9XmHdzCMDte1n+2FMgBlT
juLQ3t61Ar3jolhQfdCTpYfPIXAXzSzfT7RXcAf9HAfVmQucKPsRgTyZYdJXNKen
CcNv2fD9uB6DcOVd9dvbxl0NtZ0tIQi3owkC7RAhBo32Af7TLn+iicB8mTosR7lH
ywWl26zFTlFLTSsdRa/7klr6qcZYhwcM4zGJlF9XvaY/CpQK4yj7+3Be+w6F1F7Z
S1X+4S+gFPqepLy0rkWPsslbM1yVuR8NbTTqyyyYyOs06wqlkiN/9d+c1mRtlZQe
81sHh37xIAu8mKqyyq/6B5RESRq0hv8jnh6IZdv3w6eoKHGcZACrxoL3slDrkBa0
WQSctjjvXXvX7cSvuzaC6UhHiUe3hPKt3Ey9fwY5Gbd1LWy6FIsmJq2hY/EUHbTq
I7tsIM2zYaRU6o+ty2PYWIHxfIkv/c079B5vsbehBW+ad+rjOHoy9X74imy1+qhM
s6ibZQwrcVYN+MXfuuFLyJAnFiamM/+d93zpPW9VUXAF6X/uozsMXUE6bRBdDK/G
X6eC8cpCs5+nt9jz+PdfMzCyLYmF8Nh1+4FZKvVU4X5f/sLMFLccdtAV0ERCc0z9
m7NLJu1aUaowoEFy0YnGRwYQTp3HEK5Gu7TQb9yLfjZPuhet+DbbQ3163iABuT6L
kVucUHeBxnkuuWM5WvdaabYDLw7vIwXpganqcvqjejjYcv/pmtmStsuUNtjeA3v4
c5DYt2ORMMKriTgt+BaYUE3YbXbRM+OvaiT++dxq5DsxqtRoNCsek0OVns9Z3ylh
adTSERU5OInWx9ir2Df7oR3SqGC3tr1W58jOu3PYajtUqsRvOnQ4iiqcdwpUsq6E
NYquCc2RtODtHWL1KuiiSYFXoXwJu6SBm8UwUW8Q4qSXLCK8HImkhRAb8u11qAPC
4Tc1WWRAfmQFgCVVpC7WyNl1mrBkC+Is8SvwJJ6iUdFsEqSQBP47Ovt0oLZj56w9
uGkYUefrHU+kyHVkErg28dU4T3fftPyqzahVRelX2plu888N5//bXtaCepsSaUvb
MKPbzlfiF5Z8nd18+STAiHecrtBvlU220/PlGLwCMRCZtVMKfSWPVOjTbxdApsB7
w0ovKmfOz4f2udJNK7ucUFPrtwnALuM9aVUFLZxPPDYinlJod+D//SW2GiqUQeD5
wL87Dlb1I+XpM+BLu7/Uf9GQFYxLdpyuFhjZHjK+3d9Fx4Zb9GqGWiXLnxpeBEvd
bj1vl10cwxhnd/xPNmgO8iSvKEB2MsT4SKT7jYHR9KvfAV6ZKXxa+dG07h8C0+n7
l7ozqXamIZxBmyf8oXMqujxg4sjR8wKCLhq8IZPB08BkYxCfloqPciPW6T14Fgkt
4nwhI32f5o5hshM9Qyej0b0uIJFQM1fJvROUjsmb/JgMIlu2RXrrzzXE+B/PFJSu
mJ7qL2AYCjhRHRi0yB9O4IQIRhEjnCQ5oZ7ymVNEBYqJI9M/NeiP8mS/vvPffoZN
LwMO4V04FrYdwDucDrXt7qCFWPcSGMOaP5HfyEpRBymY8z23B+LKqqMy+RYeQOQO
07HmAIzYB6pUwTnuVc0jUgYtZiH9Aw6oYYkTDj905wC/NnplsRcWvap6m/umq8XH
drn6deHXQE+zBHlwHvaA/5AbDzxcFiusm6w9zmdb/gMf9hthstuiRnIwGSri9T/D
w0rIhfxDnQRYPZ7goQxuxqB1PO4s/9oSHYwHj8nwGA1++lINiPlQlFwrXZ0j4bF+
dN1LUPhmmtIL3Pp/LOTSpA9zUVvxLufB1FX5JUTHIhWzyzlC+acDBGuiT9LpaK3X
BP52Dnp9YXEc3u7b0qjk2lFIiaMI07dID6q6++mOi1UakR9wHEDeovA/8CweFKlN
950NDYxi2MDaGrFovvgKE1yk0NPZftYT52DXdLRHSifP04E5inlGYIFzN/o+mfSZ
1XHclO/jD6gj8hHevEfXgsX3uypubt+XmelhDAgtUyguYW0/+zAp4VeIOvcRHfHZ
q2hgqd0f5cxBuvH8SAKWyEGlASCV1Gwr49ZTmPsdZNpNLId1NIn2Oc9jCFSme3+2
b7v1tDAjNuNTjzX1GGGd2OHnx1fFefD1iSlHIuZI5INJu53syo2nsM086jhn1NdZ
GJn8jPqCpzxoWUYWeyhXkCmnyS/NtSV/th/KYu6q6TCnW4Mm9wrYInOJnsW5PbjJ
qwiG5VkVgQOGI0IbfmT7JXdhKQxrnLOMZ3pONJDyCrhNFBz4+oPxkXgp/bWzh9aH
frL9ZMLX07CZZlu6lGzw6FeAEQbzGXrsaAAV1Vm9HeA1DKV+FwnpU1Iqr1gWceSx
dPG1ZBwyQ/htlbL6SqomIq5yU51+eX0DYihZuoaEmgPydHdWJ2dTwaetX75j3ox7
dz7q1aRCYrzHg5CnwVJOYJav9bDsOYfkcfcYhkY1VSOjI0aAB2nKj3fAV6Qfo0D8
ZojyeSWK8dQYTPJp6yoVzZFfzM+kgRMF9Xr+K+ZrMPQbKZ3YKF5CMKiECQpW8yJl
XMz0aezVMiq9iHrMTQhfy0Q50lvHyf7aRqOxsA/JwZHJ7Crs4v0ATtJgrnyzb+6Y
mag93WwlhsmXLYq9J8+Sik1qNQ8K8D1+XoRkK4ZX/Cd6c9lwvMovOE3nYdrk9SaT
OqbNcR3eXomi4V33m3Zh6QI0VvEKlcWWwvuZK/c/T+A94+9R8X9GiHeZqybkG23t
7odusMLBo8S3V5HS7ZnHk5HKIxK4dq8v48t+EgwW6QVLbiEtj7iVo92stn2TYUts
ttAgWOqQ2XpEsN1mxySyXefsJ5fkwzkjqcK3yperiovq5FDY4s5IR4ydrLwPAb7X
mVoJ5nk/Z7Ne+KDPViZvxX0iz8POzBcMubUe1gU9pM+fdqapHlUCmsMuCUAt1Q4V
ECJxa7zhLkUJIm9AgUwUpho8BhVM+//bQhNmqstbBCcHyih2GAQe8TTKgiRuNKiT
BeSEK5Q9RmVnQwwK2EEBuJzd8K8Ae4ogm14k6MOJd1Z0NpwpaJmUrKwe+mscsLh1
0t9/7rfEgqkHxjgjrVbVQLtCeue0BmjK4dD2Lr6xzehvQutQEZeTLhXwli15ikRo
rmjxS0o5qWaA57besZFywi4kynxEXrKurjO59qUKeoNY8slzskWVI7nvxm9hf3aZ
Ir3xaaB4CyQ+0vBEK85jyMWFBZu1oFnpsoqvLvr80bCFLlmxGClFfs2X3Nstx52S
pncR8o3LG3HuxNPL0EPm9p6+GoI1RGGZKqgWt0jFpI5tDHZn1N3eoV/1e1dXO9FV
GiClMZFmAjdD3UCEpqIB95i2gIXUEbID7Uq4uMAcodVeyniXOCP2kME9QQI5ZSJe
K/5SI89IiIRk8IrYbEW3pHfq+zM6uB7alKJVFkxPv1bdTlP5TtOVHgpixbNS8oqx
faE71deichWeBnLmbcs3CF8XJT0b7FOgZQdWBpa4kkcZXjZPkqs3CaPzarHMwYtS
2TyJmAxbJR6j/n9uPkQfrAFuQFpGHbVwVOf4fKl8zY0eGdxnkK9mJJWDcKjzwqni
4tJKa4DkxiaZAadQdxTlH/kA9dg4YLNIT9JkylXRcpLtx4U5grQA6Ucs9efMQkXB
AKkivjQShwdZQUZjPMLuOnbhvTGHFsoC+XENU4ltVvlNPQDk/gNTyFxrHSiwXLe/
7+wHhAJLxI5dyEE9CId1ZZylbsfKPRK+qsn/2P1rYBa6YBj9ZhNlGDBOAiHGMyUj
aaYkUOW4NJushisLuVwvXkAyIna+nf6Geg5y8mb9Dpf6uEr2brT08wHOgVUFEjF6
5vYf+DNgf7/KAdrceRk2Hj4YmqowxLa+rGFVxOne/TDHfhvJ+Udn0bGbV7l7E0Cb
ZYKnKP+G6yOtth56IBbglO3GZZB34i53VUgLWWhta+XvSQdHQxWfhAsQ7s41I0zl
SOB/4KASuO/mlxrLtcrgC6DkgUxQKI2tlloddR/e7qBbsPFgu+O33AvlLyZJ6R4Y
jKFG9kJlUbHp2iIlGaB3OV/KsNLKp1wc1U0n1LHB3hefWT1gCb3uO5IBZ5arRYhc
dq4ZaBY6lKIwAqJLkLdI3qN6uvedIwRlaFfFnfXdWwbRBqkEXL9kLyqNFQnau/dm
u22eQDpTbalF0f+Rw1rOrec10MnEpKh6YN+dM9Rju2p9lJwuH8mhCTizp4kWkmoG
Z7rJXEoRF8iNP+ULnri8WDuZltWrgyUxsOGaNVQ0vR5HtLQX7PbaAP56f/AGlvka
yPhewjz2XtjvLVDXHdE6U3F/HtZ7/+6DD3rnxSaZHK4brHZhnKxezXn0bY4FGvbF
SlSq0Ph9ZbpJ7dB32xEdoIR6Un264yMZ18ChPxcwWVEf+xfW1XBmVgT+eRjIsr/J
3Ajj/YVg0d16ZUtcg0YRfcgbIvDAAc7Oi+XR0NQd87+BUc1ieBKI6d3L4ZH8N/qE
TPMekZxTe0CCCD72GSEgV2TRdX00FsRndsAdY04TntWFE9AWqjGeRewPLmqo9Kcw
H2/NHDlCWpfJKHTRGE6xyDklUFQIw5g3tF1XX7r5JacYRtKntXP6hcjEry+tE9Zq
Dsr8w03Gn8CMBDPtQEJ2DRU8kr6MJKBmY9KbxHdE9ip9iMbwz0kmnEwnbd3DR6Jg
eGdvSdoVuCGPO0PxvAZsXJR0G2wqwpAu+hsuS51ulL1jpaxf3GHxduyKICyxUDqP
2S0BxxL/Vm93NCQjEJXy2Ep/RoRU/WJ/MYenV33GHF0+B4XforEp8lMbR3UyBL2d
yQDi5uI74D45v1iqDz6BHMjt4USp9Mvf5I3s/CSXlfEKpAZYl0aTdqu1EPqJHXjI
ulwI307TJWZ6sq9i/SqC+fMhFSXLnMrbWvfa+vBc+tHdsAQ02DPUzst6mB+/HNhH
wWMRv3nsmyCpbQs02ripZKs22QZxlrCz3mta6aL+HZ/up7I3Dn5RyZj8MVnCaPyv
xH/MvvT2XPmooT4LTa7OIpclv5Vkokz/Gfn5EejOaAsf86GkUvSowKM+Qly+ASCz
V2fPk4ByVsQrqHnE4A+6toQxqE4/UflQ5mIODJYQrzVz64qCcQqqqemYenDBWzpO
Wgbxz+vR43hEc8vFtEk5VoaXn6jXtqtW0OgdjvqOBo8eKO/T73eEkgCQXfHCqre7
XMVRDbtkh8tciwYBqAvEfZ2HzN4sGOCqxDZfy1X14I945DoVqFakZADKJlAKr002
Ln1Gu5OMAWyGIhPxY4eOEzKG9YYpKmqtx/EJs+JP4pWtdibvcDiVNVxybv/i+jMW
x+Ra5Ig1AsKHKSor5vZJWKh9APJqwp4jus0mzp2dXsIWK3ib1QkAL1gWxDoSmmtp
6PIAQ8jIfetCcUEwP2ehTEzp5RkjCoKHc8zve3MxzAHHOk8JLvEGiDkPTzMV7MNS
6b5CFdL7Xo9wAH1EfyU+5xKEvRhxKIEb+76eSuI72mKB1qH2aD3HObblZmd82a87
O+zPO6eBNmPN28jGrz7and+VjuUhQdTS3p8Tn6avE0kKOPmu+ejd2uu6fuUh391t
1tq0PcO0nLLYwu2KBrOD7ebL2GE54CnAv9lHhiVM9HuLJSz7v2noA++EK6VvFbd8
/LOcvObV2DKtBo/UT3MDKWNnM4yi0fLpYXDOr60VED2UecZLNVILuPAhrydQxfXa
DKIqE05oxZeCX5cU0kr29fV5sk7dAUuRo0hkHIuNO3y/l4CN179DSjF7WeGTnVV9
peYd+b0sXnem0ZCEAtz+qVBXzBP9dFI4YbPbkjLrdxK3koX4QuBIn4+jKIbLMvg2
xW/8F1X+zwMcVaX3I+iI9Qsw7j02hMOASneNjm/zv03muVJrkrTNk5jrVFrNazPc
TlZLX3grhVpbm9eNi8/ggk1jdtwNnjiuaN7JwnxlnuvMEZrC/5Xj4qtJmkEfSvK/
GAONnvLkIBU6Cm0/vlpVafd/I+EFK6DKptSmhX7IgkeGZbg/StPaQP8msTSaWdMt
2X3Jumob1lLklbtiurr8tvfSlFlNviCmrtETICPjcsH0k9bdhcLbeHzg+zttpIMl
BSyikO7yJrRtnDOdVNwzByuFZAdk4FZxPZpzZCxbHEtMKP5VW37t13qcOjsz+Whw
MLaRy1lF/yTiDt3RoATIQCacdzWkKTaITpkLMlxhPKbGF6G2ZdzscVOLWWW8EAC0
72K+D9F6bEXVZqEkt8Iv6g9jb7RqWLVWoMTtpcEdqd7/G/gkMgvX/GF/eK9eJReU
74wk6IHnZzM91lGaWmII1GJHQuFX4GP1fS9kIC450DEAcJTjPX0mleb10K+bFBdb
q9aVqDj+9YEKsaYaDReqtRMfyLRHg4QYfIl6xh0ZsIa4Zpc9kQ0NoBl2phxrhWgC
qLX+maEuQXLtpss7RPjI8GXEegxD4KLTLsk3rKHDNxoUCJNrIswr+2pvpsDnY1eS
aUbPb113OTQG+7GeVQED30Q0G6nYJccH/KvKGVeQB1iyr+0sTddWRIKSJW+FzJ5d
EL50U0ElBWFGhiwOMQ7R7Cd8z5jrBqfkJ7nkVwrst2TrB4QtG25JiQORrCuS7c07
/RTAdCk2c/90BF5RuHsbvDop/1biVQVImI7cInl47YnPVUXuZMD+sscISYY/Wu+T
sGQsrzoJN36mxah1CO/HpaFU3Ge+Y7t8GFYa4z5mN01qIN0o07rMTIbQGLbYbg6N
PbS2a90nlhHtDR1ibV+Esh3mu1PxiuQAWql7Yh43RcNiu6tgg+dfPacnLVqPROu7
zk9CbCtQg+sVOwqS6F5mA/sdsTrXbRk+Ib3Gw7K+YgUjfkAe3/EVAv1kPTxQxG9/
3Bxe8NToGtQt8mBWUSLaRPCElwfaoRIDF5g94cgSPwWcSRSawUnnEjzb9fZDcjx3
xqrYSOAktz3CSsrD7oNMhLDVcRug028KUD28cJUFpZE4Tmk0LJmZQKhTk53miJA9
b6IFBFONoV5ZlXbSj8Mrypwd9djZCR7xtdrdzZHx5gF5AOmgGt9C8QQ+hHqleGMv
HKtqoOCuzKqGCLk6jIYLFAbC3CudDuQdrC0oqEDscsCf+gncZ8BwbwrEwhx5fCye
gCP+RvxcGIPtTA63bqZwrItjzZ+TaAcT5iFL37cwm+3oJ7fRL9qNgD2f7Xmh5wXe
kRyL3gTT8SLs/v3fKU1FHUlcShtMWUuVe+n8Ahya3oNXr3k0yyAE/9WWquaPvax/
3cyI9LMeh6kkzsVji69Smd8ZEZ1T4Aq/geOlHj7dA6RtprkXQhwyAWqPyAKz32nl
vTQ+sORjLEDnoPRAUOPsXDBhW4N8fZDfliS2/SVfIINVw1TxytGvIKXcLgCGtmij
P8AWupxmRrdHvub+dTuogZaz+B6MK0eKjCH+y1mrM8ZDI7ZHs+s9r4XhmVGRY8vs
PCOHNVB68ZuB647oYWOg6WKDAylAdoP1ZbNoEXFB7+/vbDWhGRGfOf4XXAQhPwkQ
5nEiRSIGyOynUx16BAWJSJMugi9U2R/AdCpbebgEO7lgB1P5lvzxkCn5j8Siq650
KU6rObB7qgKWtsdKGv+SDBcYBJGGBgoY/aSvnGNBUFM7lyfyAD12G5Wp6FvXUHRT
aTAT026ABdaIVB1xQeYNaXL5119RaZNeLDEMI3+nuVHukyBFlLaWP2pEDjiHZHuG
qLiEq2weFLSgnRNTvx0iltyq/PffYdCqjKx6Cbg0m0AyuOmWs028Ei1ZXvNHkZRP
TmE3se+jOV865mlMua6Tw+OKKKOaYGDHaqPH3Aeua4BdMEx+4BLFL/RSa/JoLekV
xE8nrOlVOP5zdpYjxhcKbrADm6EFQheF4JqcGDQPPu3xAFV7dogctvzCpnxyejtZ
FgOMzcOvD3fyVdxg16P1448JkxjDaWH0MrsLqJUuS9jPbTwfJ9/aV8WqhCpsvqpz
Fz+wdz/fqJ0L3a7JEnfxe+7CFScZXCOkj3KyGsojxuFy2iZdT8/nST3NJ0cDo7rN
tUmVPmmCdqS2YAI/4KMRwuRiCII2LYxmCe85xaFOTKx4RYI6m3CoJE5rlfg1bFQc
z43D1IZ7ut7x1L5/z9bKkhia7aoDHov157PxClGbEy93d8UesbJdnwMluYnQkuxn
wuOPU4Oefp/1DMG7At7/gkBwtIX0TXc2rK58zMUOMwqnB9EVCadt5A9MV6rcRYl5
3kKwy3Q1gLkimQt85qJ0qjZK3HKDPspL7nYchqTWHA5J2baOW7MXThQ/fRE8bcQv
t8/yJcmr9hfnpYTqrKOhYrhErHayVIY7G4OqOeWE5ppT6eaHxmchU/Z8hd2/O4gT
rl74LB7Ax+n7KVzHj3av2PGcvPie3dhEdqjwKNs2/y8T1QnLoOQtNmryZWMFdani
/hkhMGTlLsYZQS+54KBqeEulhVO2cSvuOgtPJExkAaDi6PgVON+fR27NYlL1Kmau
BeVERbzLoqpVZUbYGL5B2+PViZcWZ1WrD91ydGOolklqJuJ48ZHwOKqaq0xFRA6i
SKCrmtkqXFBMvkJDK+8AEdIeYgrEBeyup+3KKA6A0KzseOyOQArYehRYEK1WRWii
T0R2b8zbFgWBgs3OOQe0pGAqx1Vig6uXULJP1CGlotLXTX+K28x2uvdvyrhuMrp7
8FooyCyLtX1ikkfWhlqVaRonBBu/fsdSj/DmRkpnaC5/PLMMf2Kxt80EphzaYUNN
yav9sXO5D+u4nvExSmEsFis7DAp1xAUrCD56TrfvfnYKFTAiUzIliGB5vzTDnIB+
ndxRf+zYz1o+/hrtth1U1QCvcnk6Jh6WRkqFEgpqWP3HRYVVz++1LwwlAWd453M0
0XwnBJr6g9D0/zLrfLPZGtEj1+Zz9o9JyAl79IKezYOWF0SjZpybJL6LQ+rnz5gs
ezB5iVHOlN4HfFywDpSBXe3ohWvyy+1sc8XZjGUclLb+JGughHhBgtuqYkVTTKNz
4wzOHvvPK7wfXw+xVjgrvB4TTI2BxXc5WAT7U6WM8u3XraHV0KyjyUCOv42c/5aX
eI87lbcnLrp9Q0ePn8rmi7Fp5vIOxkPATwrOGBNHcxJxVrGbyvGPCK9GWrolIoio
yvy33pZgbGj67w/VSl0xQGRroTjK3xJ5HqqcL7YXMK1aEsxjcBUqGL1++bf1/Vp2
h9cFufNVAuw29RJM80Ig7S1pX2LXS2we5tNWRPr5eA2qhdgIdTizV4oqeAbGObpS
e/wKtGsL/vLVtbgiYK3zxJ59SQoi5ikIrZ53sSpkMbtPDAT1ufi9q5IpJLXu2pyp
m8WG0aHCFZj7GpjNawyESmXXfkk6vOwPMJ9EQX0qhAo0F2QdG6tZa/cZBSOYJLpk
TjrHD3BsxXbkncO6JcplVqqzQKB9sqWvgamYrWkSAx5EgTvP32VFVlCnjyUwme85
ldp+5XcwKk8HvlFLR6cy6T5gaFgG269EzHXmtIVCqWbw587ZyrXx06IA1Cvb0S/R
t8Z/bRWR6C6h57bZnBhUNgO7aTeaswwhwg8GWBS2IEA11LU4Yc8om3SRuH4/pWP9
L4yf1zGz5FMad8QIGCcRMUxDIED29U9GWL/OKxW6JKx5uxNsHCAhLcOYDz6bsaxJ
4rL8JaZlJwEnG55+9RYq7xNaRp7GfFYiAkpvS3gCs4XX8VdaHQEufmgubGpBjOxe
/nBSAx3ZmEfT4hTVjpB9tcFJBtYRcAqkHLD0GSN4otu8enstK+nBPmIygSmYW/k0
kkxPAyht4ULdTaR7c0usYXKK2phGortE2HQhoAFF3O3jmFeG5PjTLxs2JtvN6GWl
4/dXWtuWy/3YNQL4MguG+N1vaGJxcpjFCMoK2nwVIGaydeF+3+qoKjQWUCXiU8G7
TtksY56BJ2WWb8IjwIN3ssDJsedzV1nEFIGOQK5AyWDCZWyS1pWJCEWEFX/Y3a44
8UxP5OQSTZnoyD5WCwGvQwD++q8+9LEsQiKH4XJg45pEMULsNLKQqm7LHrYJmzBz
MzrHuOONs0Le/jyISQkqdZhkcINJ5WVmm5ZNGZrjXS9XQgQFkrJWGhIwhBLLsLwg
pg9f8lc7r6XMaRfoRZ1GsMeVFDBb548MXpQncEOgNr3xv55Bz92tYW4QjKmTXx8v
FNmqJcH/5zIvLqCO4zNSN+p3Bu2lwOTnI1jG3pOkexx/w5KPaue258VFVT6ucxmv
w8V3XqMK1NFCBEHdMBCgAfOLlXA+Nxg2gQSthQdbLwdGTueAcSXP1lTvLi56Qw5w
kcVj2nFk4Wdj/dNnhwAHE7DPekFPJXEyW/J2tqqCWjq2C2VMMXLooqr/9aVaiQU+
1JMYudMX6zlIYWF1Ifg9kP6icImnSARrSVj7NNZ4HslcnBmiClptiXV2kyGoy/iJ
SU5Kx7u0CPffUPE4A6TXcIDHU9+oJY9m6V9Ynphh7a31Ctk1b9utK7MbAKLQchV6
m5nJyGO54FfkjGx04qU/ii3tPeiiU7GVNIf4USHlDiGTUZTChLUyGmNN6V9djO3f
ilsuJZoW8p0oLwFUX4Yx4xggo4va3f2+o3+Oc8EuEhcXuw0pwmZD2vTOpP9UjNO9
wcRF6vWwJKlFtjkZpZf1myWoYOo1TFhESsMfjkV/dB1vzxLA6NqKUGTHX0G5zubK
nw9TkKTg6Bu/vsSSM6Nv3RvFrBWEYy9K4nnkVIfnI1W8HoQdRPpQMUYL1DLxLyAK
C+8g1oeAlQpUR4uoZsI7LHEYNfG+4N2Pio/DM8ofZuq0gsfItkqP15vCveMrFyve
ICk03++UC4jKac8Nmo8z/nZyFpeGfkTNA8wtoXxB8cm+P6xK31736fCbsCOenCv2
uus+dmAezrPBgqw98Y5GSZZPs0OzvfsUG1J3u+ZmvDE0jTAgh1eXDEd+PAjpgTNw
N/6ZiGWW8NPcSf+KszlAiXi9dkPIy6n8dVl+rK1jSsItxgzOBeqTjJz1oZFvARZt
DzNDYVJAfIPhhKs2a3z+2W4UuWdkSEApj0Ef0M7Q78sNOGeYdP7phRRQFT6AENqr
C6bDDlD7nB54bIn1D/JDvDNlLuO6vYJ/6K2tDeBBp5AH9BQosixJVn5JkYtTBsgw
EnLg69Dow5EZfp3NTgTGhAGbgyg+PfNRgGHARGuZaOO7RUf3o/HMxdxs5caeLEFF
XVUnoBOEoKXMIbTuX7+ABdA1b+0xvD2EUDqClMBh9QKN14pM+Y847nKRmGCppnND
Nwpx0b714iZzpRNNIKe9abTNuXSoVYYuhgMNr7AMYZUruFr5wbsCinjl2v/fyT3/
IO2OgC1Mo11+qGkPRhNgLrXckrykekHJmlKpdM4+68jQycrr8fSTVRDrxwXy8Rvv
iL6Kq8PYS+6xnaWcYJJmfdH9YBBHZFlhmPbC8khiyd0on9tb/BMOBX9DP9+1ECNx
8Ry7qulG7SktsdSj4n/Rr+4fm0/zBsjasuRh8yvxx10+yqx7jYC3FKEDWnqR8tuJ
bi5KGRSr9oi8NDP4hXm1kp8WGpLVdaNOn1O2BhnpsJLIIR9r3h5iTQ0eMKX71rov
nrxOhintk2e8X6qNwTSq9X2tdlsk+cmWdH/QHiw011lPDpnZ8eay3RTUPn3eoQq9
NMgQTv6A0HurX5o9L9Op9B26Kjc7g97OwsyESq2lDp5euWt/H1T33gdLifEIN+yE
dkrMVp7unJho+rUcqIfd/DCBC/4x0ILVbJNgd90s94ZD8myuqg20e5CLZ0oUZv6+
vqhcmOhI6wetp3MXHKKMnlRxSU0d4I0ynErTKfte6dEgD7vpdJfdNe4jshCwSckC
N3K4lXUJ871cYm4nXO67NhVT+yeYbiH1eEOgJqMKquS9SCkvlDf9oA0aGY21GkLs
+FHUZupeTw52/BYpT4x1qPppgaT36yTqiHCXMBQ98hPFQmra4NDWDjD9wVYupdcq
LpToB2yYsxX5S/b/+LTCt7Ox+ZjfBHjNaLhaiTrxflxYspi87L6TcVFkiaBBZtYB
EltPsAlTNubEomeoT40y4WjOzK1t5zAbBqZo4fUfl6bmP12vGzqtk3SX/ZYcehzq
Uw/hO4/K30tzl/W+OzHy0VYPKdtn9Xh4z/f4MiPaIIHTEhrsYADpHOZIGm/sVGjp
6TeNICjqeafNjYPhxIWpMp+k9tU9I5Q7SmUEP18IaKOaknp4E6kSKfNJxaCpmvou
kqJNxr/SUlV7mtgGFhQJMuSPMNIuo325ITFl4Pec4wPYH6qYTm0U6LAmkgF7y6H9
AUVXOJPhysNTxO5+K1GJ7jDpbTzRYIOK2QOy6D+gyC7AUK1WkcNsG8yTBn4d0dOf
8xT/F+3g2pOM6Wkv5xMK/azTfHqCJOw9Y3WZzmQT3kF4up0HtOH/lnL2dN+hWDlc
wAwenEw+U3lD7tawK0c/rOSGMw7ZykT9gA9+mQiwcHuFuWhjle13ap74I83Bcbh0
ah9pe/1KGS4QI/W51RiODL2bEb6dD0CUl7dY+ltwmGVDiVo8MdI8kkzOONE+d3YE
X/mz3O7d3hXX5yiS1WH6j/Z8TbgzdF7iW4MqwpDXJOonXieJmHwEYs4I/jPnkTBE
qXzg6Z4WX+Yv8IJPaR2Z97+68cb+OmHcv35NoMtQnb/gwY+fPKorGa+gcrWWQDVx
gDTWBJvUWepnfmrmnODjz017B/dKOr3ujX8XZw7KlznuxEyA+Rtl+/Zflh6DMdwR
KPDVbbD5NOiSF7QBISCTi8gm1f1p6d8Qvf6BZyyC1Fg6tW7i17EFGEKx5zjr+RPc
5wXfj72wHxwDEwATM2//jv3oU9G5+WWccEJq2oNREnNfupocG66NMp3RrpJpu3V8
sopIDDV9nqkomHYKu69hruWCwqpfU//Xg6SRsLM56tZ7Q8+p2JZuRDj/r/s0/vmH
Aayu3yiYaKeWCQt+EL1XDtuq3cWQVN+As5qEDZnJ4jOgUDDosM9ZsUrnyVcSo0KC
I9UUy8yg5dWDIjUcpjj7DQWa14l+zULgJlTHAX/Hq9gtGfXcZRLFMpgiBHKUWsLI
eBhShzknCDhzNihnDe+lzMLFBZgg+rGH9AhtVCjyFoKQD7ZgJZ3YlMtDuZnNSZGr
QxFWRGqA/n6O/TAS5CKzWLiiH440XIrtXjsM4t8z31aZ2rwkmMPSJFdVyYov8LtO
utIEOTdVjhWfhE98+iNPZ11q5dd4bzs2jiqnDGMcdDUFwebkJqrz8ut2Edce/idR
rro/i8giX4SqBvjexn2344/XGq8fih/p8t7M5/e4sGnHRkfofK2f+yxHt+RPOMCa
7JSlFNpj8QAwcB/hf5etzPe0XUWlrtMUoCN5fhCvKHlSqCiFnIaJQXCo2pP2t7Fd
CxKHN1uRo1/zp7y+mUtIJmkV4xa2YFMPDFKAHSCP7QLvdSGQd6ira8A/XCh1kp2C
733YCxqFhYvBn4hv9Xg1qLtVaGfoDfrNq3oR15Drh3V+jWPX8HGuOEFWdCNtImsf
Pm2Ddh8W6VbS3Yd+zC4LETyCc1YaKrq4g9xJq/x3bEBAXWIiXxwF12ifcbWl6kTA
FqbveMNWScGuSU1Fc7SmA3prh6XqhksnBJ8tunewZ97HvAhr13dr2lUSAW+MXUmH
4D+ElZ8DXdbBnDO+T3RntV0VfqPwzLyOq9WUJjxCxBH0laA6sxS8ApJK8v9pCmUm
gjcM9unGW46FiBS246rYRKa9U3tPJXecxXDz0tk2UEnEIvIY7FnNWMqhKptaxyNA
ZlRMcdl4BqgIf+zIwBmJHa5cYphuXUzonAi8zP4V4gi3PVdo1Mj///2RVfNNmhb4
hF2VBWDHmGpQrfMW0Dg9NcuahtDTfr3YnQEVkxmmNcATe/HvbJjP7u9SGFi4Olsm
n5oJu7+c5fw08934bb3YIKeqh0P5pEs9GYvCJEaoUZgSb0tG5Kj+b0eL1scAJ3Pe
7JFaplUJWTpnxWMOA/YDrv4STFJoN+Mh5bq+0YGJN4k40ek560QTqVV0sMSx0vt3
2usXSML+BwjkmnH4qw+GuiyA/HCaFKd+uFfYTtvF1eaQVIWIcqbpa93r0WUj9mEC
Xdl7b9Gzrnrd6zm5TVCS+CYhrEPgKEvZAlAAtL5SQT8G5eM3d7uogCEYufhS+neA
WjEp5y2p2KfimwfzRsmzBxsNqqwspVH7G+BFzlSOywxwHgpp2v+RSsFsmspXfAKv
bKCr5xQEKKdwsNxZD5PYestRvx3NMv0GTvfgLQZkubKw4wtpxceC9mHMS0HdhEOi
WLAMa8NyhQcEKurn/5fSzzK50jWPhsBURgZ/vUDQDPJ9gcidXW6rwqjHTAnnYEC9
UKGrCH8bltEJa1iJu0S+JUuFvArmXCeBErGpncX2LX63LGRLk7GiibjbSI+nfV4G
h2B8M87ZfDdpP44ICHGzMleXSQmEgc+RR6noVVnb3H/Kl5B3tUHPBzX4VcPCoDl3
xRRQOKZW9D4r3LIkPKdsfEGQzvL0VX1NQTQ+ZkiCpO2Rrb6+NRhmRlUBGEt0It+e
jN9XGCrS2OWxH1jOr3nXSigM+/Xuhr65C07Nk4JGE0+Jj0OnVb7UM9+/D9WdNja2
2I5KXAsqZq4J7qfIurBJSozMdpLXJIGM1yFSl2+x+a10ZniZTxtjm3XAhSSCX03N
kbKLsyRcQEpF50BU+GBnvOnsgsBLu1ygnvA1grGOPJ6a2AUYdPkRirHsUuHVusOd
lmNeNAObLK7tl9VJUPZrK/8zk0vaedn5uiUckfZuIeCW8rhoPkwO9QP/yY8qketa
l9FdI8ZDGGpoWSmGvxSCfrRRXV66umLjsSznkYoB5G0w0IBMvOdqMjbFvIVG2Xmp
r+GIDD3xu+rXfA3QHdIPRbAoKV+9GpS9iBNFwRDk0IOvnvaS99p/APOuqWasZ1rX
k33CwilZs4NrJSh2/pRGJdVgEhnp5t8T8+HhHuFTuXLnz7h4FnTYKNOp3PgfiZbh
GCxMEhbeQU0P4qmzx39rWzL2SDC4yBsM3Jie3Qe3r2peD9nHCWCR1B4jlIfdirEh
L/R4429rTBEsNuK2BzmXHHoUarocPf2T/wAi0s57YCeaqxHiRVMh/LNrY5NyM0RN
+rRxnCTT2TRbCTsiqcE9kX8D88QT/PbhDPWqgyfivR+Cm5yZf4o+rpadN0Or/WHt
38i7EV2UZyZEK1j7dQ0pdEG2+hci4CwOykC0hD7RXPuTtjFALUrROxt/IHv94S0C
4H5ECIA8urAZqp0J6kPs7oko3f0OMroYAXmMMmG2akVmPpwFK5fJHkTD+3TqfuUA
ZLZt6McNaiVLwX57FU03sb0OkceYSHOnUijaHacE7/0H+MCWNGmv57vD4/CGYkBu
lilCBrnYtqWM9knMHpI830LZPNLQ/hLffBf/Brc2cDcBFMKdD/nPs571HJvDOkvg
aGERE8xldOMv6lHoMIjVrdLZ/C3wgOnJerRS1kwlLCgVtOFfaWqkSdHcjRhhKBmC
r8edSGsBt+L2OfcW4UdScUDeGVJwT9vNNrGtfKvBH2fctdgETvTv8F5hZtaE9VTB
ZcLcmbvU+s4IRDTJbsC8kPZvnPTvhfapsBWi6ovpbBC2B8OSEj178sR4F928Uokh
CTPTgFbu7Dgkmt5bDuhV7w9f/aIM13+rx5CpuwkszKt8XZhFaKqB1zKxUMaRd0Na
x+ccXHZWnIOCGJVuCMhXwT5T4SAe46f/kVPCeYScpjY2kYbRd69boo8pn3yjojtM
EV5cAEmP6kwSJknl0ntLKqUCS0aSztlX1x3Mv8KcQAWpqOrA16vM9Lra2wJZhUIT
+Du0mbTxD6sCMn08d5cd6xNr9jLdXFFRDlrZMnYMW5RYQA4YQaUsrqNVSvrFHzGP
6rHhu7SGc4EuVFPiRReuFwsi4JIkLZ0/ZMZ8r8l//1c3PP2fp0VhwSahGPuIxL1T
BKCgKoVkDENpHUKPe4HXVdjvWyH8/F1r7KAPYmSxwhDbRjwvlSph0engDPP6LbdK
1guqZrm886kOlRB2XY9PaJpqlAL2cqN8oXADz1ZHYX5neghThXox2fNLQJ3oxPR9
H4KvaU4Zxq3sw4/d8pACdQY5JyftLoYQZsSQ5fGfnIIzhf+B41COlVJNVI8MSF14
JnXvZR9oC6KAy/EkACh8dK9Zv1uAN5FANzKIVryqNHP8LZuTlHdHnxSZqonlwSqy
F4wPbArLtjAHKRL4r31xbtQ6Tm8HxHe1b6y/RoA2aak34LWUOSoyIrDZBWsQ8EYM
ZvH8qgFrCf3ytKJfELHgzYvU8y0yDkYvLIo/Hvqs3c5TTmqrX49doRLxl14XKUdk
Jjurb6YfTVI6yIvV3R1C8BH2uK7/yphuV5iwMld09deVnQrn50rV2nB7tFNX3ZvV
2sH9tMBElhW8I03YSuQ3mrNcuSgp3Vbjm4NXjpB9UQ4j/YKYKZmQYc5CFhDnjlJD
TFV4/wA2EzpM7Hh9HmmmwzSTNtGgVK9JkeIqUWGXOy31+3h4L/9fcWc4CM0yYSSs
8W0LGAEqg3CCEB3j9BXDFhfVojXVrl7GRxLEZl6MKs8x/HMoPRhsNSk/fhj0OiwW
l9GSSpBOVK+VNgCl1aZ4e6NpTwQd9/VgA0JJG9hGq8quiIHvxFxWcv/3usp7s21I
LHxBe1p81quCckhQnaXeOVJ1WImGup63JnDAwdGH31I8GAUeLQ1xLHIBhMsLfRJV
Z09IH/WrR8zfM9Cd8Uy5ZMi+2Y/kIEAiSX6CwiIlGxu0B4Kxt9sOH89q8mA5xKx3
Fcgqj/zCRd0rDpkW7OV36RjSjGJwdv7FhEFx32Xy9fjcC/kBuy7Aw5lx+uPcAmTH
gVpi6z52hbQG1PVg3/24xAjnb0p71zGY2bfQLxNitF8HXdlpFsFrgeoKTwIohZU2
81spSDT0nXq2GY019dhP5oW9yI3ymtWR+GHiUMr8/CoBQDzZ74cwram9KDklgrqY
ScCFbLtf+BSDEMpgZ7oLW1wsTszgVNceqVvP1gWpWGIpLRn9cTCQQutzbWckAkkY
gCvcNhcV3ea/ijVZU3wIboUv+krNQV/v5ZB+sz0p9D+vuJgZqVFiafyuy6Aw0cpG
1XuAq5ECCoZ9Koxa1dD2ukPUZJjEJAlLCAl+BJpu8Pg4yRmwWeNaPfDirpN72b+T
b5xdIglunO0Y+Ld+j3DXKqr1Fs3696IFN0bAjpwCMY0XxqQaxjWJhUJHjiFqWFz5
6tuY0UmI2DLuQFBpJ05u5ojboGv2YGl2c3t7ULn6ppIGWJOVuzdh2nmzI3GpqyZ6
Z1qAwIKcLSAUQo0FsNR34LJHqixdS7z+1vac7ZBHytxnW1ok9JtAycb7FVD7F/+c
eYwn7kvX53bvQwi9YN2v8V8pLMckfZwJ0o0d8NHr0bf3eiS/jqwtAaX50SKLL4pj
Wxq/2nS2ieKhPIB8hbd3H7BhEoumB6ghDs7phsSARdFgU3ycrLO2O8hFrIUaVgf2
d+Em6xdx7edCkgT+HMOmp1K8NdTSq+cEWOf6x33bkkEa0NLGgqWnqKBKH7nVwsVW
ROuJAwP0brhMvKmnNRunFvl7jsV6YjSU5SjmB0ZQJg+hPNR4DBFNW6QxvDAq8rPD
mLUsN7hLojj+8ETKKAh/S/81QZZM7xPAIWsgFtweSH4L36NvZKgstemBy1ONkuuI
zNorxMjsUnmPkSAxlipYA4j9a4IOat3LLTUrEceb+xtbe84UweHZp7D/nt1iwUAs
3KUAMNK7cC1kfHjirn4YvkC+OFxscqJIs0Dt/gkdpGdiu5EoNDOg6mUtltE9vyAZ
Pq/RKa98rd6USleIlipzH1yRCdmJ99cvkq6E7CWttb2EIc2qRgtTfETlSCqBbrs6
gZ5Sx5iK0fpetIJdgsBNO7yGsn8sEuG5s6y/z8vtAdTGbAzT9Ot3xTGvurr2spbA
o0P3xv66beM3v+eroHb54pEk11PbM3d5IHMT9ehkLtdQ73fPZbiHYIL7wzavT1DC
a8yE5OAyCx9MrHYG0+yVjGHvWbShIvn8pjbENTsUcErWRGqWk2j1oTEtGOOVlVZy
NVdPtfwl5YBwPWrbNT8zKCweqOkfgBJOMtNjjIJf4AkCK1raBfjMZoy8bq2DyYwu
Q3yeJpBfoSvlQajb4QcZ8C8PfQPSzXjwd0Nz+2/hrpIooaItalbYpXfmF3MseNyk
E5BU3A8LuNbXcDxxrkU+FiRbMBwvBs97XrcEPywQfNfRL3a4WAoaxnmipl+Gkg2w
lUer9bgxb8adWq0tTLtzP3bvEAH3uw88vpiOR8+FjEHV5ka59SZRapyqV4i2CUVn
1GGYElrMtS9qfuWpM5ESjKUBIu+w7J7ibU20oILiqOTYKmtozmfxYfxpXz4VeeNl
0aGQQDyr93XSbgsVxTGqF7669pJwie4SiVXU9A41CaBrq4+ZTEydpWi3YjnIwfpm
+O9CN0iDcfhOzM75Qh/LSpXGrKSXaGF5x6e48vc8EUzqzW0d/h6ibSl2Z3iLXPNZ
xqxMXY9Zo59Z79+5hUS2q4ukUGMuzLMEF8wQv0dYRotm5WgaTQE8hdVjlxriEbT3
69XkIaYybsfKVINkOH/sXnK8Bb1zr6jiIrI8XKmMNGPhForZa70qwz3SaDISJFr4
bt5ykmiiaxCfBns/IIeJfbXOgx8EErWFjgYJna52OpEFn8gVnDr3yvcZ5HM0FtPb
NB8ce9olREU6lhaTjXm+oxKX0A15KWEzXJO47R43hO4vYG3EfJgfXLZ+RconahYJ
pbH5IoaxjV7so9JXhpHNfZ9b04EGIFWtdpNF971hYnS03gt1MCw+rtvzqVAIQ6kV
MlTwT2hiaWJmpIJKE5XGs/THkGULNdtB1pVEmqLBapDU+WU4+DcCkKGiXJKsWxm/
XWvVlO6wSTq6+L1cf5nt9oRbKRzRR/3+pVsfl12TKbieVLLFK5R8oHCcb9DmyJRv
GHGWXziWr2PrURo9M+zduUP9XW9iiwSwTOjEYOZvv5lw2phCPWKm+elPWiR5FtAn
0J3r8nraRmKu4tHEaBFvWLBW9gMDIhahvC0pQVD0q/hXDVxFrUHRXvUSzBuQ3KJb
e0wDAFNkWlbcYqu0ZYk+79q3YwNzAC3cw4zBbusdmL+0F5Q/buCjCeABFp0nnrMj
IZT4bFx+gYwcNEBu2PBPy0wFcasZ2xiaLqv7RPYcNMKtob8+U8/YmQgmNHH0bKU3
KEonJI1z24c1Xp62KCzZfVKTUs/XG7l50G1HeM4Qj+wtbgjgZGLcxumhNq21L4F0
LjwFyYZjZfw6CnUB7hX9NKfy5oSoPkXQ3cWmTWFA6mYVA+skleYFAJDRKqKKbSru
Bf5W4OZxpfc3h1cAe1sc10UMvFCboXKORXOsEK0kiw0iu87Fv36ij5Vg4qinQk2a
I/FMV4Fr1gWUxHM4T/uVwaXEyzEXsw3C6i7rb37TwSMffqBDzQcHAoqnIukzickW
MCKWOUOT0GKNbZq5MCpJFpj/F0qAodlo0Pr7s4XshzxjqfA9EFW8C+c849S15hgR
V0K34sG8DxEidIAbm7QEGUlx0rIvDTpPjARH0zAkajsiSINAUmdoY4tqu2dce0kb
xeKmZh3ScAwwNUagxUEdY+KM54NjIz5TBdyRClfBeSKnzJAZ97jSuCCDue5LFNSe
bzmkI6DmrqZT0J0m7m6IzK1qq/KWB5HQ2HT00I1i+qBiE26zHgggTlz56bticxe3
tJuVQxY/hjMPw2tAaRC8glBIFImqkgiAO5mZRKuACp/JPZ8l3h6Kv/H/ohNv4Ccq
CBlGyTWP2koO9h190UBnARALg5c4OfJwoopwnjDyYx3YtlOtSVLSB8/dyB8TuYG6
EpJgTLAijjSo0ZwVlgF110EbQ/5eIvxyDe5qg80mHKmcgZEdoB9euEDXqCtiA3SN
n95KoFvBCOtn3IdjZ2lDexdC/aSMrej+jATMSx/BH7l9PGtgDICtf/8xaTUTKBJG
kJW5jUVFF38x2QlndkthtfSeys8O/GRGmAFHc6vv00Tco7Ru0NRy28OB/C5gUvlw
NH6d7g6l4TiGAOURr13qwcbTe0G7ZwG5cyUQ6k2NsZ2yr3ogkE3g43JFT1+O1xCI
vQ+J1cfGYUIMJPafa1q4Bcw4M5Nj44ry36d9kJUube1y2JGqxQzeHcvB7xofmOuw
bRVBtemWz771rvu9XRY2kGvSwl32QUGhXS24dbso33tGpSaqwrr6BQX0PmVkGvd8
dvgpbPr42odMw+ync1gX5kEm2S5BHv23KbA0Z9x6ejDmsJuMQU8GubIFwjE0BMAN
Sq/HUDUDsQCNQ+foOaf6TK/saE2ojBfAUgME8Q7gcL/PIXwH4fk8QZWy2U8tM8b3
iJdRTDzGzifRRByUakJ4M2DdTmV75XIQjjydTOdRx6sutptf98EG8FCxbvijiz94
poHUgTXgqrv6+ggVzThWJ+aNjRf0CjiYGN+JdTLJeCy6Y+q5FoOkFiTiUlbKdO0E
91asZCkmdO649DmZCGpYYVcsmIrUvhfjOYxKxJwRqYAvgId9uWFPRgHZU2xtUsv7
uPs1iTwJGParZ9EfPzErujtHaWcve8pn82PSBKUufDgFGzpN9nrs6VcxIOPjGTRM
Mha1JbbecTT+sFmX5OVD1sGPbDff7gUBGEMCE80hfia0a9n6s5Xjl6qPAqOxyc/r
MG3StsTyGZ/x9u+U/R+V2J7UhN3ywUCmwqrrv3H8BNf8PVIBtvQi+ZnY8wlt5cEg
WXz9yxiZCzTKty4Lr7bTOaVp2FqAgyaTey/ZswKhgdgXC4fXnpDF3PvfCgA3L2BS
VD6I0J/DDlUpR3ZDbqy9BWD8mKuKtsGl8osEr9FeaGoEznGVXG58jsrC0a6ju2uH
tMPlS3Yqtc6VM2cEL+OKR9ZMQEgDM40ibFlHXRj276i4MOC4fyd5lVoIBozHsZZS
u6EcRX78kDyYVz6HIWE743lMgtiqSafsl37+KDkHvuCn/RZjK4AQu4ws4mdmQbMy
74WaAG4rX9xLaG4CvGF+56bFUxsp96afYbB55suUc/kTkrxfPJgi8xbhcfFbSlbt
xmpHKGMOWLL03hStH/lYwmMAvKB90LiYtWIvgqYsle5BlKshpbz+KWP8TQ4NpYOM
GMimYbIFd8vhLqMYd/jif2Xv6FH666RwpFj+6C3Otj7st31MGi36UUjkfg1Yjxw3
ay7uusOWEEUMO1x3oXW8lJZSzjALFjP1rCP7JOi94LqzFc7t1AyARcUzIYXQ0n1W
Hp72SA2K0Icy4Dq9EmOKQ2UBt4Bgg+HBn6KIUpAxMQKv48JFksL5wHWdFfIAJVXp
7fUSFtIMx4Q6zqdz9roZoyvyNWgQlmxLRHd7n9YlAn7q+ijNDiDJU9UwtO1BgpYe
y2T/kA5cSKy9DLvrAgWQVXjvNejrIbD38GR9B5jOmQQ+nQ5WA4+jgZjYWockPH8I
Joc/T0M14nl2STT7Vww4PLQZW8e0oinhOMHYGjrk9fdXJAdeZFGqb6W5I4iWB9Ph
UYHXaRrwi6iPurrwmliDlWJPxicltLhP6q0fazPOHVNoPdCDUymvmsrYWPBWJz9n
XGZr5ANd5Y2Ux8qJOjZc2OYBmyIBsw4+sYo6KZeiVWgSjLtQpo51glxpHYr94HWp
RJkZbne7sD/84UQmf647HYP7m4zyvLRGEDuE+LeqiIz+hO7A1f4GDX8bEMg1q71j
NPaSEEReUABG3OF6UayxKF6DlCh3MQYyklGBq+KB1WbTd6iPFWtPn8Zl2TEzi96A
SI3Tt1sSZywpBQitr3br4Ke+JJ29CQMLlA3uuavpYLiOvNsByfP47TNXjdCouY+/
yo6XdGCBqgN/pvlgZiUu9YbQQe/t0UYAHLx3W263vDgFXqKKpmZ5JOp/pBwJFxyg
7xQc2K6eG30OYFuleaW0blG/oW+gdV6lc0K2xgvY2qAYNQ75Sds5Mo5N5u3nre5p
pj1eL6dIQIpBWgCDQBzK071zXez+beQ5Y7nXnzfcjc9ZGXG4QvWh8CftD6uFdg1Y
2DssFAlcdE8WOyN4hJeYGjNog8ecjDaTB6/5u4Q6R7DXR3IE1EiC3TOdTa4ad1F7
I9BS3ezq4gguIVfEfGiCaFaeKbz+hxzSbCymxQX75iWfO8Ch2lPTDsKCJYYrbWRx
NIv1kSPLkdMjLHQxa9GMuuVJUj/h7lECN3XASAAGkbecehTIPaLqCe0988GZDAk3
6zpqv239KCx8JgzdshMvfQsqBUQqPbQVgVNiVJ4eQ7UE54Ufhw6hftTUuazLEcxE
6/o+9uCnfsaCItPg7QIPqGurgDwZkMUY24Cro6YZrN3LeOHxOlKj2Ew16U1Bid+D
B1Tjp4azKaw+8YSgi++Xo+23aYA+sJDzltdv3VVfxltr7ZKyHWQJ+jrDuj1x/Yn5
oSufUfF+QvNNQjEyKDFcvgDmbDSTdMUhRLCkDaaSBc1yUDvE2kxJS/FQ41E1p47U
c2TThyvvGFFv7EvfJRqYvNE7ZND/b8JVO+G2ioG+DjuMivrzxsr9L3vmW/ydZBZN
ptCu3Paeqmf0apeA2zfseSdr1/ffIXe1WIQX0UlqSr67NsRK4+e4b+tZklNVWKcQ
AGZEodbVsOuHH+NU8389GZxceF0wsR9ZxKhEGVNFz8W0IADFjQ3ineiRg8rE3kfX
21HVO6/6eTaXdsgotVv8CjfkcicJxTdT1I0JwxwWs8IP2k0xxHhmTOcrtq7BfWvk
5b4DGrzsOhjcZO26bhSKYHmilBFCu2fFFDopbqviajx8q637/yRL2Vq1mA+7DfXV
A3VjLHKULfWYFJeEcNHOz9t1pZOOvV98yejwyVESXWT8zTIid6cnzrHU3wLJidEN
sL6rRkkfwynsbk+KmbjyN1cMt5Hjg0KchDh13KvBhN9BGAMBtUSAq6lZlETJQ9HL
CyJBrAMSnm8umxJnxxiBEHrJ8soRln6eWBDbiIMMqCEONc97m14EDwugiSGA0LTT
8ubcL4MP1NYkS6DVqNvdnfbTFlyNKRg/lwuRz7UcVtsETuX+3CBc/O3FUWp7c13A
GltIXW0cmuAa5Xi19KPct4gLAfHLdur0TsVAKhFvC6Ut8nTD0ET+UBWPkWPkL9Fz
mbUCIq3ujQQpd2yv/H8i6C7UdMe2yNyXw0VKQjari9X0h2WH5DzkYXdM25toV4aP
Ppb8i23UtrIywjdVr8CglyK2RdLy+GoEc+NY+vHI7yTIinKxXBPwHja7QKAv5WBL
AbW139da95sTwA+ENfZv2LjNJhuylLmUmBRtc8HGxEoBiEEg4bpCQ8TPjJmYgbQT
sauI+hyKGrh1ar6RsBjTtYXlJ3VEz9f/R8BuQI74haqsYSAko6qoahluXx68MFY0
COaOOoIsJgbOgqx5Sb8swHLlG1JBAowHSb2aQmSCf6kQsQWEhAr5FXtExScG4OOJ
fl6AY+PMIg+02o991wd4+M+c7sbjppLGjO5erpnRlqjy1/duBucMHFl3cm2wzL6U
BiUVw35ia81es2K5ILH14vSJOcOVWaRJr9Au2n1p7HuG78wBQ6xOx21X8NRbiWBI
dOSHcGpCF6n3iBczi0imWBBKzLy+7U+XBvb+7oQ4EUJyQLo5jGB0MSn4K11X8UzG
l/ISgSWlOMYhkhUMeg7UTZQ1JY3JTPyLFia5tqoxxRA9K25Lc9n1Ll3WLuESHp1G
6MYdh4k9C25dgcsnuro4V9NQYJDP9/VaV0GRxL0wn14fFNhf5JURdogzkNY06IMH
VP4q+SoEB4phWJtzubeY+POdaQnul2HTnExn1CxIjzR1Lcp1bYmkeh1mFep2gKuw
dVh3vR6UYICblc59X4yWwzaydoJSkonsecOqRZfHr2A7qMnkxkJuLD21jSSB/aEL
MDaWOnBrMWdtCVgh5hLnKRxsQnrE7q84X37stKC3VW90Di4f3nF8xqRJcvmFc1/O
v8SqZa6LonOokaxIZV0DcikNGSOm7NtPnxBOvgchEZJ/U3qKtCaZ1Z8EfWfaSbwA
OFwArJtQI/16baVA6ELN8G2SQYGe0tiRcjAaiK8EhgSF729FcPhEnF0Ng0RVisSE
0LmryC6gswv+K0HtQmuqz1AlHpo51H/O08LtY3w/s59kYpOT/ZR0ehj+xAKG/ugj
OVZNyqZwvacmf6xhHl9rbgrA+IxUowtdSp1toVvaysqAKX5NmV0gEzqXdw9dIvKx
2DnI6OvDuGROqaNHGehKDEVNxZHqVoiSQZT+SiNSC52sAPAQfOPMU4mZUF02s4wl
p/lRTfCe8eTK1jAHVj+M2jM6+n/nI7+oA2FZfr1qSam98tD4XSKBtKYolFAzFa2c
8gcWQwrJN/fDbHeQydEX2i1jyvsOKbmt33XsV1XIPgvTdDtq/hhdoKULZxCGqsCX
vyY1ZXTXPiPY8hw+I0vbpVTDk3LODd8CPsxlLtBTiS4JJ0cOnrxZzg1NGvewh5eG
DYTyZtgpRVunsJgKxDBYm20u+702HFzpqT75jZVrZlZXYD0VYHnIwj37lDy/1cbS
UjDkUubeLqtd3dSvb+BL2tBJYomixnMIKY06xYSb9SXboFywbU9sIpLJjJch9Imi
wcn38j/MsI/Uw42Z+Hnq0XX/03CUy8Piu4ZTSQMYscN6xi2UvUe5nKQzDhM5A5Ok
iVwe8kgu+YfMmw0UJpwgSw08Bm5PB35qkTN/cVdxeNgVVMXit8nPdGltfcCoYF4E
bekMVPlTpmrhGxuKvsK1r5plcm03E5Skdpxmj/5L9KcgRiAlrqycCxb8ftdYunZH
8PzCuahQvEsNcaEauC+dFxg08tXl5d7eEpUdVX+UJmyOwYKhd8qw9lEHRLSVKrLH
K8rjA7fN5SxbfYlLDb3co7bmcrXimlpqUhBEW1NwnXqrB+Lv/6GM1jGKqxkmDife
JL5xpmRPS21htBMlzBBULBc1OIi0RQG7nY0stvl4D3W9nPBp5VSAw+RTFkEbWBzX
jquGOcHXdKDtM9Rn21YC+HovzB1hJS1hE37XQB9r4ydgZ2pSc9R+NRhZ78PAT3K0
AoK3uc22FQUJ3HMqEKm28CbdnWFgEH88Xad0xBCxYzGNlkbsiNoU/FgPLunQUrcM
sKO1xGG56ED2Pepm9ZcDfH+sfX1WwntQWxqAsfVAX5F3fpKRvf8iAiW3C8F7GlD4
msb2sjTStF6frtJCZ0KUn99EmeTmXbqzOvtwUVLWV8GvWLigPcNWY3fpcklJ8UyC
wwAZr+TQgUCjQFewZHAqtW+Fn2Tb/o53rjLx3w1+nb+uqO/zuzxcI+xSVG8RBBQd
mgIQXgBPGwUEmTWakYtN/c9gXtv+FcF+BmgJ19BRNtG/r8lxOt079wgdYsPuE8a0
gVpmiXqLh9529hP7dtvRG5SlUBNUGY3VlD5RB1mj8K+M6Snmy2m8B/bPR9bMczuz
zHiGOc3okb8c9g9T4hi64ugtgegzII689LgopuGthVyZxFEd4RcX778h2HWUZXhb
yCmckh7+N7GYST0nWXGee4T8/Gw6qU4K67paGnQ3cen3wsAcpto3N3rXHOm7Wc7E
96t1E6l7uoeVcYtpYLAgapXdePAUgftpcPm/CtkD8qjPykdFzOC37Y4Oz7XWX0sn
pRtqKrGryHPhRmdTj5yFW0iTZkawKR8+iAnWeMPsoizr8/vH1Da6KgkeBHe28K9q
ezsfC2i4ZTXQgKhbfIILPorZFerkKq+gTVpQXpTaKWBnfKsR9P6esUqSajMQCo35
HaAKr76ksulHemzMtLadj2gv8PVOU+ndITLl40yRQ8ipWYdQvs1C4sQ6Bjbi/Ddw
bnmWwh3g5/ZvEr31dk/mCP9XarXI8NqXzlm6/b2KeG9x1qNv3XPey+4S/6NUOmKH
yYZk2uk2mOtYyFhRYmYr1BHOjV+4tjZuvxDa0fXKm5v0BIA4JLrz6ihTYtoe+Rtn
WGcTiRGd9sSKul0gXetLArkccWi/kfXKwSTJRGXYNkNYrg0hTE4kTMpVexi7ItW3
D60epONX0OGyyQ/yGA/nnWakxsHv9VJ1IL+4FvdNvpolaQjRnNiWF6nuT3Ji/JZm
+LL0ZbL4Q+Xfmm5QuUQZUxGeU05HXBuUK2Mlg/NoHaAPAS1HIi1DjLktv7hfU1VM
AIYL20X8cPq36QKXK32tPOYuJ5mU97G/PfBxS4khoksJhtvSCggMw6ZCU9pogJsC
dh1g4F/4ifzX5GQNV5XDQFvpKpLFaDzHxc8XiYrP+uLGgbBAFuctFfOUZECanF87
XXtU79hMlxR+QL2s1mZ2UImJ4FxV5DTEIKA69wEkS8xTVVbscoY0vwTdKMOcH3oj
YeZPRSFNmV8tcIV8LnS0dbbJTpy75pm5mtUznxjU+cRhG08NmD5yzHPTYqEzJHcN
xKHfslarS7a2Y2lYiWEvvCwuvdRC23JmtndRzidLOTRritVYvZB22SVcCCLPZb3V
qiWwEUSPJuUTcm0jTl4t+W2I8LC0w5/i3RPIlfCiCIGO5g619kMkdPbs9PD4NELD
jdlFUpjpYTkAzSoNLF8DzX75nV7TAa5Bhj0G3eNnjZa3Nt0NbaoHyW9gNX7qk6b6
1447AqvYmKVTSpk+XnOh8FgWbh5yAU93+i6E0dR7AyiFry8pXNbyVkOwOCkuD8Sh
/nlbbF5xOA+xsewgAelmMziHcfeeI/zEROosTbKI5f1ezqmx2uiaoqx0/6cGn3MO
fGL6dd7d03xeLYt6A0ubxm0jeoWH1HVyK7FtChxecHumQjxTP770myyblYZksTQz
vgdAeVm8BKwHGkVhwpgeo4eCL1aGaci4W1gCGJhx5v40IGfIOPo6eR7twiPIvSxl
ZHkEGLAhmyjhgnnzYqlBr3Tt5rAZfyiSdsNdYWS9O2w8d8y/AzhaKWvoE3+r6xuA
nakK5LE+8+IQSd/dvXFJsQRngZPDPkGb9A9dThc98Ji79HicCVxPcQmXJ4rRAtmZ
qCZigNtAXBYQOpxi62ZCRh32a8CcNVpD6x8tvNstNkZ8ugTLl/M/UE0M5DMEpxqm
9fH9SWJRawItfDCpBg/kKprE9ltxeQ994GyYpUjyrzgU8RxbLKkbb2KBiiOv+dDB
w3Z8mgyO+Zp2awmHNGhguc+X9F8awjYxZq72YGk+NvMGDLxBZ82GKQygJksXz9Vf
kXgzEh7yEYHP9z4ZEpo/H6PnBx7yT1zkTlpiKyBfzSd1X3mmplvGRjcuBFtX4DKc
cvxYdWa69PSXxDlLWoQGz8I2rk/UkRwVYnHdmeSNea4EBKLd7yhq6aa4PamRRR3X
uwzpak9joQfX0SHFACimHDvf1aiAEvfXBSbFMO29m4UZWPp2xFP+BCzZ8ZaxM3xS
b6nRK8JtDevYnOQjJ1LwbSEUInk+X02Dh+Gv6nXoSdEAuFCvEyh361U5Jfblq1GX
YLSAXnQXA6IMFcijHnVTPmnBFQJ8IPVCiCojAHj+oFp/7EJP7Qps/Y21IqZtyr8z
WCzy7SFj1oeS/Q7UIvCgd8IcTova8/dge/O31uQSJioVM20f6T35/DYlBIFUoIUg
LVFRcKYZaK4ZSi+/5ElzFp1Nzxer9ecDxL1TYtGBt/6uksF+It9D/yonDAzEeIC7
aRxC/SzqLGTVe02iag5rVRJVa5aDejUt2S5izXRN3eClJ1hl/cqRuw3jRS709maD
rx9nnPFYSx0LJz4AV0gWtyix1QtdrzV9APx7DZ9FDOTaQhF6LpiU0rruWqtfmipw
mMmwBlND5xCJ78yHM+Zt2xnV/36M9L1TEHD4GJMJOnqFbBQDq1CXymLVU+KCdHvF
Z4Cec4zfiC5k41zbbth1rze/Phvj2G6Nk0tFkxmNqe4I/8CBP1bs7vOpzEjyPGk0
iSxa2k5Fv0IhZQYbN/vheL0ei/GKjYOEwbOLHajJbDazyhhOFdTHowbZZ2GOBX2M
aFdOeLSr35us7BedxRlXosn69U3+s8XecSULvX4IzyDj4oYFgDUXlyUkWak47SWE
TIIBtUyMdf0ZnWeWagvUtFQ++jqhdiUUkVm62rLTI6NYSVKtOXAkQ8Rs1IOuDAEb
A1XslXAoMlmup6BPnyc2VXVLBPqgOB6BNSnjkq8Bn8fdro6Kqo/fQYCCYRXO+jBS
pnIwAN7eCCJK/FSw0BC8ck6PHsQIWtToewm6whE0DUmzSb4ib51aIe2cHDIVgm9a
dkBeS5SePDhCYDG67gesz5Kfi89tAMvqFkp4D/suCa8IDMEZlWflCCqYsobxornB
DYCJW8jnabXGaEbTb4X4QK0ZbkQv4csPk8kAsiIdhLPP8GlAinXFaV9r0mrd4vhN
LBVyjbidfzpYSIdLJk650thux0gRToZ2UXGc2BQ/bCoEU5X6/Txm57DT9/lKmUu1
wg6UGPZK5IqHXQkIXkd8c+xQkf18C7SfM/AffdxhXdZiit4FC662rs3s07Ixhhjs
eqbYdPOW0nCwx5SusNirM1gzNS94HdvGCz7juzvsrEiSgvDstU7NSYDvuAG98KHw
oywy0mQES1cwCrjOTBpNTyAUE1DmClQXt0zIj65x/glB0giXczkW0B1wBsUpSMNc
BAt6u8IqEU2JlTXOC0IwseQRfkdDk1jnWeWzcZ8KAlwYxBH28J/lvB8Ssl3FabzK
Y2y5E+vp6tugiUutGZoruxl95BuVyrJ/s8Th7adEw4cff0c0iS5dOCoGpET0qS1J
ra/sv0RAEMM4Uq6Q4FdQLCj/zPlia/fRimvIvpdosx9xE5+DVZSbfBUVDwiQiSdn
sBjYY1sLyPhiqUUoL05sv6VMUUt5jbXf8I0+4AFhT+YlT3VKtxE6CupRsiIl6r3K
P6K/cZ5/uTFMMJJuwpU3+0mJAtQNO30kNfXZscA9gZDt/7LaL0U8bcUA3xudBw6S
gFJddRGqAzxxXWIFcUhaiPc7bwUNwKFcHI8XhF3ylYaYLKmTF4PwVwP0IMadvwls
MCUB1UAWm0kEGWvNwYXrH1XvZXvlG59Mnex5gKCaCcz8t0HH96JianrPp2Rquhnw
EhCNs9WgQkJUWK3VjOVMPJjxmaZr1vcDKIpR/FgdpdfR9WnpbHhZ3ssInUat6+9D
LwCDwUCKDr/TBgERSxSt60IZx7gwZ4kHr4p5Q0EaQSgneeZvaCQQ1Pl925H2kYAQ
TIvFm9Mw7u+HUqVo6g+d2jlPkAOWyXx0O9VBbruCts0ESLSytoNwAdwUAdAEc7wU
T1sKKBtKj3Ere8F6Xy3QMAjEIKR6rLDkIeWUdIn+LOkXh1EqPrVcxeZJhEvZhg2L
hKyTW4ayenpXxzcZzXl4m8Dy4aHPTUAWb1RIY4t4MKFVu0TIm5BAaChJ+kIntgU9
YMo4xU3AXS1SwCh7e++xG2eN81XzSMstqdwQaKLr0fAXPVCFM4QB+2svuNc3Mi97
jHmIpi4bpWKd/rGsqREOnO22em0Dsy8CP61hNZrZCtmytZYK2GMfMxU333NSlcER
joIDP9W0urlZ1ys1vMSEsIvF0gx/r/WOHhXQaEwEWZOhJ7hnUFc89vF7xeOL70B2
WGs3wMTI6PZh1Iz10xVJ4p2sbpuUM5IfHYFuF1IXlOeLAYxwYJneVT2P+n/ecwIk
DFHLQhWy2bIPvWCDkz83giNqu98sM29+KaCm6yi27fFOVuZHcboOqHtaEd2fRiu0
tVmkmnK2nwjNy+mWMzxzcFvFoddpVVn6wx9NLKciOKHZfxUgc2LJ7tkBgdksCNxs
5gGUXJbvgVZxtpeiWMObuzCTrXwzFyIp8JYgMS/qR03p41owes74EDJxfsD0YVA0
A6UmJuwP7lItWrSArniPSlNTO76/Jd3ytfpqH5XiF9DmPY2Dy8/I3KMpES9q7z4y
Grrvz05DzqY1ZLGkG0O6jNW0+m8TyqfuHqb4QLxAlVz/TJo7vRpfDw8hVDYlxnbw
3Kf522aZX6GvMOXwxGQZkcj5ST2CLuih94BSXpqxhkla7IiXfypqnFEFBEZNuAGF
Yw7EVygkrx5Ef684qMErvD4H5aR4LqxuPLPoGHgDNZb5h5HU34KYgmjZiSoqqbSv
wUWX03O1+WVnwce4nj7Po/Fq8yxkJL+v1BI9pmjlNPUKoOCAV2zeZFKMZwk+KGaM
LGTCAk3uhQD7cXPW0N0lEIWz3uvl3BvMBSNoygkSHlXPCKv0NGs3TmYLK9AoeHMX
DF0B3W6VSxOwDJOTmjZZZhtcKgwNdT3hVbabYBTf28rdplj0jZ82rwJ77k2Qvx1x
HyCyIA6Cp/SzuxgeCaX+jHNNRqC3saTUeXZoxpAhImheSC8fy4WZLBKhtnXEOihk
nLXqwZWHtvIbPsR7UYyOM7mZm/J9yWNvVFbBA5xIlKP/i+SeHpQQw0e/d1axejo/
o9fazhpqIGoJaNsDAO4W/5eLYOKs5N430WqGgR0wNJIzzaU0OIubtKKXUIcV3EYv
i/cxr2ixxjbZ42yMsUStrEvWedzGBd+dVYauPMr7TQXAUjgNUAAc/pOnTGqSf5vN
BfdczZuv19dLQ8P88PqK/XYvFQ3vsKJHwuXKj9BP0UN4e7+O4pqxgwWZlr/GLOPb
Rai99QFJrj3ZaVZs3o4y7Jupk8Gf+lo7R+IMPSvYNLlO4R1BLBJYaz7+n+vD3tXN
DXD52qPSjUoR/BAdta9d3ooOdqFcVdQKOPfWnsFR0Iglv+727Wf/LQI41kNbIKFO
n0V6BIj+sIXRWENqFPr3RDIo0EHd4/o+LOvQ1nHMakd1+0gy9LZL8POwng3Yq4Jp
r8BD1v/zcfSInwd0K1XfY0xw4E//7jEhDiqm+aHm98C1hkO0lDTbbeENZHF979Ew
UNVGeK7z4odCCUZdzdDwvbBsugz4HoiaI/gnSmjLCK/XTuEL05eZk9eMbw5dWkWT
jfApDW2Y0GuspDpx1kpKODPyxT0IMpyQyDPRnXVZAYDIuoL1RY1KpEEycJLK1MWc
fLhPN2yLcQKZQTLyRC07RPBizoOe8dX/21LuIbueAQ61fnXMWgTdd0exiOTbBeTJ
vzuUQ00ICrh8LTyfPKv7CNo1taC9chxo/eiIjkfOUEdhuT8+RTunSaPsRp+NEKHT
3mgf5iUtOeXp+sNbO9cW0tsCSyPrzwJ0hqlqNkEXCbQX5PAQVAVIzA5+qXfvST0q
igD60n728usCesDxW5ZKkvySlQqx90zd73jyFinaOBNpFCKQxld7qs3NLSQkx55J
JZCbpTSyWHV216C1TSr8ayz/vR+Ozo0WTrMO6g6aq9PXJQKv3ImuNLE+oYjCHwfP
O0YmMHWxW6jBr4GWhp6uYps73WZ5juFdy6lhKl67yrGdUpF7DaG54R+9lL5xLeLh
Q5Y6zYgzY1X4NO/2RrXuA15CFppfjF48wuDNEsbdxHQ4GyOP+B+sepLhIj6d4+k0
KrMsTC9yl+JqLR6cTUbvHqZCnLXskteBgVsPu31MItvccZa+vrKD/5ToEm34T2VZ
vFKrqt9zL9GYq3SfR2jClQXlwWqglgH7gPunA0tmImLsdQtvowEFWYXJYBTdshy6
OBiEkYZx59ZVhyIBnhECT6YvMqoBT7Hikp0EkAATUCVh1ejfp8s5UaMYD1UL8f6V
g0XQkS8XVSIbEdvOjCgXiHe9LFdePwa+NlGGB7tSNk06nJIjIGdk3bAACwoKe+B2
a+WIM7bRwlJ3V1VilQMXGc6h6nOqL5K0Lk/eC5BaA1KH/poWzIUQP6MfcZPZiZBz
efDc/P6mXN1JD/MziNo0LKeMOMMRvLacWEiu2UhvTzYjeN+NwsNzQiY7Aq1iRLgB
LgTiByaLxEor6BFUTccT3ke8mE3jsUHjrnc5grlVVedxBDMCM+/d50Wk9lgfP7lN
D1XqENnp574HyCnL3kaP/MMEV1IGCJb7mSJ7sBon1uaYGdheyWhvTe8JcFcqwm8Z
jtAoexeicXsSfRfr9+JDefkU7bdkvYxn18ApuRgOEj6K3rcMrG6LGxAhhBcIf3pu
Gh0ouSxf1JELt+5CWNQ5bkflm9jJU3IBufaYkt9NW/WpMfOpuIHv4mFepSHe9koE
4emfttoZpxKt+nBkHRcvi0ScAR9xow0BCTitfRECtiYNK4xvzbsyt0VD/TxMo/HR
pdz8hvWTV48kDE/WH+490q5Rf1xVNr8GYf0jF5hZG6zKWZirWxW+QmjWz4+gV6V+
/Z8ABihol32cgdBvqCV04bFaEILFIZtNFrjKgwPflvWMquNy4OH4S36scj/Cnbw1
NYqO2v+hXflCUrJ28fkKpt5MyjQ8W4RLD3YSWNbM8yrzrtz+NZbQSZ1sePxPvj/r
yenIJWqJfCZE/GKiki45xkRJ39dA6toNyZUlpav6sIWj7tQieZZDajEY1c8ykWbL
V/ehkdOH1etRLBGtFXPiwf81tYUA8r78kIA3uKlSGatHY1H0xDmtzGgroPDxUBPq
fscpK32wrT4+xGoE/ArmHhnKrT6n66sPv6msBBInJePFF9zpVeT3sSma2OkBwqR8
QaBxk5SNMbnOKP0hu9VoFxvd2HpIRrZ4GJhSceB6tvn3AlIyPbElbozw0orpxBd2
xVto9YJA/v+mKPch5MPqT0ZD1Ib80p7SOTNhxbfmS+ga15tnWk4a6mNOeHGkj1XT
fatuMr0riNiiSPbwKO506QllHIa8xufiY2Ys5tc6C0VHfgB+zHPzNSOt+JcX0PoZ
8tScxpvlYZ0Ia1tHG7WGfJ0owmrANb6oT2rRS2optXpPPqc/9g7fe4CoKpbpu+gU
dAc115Ebx0L+Juf+0PftCagYpA8To2dMUQLPPBrk5R8GPaH55euO0F6Y1xLMQM2v
irDYqjSrD7VPY2ByR25Ar6Ne3OinurRYZMwsYeBdcGnVvadZKsKVk+XBSCIf/8zB
382pFn0boF1CAmWdYJNTH6F6YhA9Ruee9qtBvJ7ffvyp57uqlf/N6yUtF6hmRdCU
/VbXLRHbsRBc1UQIjeGo394YLHRFOcd8RvgIsLbg8mL4Yy55JOGzyDDlixhELEI9
8yAs5pPp+DWKtvuc+Nn4+3R0A2/28avsokiNw6067C4SxLls8XBSwPopkiNk5Civ
McKaVFSeH5OGTgbvCS1dYy6pv3hs13XBM40h9UmjHVzhacbYdkx1JwaJi5ClBZ0M
/ypUTHC276eVvymHJUti85YTc15ouOItGADC2cGptqEuycW89sx4C0TlGwNMXjqW
sbTKZK/jvejmk2qmiSHXQW4DfrYsaGFBPajjECG0fwoOnYOxQjAJexwM7njj6FDB
EomxgQZ9WW80FK/bgXV51rPyag3WQok5SMO3TgISxLXUVK4kFvUgu2vLRn+TZYvr
Iy5py7XZ3tcgE6vUEFI/L8UHOM0W8YZ45p+YrDSLeAMlXZcUlsxLvNlKjQRyYrYF
XEmIK3bmHsFRFXZWUBLuhls4Eyxrzv6uMzJui+upJXXMvQBDOgSSioGH9GhPpRRw
qizNv9LKh7Vf8lmqtDkHNva8uD91H1rzxK2SzoNFVLHzvECtPlkl8SJddTPw1D1N
+v+v/GGToDAcUv1vywcVRa1IBw9CPtLKCI/eg+i9dx8XxJTeBLJK9hzOFlCzeagk
JF8Klna00D8ay6Uob3l/IdPuW0e1s4TrW2kZxj4oARGUp48TgjaMHpLUwq5Uucm8
n+Av3gPMIBrMDtZYdRQKfRWyTPG/FPaIkpuE9ctV97JPtyzjPPPMsgHn36bP9E1I
vmReK/XJoZyUKnYVNN5zOJj6oVJhvqxOheiifTaE1rw8O17V15rH/eGKOMHXqbsL
evnjSAiVR+K2DgbOP5iHqM9geiLEJ0R6AFjEoTv/6gdMWJ4PK86a2mBYgNOaIEFF
/RTr60Ig9c+2j9Un40Uy+ZLdKrEC+th9Ty9rS0IyqwAmsolRLEDk47gWmTjmN00B
eDzL6N781O30+lOlLVWsjqr0DTrio/yqZa0ys+mEXlmULhUjV6G+e/mFf3Z1twgX
Do27jeE4CAxuRl7pvg4hY7AafZQ5mELbJE+ddAmz8HQGy8wDLujOqJCanRiRbSdZ
MewlkZ4xfI5+Seuk23u6Bezw1tlPR8SqxEx1Uy6CR4miFvk03/tyuOXOGJ9WgcWh
DQOgxjKFnua7jkvkGpNNgVfKX2vvl0U0Gs/W/YUZj6QToEru+NliY5phCGjPnc34
tUGTScd2HfUyf22AurVOcrOkEeYrSvmmfShYcOBtoSnbnTDIG9bQOPw7iU6wsuPy
hYqsYJgjjrYuTcRi1ZZ9dhLrpIy8lGnmNZBL4nkPi8P2AzuEg7YQbY1OTQZ2c6oV
FLwDLMyNHTU3uiZX4xpgznePeoizDmnxB54cVPy4jVTJX5lpBgOZYVyPjH7bdEfQ
6xQYJk/FB40LnhT7TBPuGIbe3gVuXD5h+kbBrCFYAVPjBdsxM8Hu+N7Qbfzf9kDs
54cGVYg/1CcNyBWFKEURpRNnxVUkr+Celn+WG74dOKafmaGt5mGB/l/4FzstrZhm
b3xTINolYq9LF92w0Sqx18+BT3jhD8AaH6WnbPyq5xOdjepBYPx7dJ1fQFtfWJE1
U5Qw1dS8dcxRng6OwmT/vBjW04lt3TYjxvhAZ9QeksXZSTa0SS1Z0iFCHP1aC+M1
EYvJ9pX+Ino2E1WxJR8QZjQX6VAwTFRHizVA7gEo7QrPUOqhYrSBRLoD8glN2TtH
iXoKIVYQlc1DwIJf9uxNodvTsJfjQZOb3TVTQ8cLNDh5FnHsoweyXEHgBz9juyEU
tCAogeTUGeMypF17n7ErOrjyhFxUN9cw6Cv//JBf9GOnOyXQCwXhlvAAx57h2JE3
Ai2IDOocVCvfKuBEK0aRrZAthJXCItgIFsTfl9ulYMJmpgZtiu3l5pJpafjRY6aU
xdzYMQAvWsECn4yfn1HCzkunWyEBmyCv+f/W6dPopLf6fOwex+14zRNm932RvVfa
dCqY/TH+f+m90HezCyAAp9qQeEHFyrp4A5funqGnHrJNivyyvXfLDXV6uhBq/dzZ
Z3052UyciZ+UaUSe/VfSU8aRJ3a4Vi4dmNMd7G46H8XQT9Xe905EST1CeorZcnsD
bz8saUbd5r6B0FdVXZlzD2fnFmJCujdFgd/zhtKaZEzclz9v4x5jB0AANNgYwfte
250nEZSST/VpmgGimjCl40NH4F79OtuqrTw3OZpmxD8YdeSAufmAm/PK94FiU71x
wg6EROFqy9n9V+DFW4StnlmKnT2Sir2pQBuedWZtMGNlCFHwq1ldmZr12wR/E6IY
gQpjtM5pGXW+0ZWVsjzR17v/0SLBHsJeY2QRmH8Piaml8S/tlQ1S8VfMrNSxiHYx
y9nkauw5ii8sqi1E7/RB3vPwmugc2TWAPB6IXcFFuhJP7UjdpV9F/9Mn/OvM3LVI
oAcz5cqZND2pvl0JJ07vQCqo/KxdrTHaek+r6hX7JLHXSyWeRz1tX4YI0QK1m0Tp
8vLDQtdB0+zq8sj91daVPIqOTTG6u1PG/2+Xaxc3KC7S0vVAfI5RdfJ/lGi5oen1
BgII4Lq9j5p7CndQeAdqedYfpDDqHFppeTxpfOCk4C4Z6z/SDabMnxrfV/H57iD2
i4lTFnGlw6YmhhgOl9piN8MSkVYEaKYX0zFfUaJiKBANzTiyD5nvFoEN1X08t+Nf
Ub25cw6+2V9WeCRyrYvemawXRPH5+iCpm4dm7EgZT5JE2bLFB9A6dLYS1T2Vec1f
o05cL3OoNCu1sYF0BfHMo6DZvMwwqdoOcf9jtVY6FCzE8by81NL1BcYpH6Ulu1v0
19SHRp95VujTmbZOvjr6jnLpJNnKdd4XI/OE/ePmoloEMj78VARFKRY13D4a02Xo
F4R41OOliT9FR2PKv863x2WNK9sjW/OmX1ksvT2GuUlK5ZS1d8lVWzLSCgey39yC
IccJwMBUEvPDEijwTYJzKFwHbEWyjlnwsAQNboToYPrvYdnloOP05fTYN4jOEB54
FvPFIUwdvBKz0AyFO/qKbNugTd+qe5UAfJGQCijk8Y/rWx1eNG2TU3CB9OhVNkOr
0z9mzVyZIzxUcryQti1intWd6URHQkn7ZGfen7eDmGEzGfaCTxzLxb66SppFGUmf
CceFSENBOBB/cxUugZ67dCl5aEZN6LLvNN8vRJ0oisR355991eX+zE3f7ID5pYeS
phrR8Q1aQyQdfy/7/+CNlekqmhMAKjFz8X1w+6CXVsMZjJz3HwVU4UPrIqtaGpQm
LES63ZiMFMvaRCUz9MlHhW7Izv5ShW0JLiZVMADAmRU36A2jpSoW+i7uhP8UQHQX
KmYzOOpVPGseT5MIXX1YIDrKQa/MZoNCgst7GK5quSz/yl8ZQw6XJwSvsRfOmRE2
O8/Z/jXIQYx3XSrBY7tCglOdGJ0HXcJoOCUtZIP2URlnyoTEkkAbLRa9YTs+Tr6X
fhfilgV1vC6L4KS+lx1+ywnxOop1DecOBSsuEKoolJRR+xLKtQQpFSe3Al0rtJZb
xikJOHQAnEgG2f5YN9Gi07MEo+eWT3tWfoZCIemRD+5pVp1eitQDZ9Ytnky6X1G2
4DlbDtXyJIiPIOEgTVJSytWzOwqCE/TIh02EpCs8T7swUDro+jPpMp5N4xLWEwsf
BzJKaBt/ZUC5YaHFnN+tiM3iMn474+uDIhzdssyCrPlM2mRy7Q7kVvXZMXTZIFlc
lvd1CZc9bAUGyB6/iiUsU44hvf83VA2yFdqy07BtWbzVaJWy7cydo69X5fWKmHRm
p/r3LoNgRavOJBOx6e53yUU5AG3k3dJbhBkVkOd6VTVqu3q7DxgWYmzuXBjuCn/8
C3nOyp53xVxbFa6Fxptsp2zp2CoA4Z6eihKaryWsGaYXBXd449zWZylil2RL7TPr
Ngt48IfrW1bohXu9pGtci0p9iKbR6p8bG/W4gux3JHUU4gl+dS1eptTfsCiyFMnQ
9ym220os84wP64PakOO5gpBHf0HIDv+r8aQ3i66r967Hz6GI5GOxoWPpSxsYHA1k
hKO5JIEc83bklCfZuuqfca93R4+4ngYOmDF9UfawxLG6K5usVVTgO/0c3RkrHpTc
fZJdlwEMZfPFddlEuW5TfBGZlExXOziAlvQdPRDM3uGxcdslfMLMov5dOs/ldD7+
h7+EaKInOMedM29p3rcFuWwMSU6AtSIa1KLe7+ATREss2YfpBHeNi/p46ykQTIMG
w94uQQvSy3yzAFbj2XGt3KhUWPfURBweeGeHFnKyg/wadieEUX8YJOKM17Ton9l7
V4n5eehq9IiS+0u8q/OPbz5x05apcvaY1sJf3N4Lh1+xyP2pjynPjp1W6tG63Yj7
RasNr7Kt9jCKJMvat7TSM6v3KAwNwx0YJSIfyeqNd1LKtWRsdsAL83vNUZ7WDT/E
kzP1TNkiXIaXXeIlZYodk1AwNDxjTFeKUddhoXl2ncyzzDtuk0IwSTaYndU2wDdh
ieM47m6mMG2W8LLiF5puWXRfs5JBeiIwdxMAyUcuujQTZVLBT3tZpKpRDbJqOk8u
VUpBSOtxPo1bsW3GAVI44Mrc5o3yLh5PLKuqynbSffmv0wu13YnQzSNPoyHws4Ar
w0GFRTVZ4o+XJWbyi8X6xk9FABRbryk67pRrSMxldZq/ZcthgWTxOGBQIDNmwdO5
RpK64C7AsfE8zYDPw1+n/P9pUmw1kISwyppY0Hc7SAJ/I8HtwmhoIfa05GHjG7EG
SBbA0bJnVuth7sjQPzVlWQACMjcoQqJfCMjVG8wHm/ajsuMKdFmOwlJLhPXhh2Pr
iA7GwLQeC7LGaqhKIzc52lbm/eXCwrqXF560vVkaVCyPdygI4pAtlYEdj8BETPyS
Vlcuofd149QD849+Ro1OnkduZArh6O/xWne5Tx2j0ZdQ/vscfVajl+96sjclL3K7
/O+Xn+hZG5d+kiPiw41R/JrFZ5LUNu8BEIz/+Hx56bhkxIZSnkMEMy/V56RCav3v
Cm//nA91Vl9z7GH3o5MwZiU1CkjWV9VDcoYFi40SIk7IumYq88UGc8ZtKzW350TO
D6RyZ7PPZ5uXDt7BvswiQ8pVH9YkNN/lhIm70mq6H9Gi63KXvorNnMoF5mIJ+xfe
xFePcTEGyA1UjRfOs9xlCzZUTctT1jTefikhZqUcqpfYGAbEx0soX7HzmNygudr5
Chf2kQeBxNIu4eZwdebTj3OpdOcU2azH6tCG8DmDSYbBgJ3pGt+D0rEGHEububyq
L35s1/mqQPtFFLQzzpBKFgVrLOAgOdX9YTSII3sX9Jxic3MaH6DhJ84+HMrWY6QG
fvJc0uQMuX71OFALKilza4l70fARqIuVx22Zv53jo2YV/halV6Hk0U5WGyKmEo4v
QTL445h10wmGzIl61Pl9y+UBtyL38KW+zHphxxTgltq1IhZ5Dx2Kw5bcSPB7JDdq
aaaBFVmE4b49JzxRusM8BD13gD7zkR39+BH+PCEIIIuD35RMOhurwRP8eKNZcPA9
q1fS5R3Qvme+01JRWlPHvGHnvUo7b67WFLiuaSjxF6HnjwzK/NPKBhogsdsmzboe
bUDQPDTGIvqFlLOjpfsqyrFN3w9FkAlgI6XqKfVMEklQY5JiHeqZxt8JqrDbJOOb
CWi+zfqGSzT4vzLwj90RoBt1ijxO2PrjmcKpcrd6iM0KEQTLpNZMsmvdkg/f+gc8
Rzv1plKmjQUOoxl1FVGBm9scjhDtyZGalQrKGpp6A3/YOw2OTs6hhiqaNRcnvJkg
1TqcJjQfuvvqcR3J7qC+ii6CnDBjJEjpgEGq5yW64ut1himn+MChLKu4BGuSmBvN
n14+gi+AoRARBhcCB4hDIZhhm39Nz2Zx59+1HtDbEcWp52P3ZvZJz4jPIkcKUj9N
EP9R64djM2VLrbhYAhQsi3KG8zGOj8cBg16t+w5lp4GG/7+tQNDsLbnzttoYxFlz
BqhmmtXtj6i6XCCvLF2As+AKozxVLsDYKaispTfuyUrMDraIINQ7Q4E7NUmpbQzH
X04jiHS1rdOwN0wWHftEjQT5LoWtyhSfAVkXBzalCPEexVtvJBMbwOESjhNeNMmU
QqcHM1obN/sX2iXTo508M/JOfU2eje41Vyv6mFAX4AWZJpTXg+qOGTuGfv8Kc+Y9
eXdRHqfSOv+juVjR2gdAnYqrw+kUZPnpl04fJxi/BDgFbM47K1pBPbtAuA2eRI7y
jJhtS4ON1pQZD4Lv3DMFTaxLQ81mpImGqLtybCAh6w8HqyeKVeS2tlI5j0jhzK58
/0RiqIoUNU71p3CgYOMQ0fQjyOBCZTodtFPicuHPkHrVtGb+zD1yAp+Jc8XcXCvo
3NefDoANOa2jyXnO7QIfwiazrVhMKmOSgsA2ua9HhYUIzyGIppCw7PVVD+m/kN5A
OdNGyrKBWE/Dz284x1EPJIhxMVhPXNTquWRbzIJ+Zlv/Nb81SVERjSa31AdzowNY
EZF0CKjKg4PIsLAf5qg/ekRMZ9r7XxU+Xgzs28nLuNLs22aAPV+fd/rqFTCRqqfe
/tJUKVGoocWtduW1NOt31/MbzG9Zl6/6GutA0ntuL4QLCzRv8+UDbe53Kx4VFsMd
MXp6iQ9rkniuT5v8daRRX28oPub5m4IzjEKQT2eEeWPwYd1aN4vclKUaDXnYL/HJ
Rg2DESLuEjN0v5WFoxFYVos0BPFE+TB2EDKBpwd0Sb2o/Hzk8EBVeiasiG2OySFA
FOW9xSFnKe1CJy4Vj6z6iEBG8thT7LpKCAWeE8YtYnUFcA07PiUpJy2aV9FSYF/R
S3We9LM59Sj88O172UrVsQQdzo4by7h9Lq7SeI7ER82VHXVQ8W2uTolRwUlSZAlc
BXTnyucLwXnfs4+39trh8XnxyDGKZ8+pR6OyI36bYSByezErOJLK4Abe0Hp/qhky
XKBlGZUo2jz5TWTYYFTBBsLeo18ENQHtcXwWJEZvJlIoLkLAnzVr/pkwUOdGfjF8
K0/DquWhjRuHgUODL8WPvAiu//WQK+GUGJ3Rpdxx8AR0IV1MKFf3lk76B0YNRND/
RVDWh2YrxOIKp+ZxhgMiaybfPgtgZnAHXWWloIyvIyI509fd6PH3b6QDwJkbxKqp
kLK/fCrLcxnhoDfYJcOQJCZTGBWaJCyekHU2AZvu3sOXRT8V99QUtQ9FrPeQgK4D
mIeAL16HPAwOcXjDUk20WQfI4fXsYBkn5mIuJa6lBVgct5WHu4UONew6eRruDwnI
Nb2Sc20Bm+YkxgVyvCXn9LEc2HwGisgvMh77CedHSz72UG/7iSdr0l6Din7sq5az
CrJEmPz9gQB/0+oyoDGyDUcDqHxeB6/MCVaF94S6PoO4frRqFhN2Nq5mVHJqfj4V
HMPlQ97XIZbBJsTG9+QJNosAMizTAA6JxEhsPUqlWWcUXrT0oGYie1+O4wzf/eUH
n3Boui7cJ5IAJW/LDOlJx5Ab8qKHvSl4xBY/H7UdehEFU3FwoPxnArgTfNrOTUZb
FYYDVxF/16Nj/ALmPFAQYFPfezDAsN0M35x85wtjUzWrMV60wZe8iFjFBkdIs/L/
qEnjjEIQQj9PCkH7j+gbpwQU1nFYi5/d1xRwENApVYnQy9wNXHq62CEyLWvn7/0P
qWkCKy4OTZsTjbxzBQTxD4NkKGj36X8sHTUPZ3GKFzpbmS/eiobQJHr6xaFktiXB
WQsMZt26XakNgqmAgXvO+ke9E0XDD2XSD045JRRQ2kQCP7lhgC3FMxVQjhhMA7Po
rvhbEy3jxy9uvlGIE1QpRPAx44wMNSsPJQP+ocCbx+AWrbvJ5Sv+4iOVHzoK7rga
iMhhVV2El+btA+12Ao0Liv7Xxr5xKdMHm9je0nQlc3llpXuoFb8xHnF5lA5MBfBa
znWGz12frGTRGm68UOIa2RKivmjfB1SUVmGorGaRgLN/wyWV4DDby0IfU4Xr9mrf
WBge3gfzvs2Ip40ZIYUkbwz5648y8KZmJGFz4Ef1wk54ByyxH4ep6wGDoPZvaA/1
+8Ek9yMiuMmcficRb/Da7vg7I40sOXnZNnEYcBOkBd3A2qbi8pfgo6uRiVwJ2BcI
T8j/jbfceTu68chJ5ENR7dY7c7Yxc+mwqiHHBwFSNbsaz5GXGiByVIwWwSAfdbis
aHU04O+E6tc301LP64MPG8Da68L2+2habo4+PqD+bMNa9BoouiMYJUNPQNu9yrEM
T7c36VcAQKZuAE1BSooyNx/5Ebgu5j6x+qH/RagcPDtz5A22sjPNXnNOJrhN6QkS
Dw3qtXUS59ta37t41lrI2C9XW0ykYp2eh6/ORfFSKJ5e/ec52W+HiS4JrwFPYNqO
W/oW5y6k4RCr2ss+XncikPJuhB2/dWrZgO8AV2H4Q+VQUuXfLVBaWzERu9JZ7+Mn
ueg/P/86DBCmUidvMGm/xq0stMk9E0EQHcDyaWXW0riq5NdMpSta+kvyD/koVJry
MNCne8LxFiH/W5HcXnb15sKbxfcJaEBtBrmsoR+QmeFVbXRr70ST8WooBVnA+pEH
9Z3oVgajUi+eZGYftWxjL3TxUr8q/gLSW23Kol9hNOuNM91/2mqWBmkqv2SR69sV
eC0M/xS+VcAXiwrfkoD/CFkEPK8TPuOnV+ehBwjRW+4U2TUUREiSh15ljH08jBFc
ZQjD/r7qV4vwoqb9C+EViYybCRzIAReL0kirENcNHfRfjFsmnNe9MCBP3UEyArQz
6fA4vj9YJG23UWQdJNVf4Ejto50iuUGyScpB/oiGIirpwHpVt4oSgt48QL+S8tf/
rfPpcXJQ48VmmfXDd5Pbt4nTkNKN79SMvYyKKau4Kw+jLXFfVM+gDN2gkGD7og5F
LKPVXQl9eNem35KWHmN3PJ64TgfhCRZGpEaHuDCBANs1rztsseWFJze0zg+asNfM
baYCLjBsBKG07zUjYvE++zXUUZOPP4hVB04i53+qhsydOZI2OCPOqq06LhSsThbK
JCiNBJL/dMCCo4VfhKzTSK8pjZVou8k9h1VHr+RSbsow8UEATfYCbjVadI5nJBAw
dkI8qzONLO7U9QGJcY7kY4bbCDgE//bKmP6Kio4x5s4ZQ75pvxr/4lJn8t1f/FJB
rXJZnejtQT7bD7X7TmdO0sd/v4lXLsCtNR5uYgOrDj7gkuXGF4f6xfwnZ46V0tyT
0S8dkbNk/HBI7Q6hsfqb7d0TKN/VgurfxWr2R1VnKOhQxqtobjopKySdanyyFRiG
wk5qhV4QEyR0BRGWR0pI3UwCDHvmERjI3+at8EWxVfgLN5VqpTFHViMdgcv6fiMn
OUXBKAqosB/fGV2Su12zYSWGqqaqb2ctXe2jVz1KD3rD4ZRK/nfyDk58JJ9XfH/Q
ogpBtqJqisi5su5OPA8vCTvQmShlpV9nWZHSV7WiR44lVaHeX18zR5nalhAQv17V
1RbwYmNWzBkgeWRRsop0/CUFi/zoo4Qk0JJ2P4MEZ6mox9v3IsM4vSqJ1+pjpcLi
HsN7YkgNh8NewadzXuV1i76C8Gq4ormAE8YuMxCWmvhHY5DBP6nyFgEB83t1l/kT
GUs52GzKHevKkcWv5f1B/NK6T+Hl6JJWaALQjjKaSpNXTWqpNDyChqO4Vyos9UZQ
r9cwJN93nWxRt5JphOzKADgVcIzmuW7CTWp7e4WEg54jChZ8uU1xl7mZUWKURoiw
gau7dSWtvuTFZNUF2v5hKe6GExc7m/S85fTdbyJol9HXjPPIwJ2AzuPHxQNAapL4
pQscIhR1a77xV/d155vnK0J1xJVjQgELJh1TjO6MTYnl41l7p3WZwFjpGID3OdvI
dy3wwurzBcMlJrQbXH78qiETEAygrWJqhAmgFo9wX+9aCBhwCjSYNMfGI886grzE
Nndgh6WC76/Huxr7fIouLdOda5aUZQtXZagR7rzIgCIMsn6xJvit6NdVC5Uq6m0R
nsY3xmtc+zUGV1Aw68jGpazWBRKdSSNXvsBORWy00gJrtK9YzGmMKE5KVbsCwaA1
mkaqREiJPD8sUOufnPcGsT5ey7DxOnZwLnZkLmsjgKfIiwsNc9bpONfaVM4dF70k
owfekvEJQaw9vhAoSsFX0fp8Cuqohy/pwBkphyMy1WUtPFpwl+Mva0bYVrzKHwBJ
vgyQD5oENilQ8NJ/qqGmwfOiwEqdfR7is/ARDBh/0WNL9zocWIHUIoT9Re9it8mu
02XH+h9fVJEjyPSjZ5yZ0J+f6OL7nvnAB4ecN3QQjo0rEX42B/1ZXnSxAtdTDbvg
TuMik73/nTPgf1wAeYa2SRq9UOseFlTZgp407fBocBUEIqAxpKptN4LkIhNYJhcF
z8ezoDZ9VrQwUSZeDwmcylDZTQILABAfhgaJgsZo+zy5Vt9NVmI2Jmxy6jfgT/t1
eP2OL3JtsXUi0cehBG1MvyhWWHS2UWWqY6tCY8h4QdOjkTl0+4/wZgToxA3iGBdO
N4HmDj1z3jn/NhX7jGR7/c5mf9Hu8JC4SJ4KV1wnViaPQFvZr5JiYeD6PDSbUatQ
vkBg721/TF4eXwZikLOj5ky7LDb93aoLejZsb1FVdPsfIHzbgvKFyVx0xRU0tYSn
4ZqOLFQzmNZBo5Y6MSGwVGHQx9JrUBKdzCcOKt1OS1PflZkThx0DqSWkxRFQeFea
T+hK6aMARBaDlIPRIyQWyHVwjoi4c6B6b4AhNLz3DNAt52pvtnXfEnkCaZcYLkYV
/bZLfbYP8wPxlEDv/I2yHYzFoqpTxNjzFPro0xMrutxpCi1BJBvHTSjou44CukP3
ETG8/GQcdgI15n2KBLWGbcBH/h2PdCEH30XlTrmZ7j+Lzr9m44B/cVyW/lf1mu+/
GSI+RHMRnsKVfTY3SUvsAFYoQlC6N/ECjWqDhId1QHtvrQzu0aqLyuYOqN5LH/wV
a7o5+B+HoxEwM1TgdLeB7bOPqH2gB9AvfPF67i48TxCqnXrhBX6c01AN0JPRgvqQ
QNL8oUd02qGmOzluwufMC9Th3Rvm2i7LVPHbJwIMC9W39/KxTtZQ/ro+jIKrUFFL
xU5j+E/7rxfUmKw+1Dx6r0GP02GF1vDia52bSfpH9dzb25lJmGM7QGdtnFCj+cza
vbo4LcHgTs0ftqGARf13iAI1ENZW9LMd2+GXTiRweQv3JSnewnNZntyLZICqXNO9
5/7j6xytkBT6oUx0NOu1OLh2QIKiORM4fWCMjozSfbXYjROR5d0vHyTIaNY29oCa
OB1HJSI/VvF/G0v88PL4YyOGbx+A5UF22QjN4b7/JMvhDUn2zo2FRZNdBOVubdbR
tzrXo+eb2O1tesKuRXZ/u9+EBKYb/7eDB70lfeEl629pFAx6x1VXdiN0UzN7XtV1
VVogU5lc76aqmdc9jottscjv6ahucKQdT0+egaftdwl9dymNH+I7n5AfxQEenv1/
2AHz0QgLAu0zuWpTAd62WqbrJOrvCgfqq9COUb9QKoLzCgXuC5AKX3AdpHLEQlJr
L+ZqAPFQjXM5S9BYmFfXzFcI7KU2PrJaKKGFsBzBbpr9ZWxxsk5elutUlmM/GnB8
0rR0wn+rsEjXSPXC9Cf8lW+r/VnNEbBT/863lW2t7WW1izSKjJOjqcnWYjLAlcWm
prdi+gaGa2kFxoiMwK0CftR0hI4OV5VXi/OibdUnN3GdjnJZ1r7hr7EULUF2vJSg
Xs/jsn8yS26PEFQvp1nZhOH2K2RKSDIeEsDO6g4PMtKdAKILtuOxgy3+oh14I2NC
UdZFbrsTf4kY+cpoBSe2RxWnkyoZOW9vY1x0q4C3ojKm89HPOzNyqDL1gVb2JEVy
FBsQ/KTPB69mq9tm/598yJORftfSH4P1Vs8djWCsL5+Jjfh9s8kk7mNRpaDGdbab
8MEx8kt2Ygk7QHXLG+Sb9Pk694vXVTJOFdsFwYam4MFShSOcMaLGlgWvi26dGCCh
+uYshDksHaSicOpDEGyFSaSBhr+0hU3ehb20PfKT69A+yPO5HN8ZR6/p0E1R+tew
5uJMc0gWKSb4tyGyBDpK5dZhvcosZqWJO03LAyck9tEl9KsDxFoev3WCqeZSADOl
rYRRgkFH+qKgI+yQ7ugh7BoZAvoM/LBGQtEj7jFcksbgMsQYXOvfnLgYzdV+d3j7
VQ9gNDn1FOy/XjeUZ4UAR16yPyZ3uTFBeVVhDaXTLwDLfKZQPSK+KKvn8Zxxpyhm
mlWzUzDfcPhLctaLpA4lW9MLHikHoMX1Ae4l1cap0IhJD6zK5W4mFyyO6xb5hJsL
NzpMrCaIxiHFG2ZptQ66a4wCicrQP9MAAK7xz/ljoLksJmfwP/C9Bqf6+AswiE/6
8fP7cnEML3TDrGWpRb9atY16GTYUhbqcVlzdHBUivyKAf3lajDfan8NzOvuDxLhz
9PhaQ1OISPNvJNIGy9zCzgTmiD3kPvozZT4cOJ6WabxQCZjLlkq+WVvbrMy70t77
8/pFUPHQr/gRdAU0LLxsbDrCtKi0uwflv8c7oEdGOFNx7hcWWiPkMNYb5boHC4Pz
L6rSWG0WYapA/GFK0zZqXPTkfW1C0QzjoO9tJ+d0IkmGjIhrlwDuBCN4N3nE3nUZ
7FQssOLCgnp02RYeqF1LTMHJSb4JdE0po8EnmIi8TPH90qSQgN6dC56BvP/pMi+G
iuW2BOG7qjLyaTzXOgnkL3aAq4AEJZc0crxBsFW2UN/6DqPcfavJNBMz4zs9kpiB
L7VagyvKw3j1m3n5fnZfR2A6bDMtQQF0Mk4HsNJdV5+xjpTP0bbYueDfLKtrLtCZ
HX93QVR5HHpMbQzOZC8q6AdX8HQHj7Re9jv1Ip5gozQf+PwwHOC1fiSBIan5qJ6a
krtMtHQfIOhYmOBpR477kp6PvZ2ebIFIV9hw3wwh0OT5nhapJbwHweah4wYiF5mt
Sxb7LDh2o0wA9IOQ3QtpC/9eRG/OnfW0OaR0WVw06HwymJ7B5OWCTO7btXKzfm84
u5z2jnVCFRuCNQK1nR529uMUpWsJryc6G+NL2hrGkzAj9Sam5jhD7X0jBWTK0MCl
h6auO7YmYnSmg4zt2vXjdYaeCVvNzWV/yM9rTnVQTCITXbO5pQgmApteKoE3SyFd
Fkmj3l/8uZHGBk52E0YClV/x/picDk3eG/sEKGo0JDIOsv5bmOAhisPkorNIIqM2
ml4GgHXVqo0Eui+Po7yw4WFXI1JHtBaRi6WkCzHpfJ8MGMlNmK8FqyWgX4k4blpm
c96NNYksc0kUL/uLNhqO5ZFLJEADyZBwQCbLhnv7F0Cat+X2X3mboPEzvVa2J8Oa
q6F4WW8LH9qsVxfaTdMGRsujtPVYznK/GWt2jPyyQHqpSZ5pVDhCYOBA7/KHFdhH
kltmfElDnZNku9v1Den5aBRT/isXkl/C+2linZL+TdTfW/Rv7EWy93EPV4E8hANe
VP9G1KMiUau6/LJu02Ry/shilLjeFgFOJEvzx42kkfb0nbXP0mIoy+J/R3oAmBQD
y5lXH0W1dtOtcGGwwk9C1YExtZ6u2Fffilq+vWUR6tWccGRq6quZl7wHx3DEiCcF
7deRwoMnulMQAMbtstYov26PMIcfhmMOcvKF2VxO8R8FMkJCRaI+m68ZxVM/au8P
lVWaZga3M29NpQfB2tY8pjNByxDVYCYHx7pdjSyhzG57h26DHyscN20fG/Vs5rCX
wAzVXr9gU4gWoJDr1Lj7/reXKzTLuxxwu/M4xS7xudClKz49hFk/G9Mr7Tx3bhp5
OLJSVLha9LM5gPH72uhvRxx3kHPz+t12ou2M9O5kHbo4JpH2owoWjYSQBIMjW7Bg
6ulJirQrItUxqLIC9ngjgRs4wQG9GI+o5H7UvjTQzenhVR8aHbQYyOoa1Cx6cmNb
BtArPwLUqVpqw+/DERqU0a59Ktd7hDhdXYnMjtoaoq+rZ7nhOaZM4p3vZeId7TRR
jFUHuVZ6S0fnE0qbIY+YF6nv+p6yTdAmzI8E1/ENKlZAQb7DOcB6WJ7A1JZ4kjD7
Nd61TBsKxIFU/8ZhFViz25lmPzMtE8g7tmu+TSpPsBKcHtOtl5GaomG8lqnOUQDR
kcCHLtgd5oOabmsVRLMmuxsk1bBb32+CK/nBeWbl++vMBbNjRqtLIHD3FE7+F9FB
TrZkmejHNMetfw/7zHB4pM4QrcHk6pDYLyTDEo4qtq4SJUF6QN4+2l8UeR5iPvAK
onwSVPoOa83xhkhose0Jig+6WMOmBdplf3ZTzTFy/oeknSMAIvBrvPAgHkIiFB1v
yQLBZhAc6q4ddkwfU1NKfJNqRZRQA6nVFMRiSt4u3f131oHLueoxZb25qOhlBhRD
ua7lrnWMDWDNhuZhxt+SZ/+iIpnlkX9V1zy/G6c9DxU3e6c0DJC6zjtH/8ZTtSTm
knguaBRAb9m32mYFme15X5qiRB+CxN17z4Ms8bXl9eSK1uV663g8P3Eb97TVmvth
1iaLozaefSkPLniilt2lqbfJKOV8vQvYbGyXWJ2scOs2vugoNyT7Ti4JJaQCmY4S
u9O9ZXnXSjj2EYBViWL0WbWC9SCQywE292J65uTh6u1ruzWFTZMV4+Ggf9mNAnDg
kjI3eluQOKfh2xc1vxF4HsmLHadDZ1Ja3Z5nGyoONcQhTvC9h2Y9t5fisc5gsOlh
qY6d8i1QVeNhRlpzkHL9XUkN5Gza9l6qjUcrOhoiV26o/2Xl1YYzf2MIvGDcV5kp
xsYaXhjyzeieijVwOrdF7yNyeM5mWHkXqEp82Xlaw8WUnhClbd4yFLbW13z910Hn
7bkQwOLbgrIp6rJs8gt1bTWz6KTEyWi0Zk567AMt+mwX5QTCFkrhS4iXSxmBDSVz
2AulpA1sxzrIKJHmOn0xHIcawo3yFBW8pFvS5GI7CMdbwXG8MW8rVxze0sd6SAYd
GJeCmekNh2grpcSTBuFjZwCC1uB/XV/4TWxV+uHncWzU2TS3sRgciBkrGThb4iIB
ISonZ/pMSmsdXn5uYwU7rA0Nf0ou9hX4aSoNy+QAKrXredvMCi2kQ+FSVvsMdkjV
IqgY26ro0lcq0aO2XCh7K29C6UALm0Ig+UDkvD+BgPvQyv2bJUd+DFNj6nr7FHaA
uGEW06ZxAi8ehRSCmS18UTZFN4TNTpjrJbCMX2aa9HnX2WV1uvVShVzWz1vbe4JG
sq/Gprip7hOLodBjaPb9bRaxvqpUBPxvZ4JURr4UuQgqX77+MGQ1TqwG8muh7Foe
fboiYVTwyJqqztc0N1z4RV/TIe3GDiUc5YVOpkau7yY9WcvPaOvjzlyo5iBD/btw
PvdX70jDlGjfarnP5lEAaP+j2we58MFLB+wEmLpIjg2d83OyzWkkCDj/e6MGEtUm
dpq3WaepIthq5pACy1LGXVZsjp2lyapI6wYSECtrkv0jVkGN792sJstDVjVFWwcq
/VMqbXHOTvEUI+8MhO37H/rum3bdZZl5p1Rz+qBHvFGWogrgmHhl+GkVTLCLYEdz
BzPYTgbpb71IAcHjVYgMF/JWL5Px8Y2hCSpdIZXDz8pBWZ9GeDFpAsyI3L3n74ta
tkmDSbi5RD1+jLQXXPOzE+NTUlGtbgzQ+nYW60WS8bR3DH3gD32elXEmDmUojC4W
gD47NdrsjVONIZIl4secRBQmoETgz6/sKc2Mzfc3FqiDau6LFRC0qS52pNZMsUHw
ntSRYv8rJPdBvKEYPjK0tcdMAfzC7LrG9k6zL8GXGkxIxAjqFNp2HfkPEnb0VElz
Hp0AkBEW6ZkAutY8bJsDgoAiR2PNdJySA6UugBKZYetr4AJ7mtWbOR5fx6UrzDy6
edzFlWYAsVl7Bd3gLQ33tdH21PmPlUdIfEcLKL6LCLOpa6Cb4b0aTl6aauinhniv
FS56sxbVa00tREJeSfNCaMgvxJsOONj7zUOsYUXpCaz4zCol3eYcGBqTKjgzAosO
YfPJLas9iOJePenZ3V1FzXg0LuVBQm4aw/YDqJSAqrmRlzd+Vul1QUAtQlXtv3+h
ItrNob80ezBO1IyrS0mmzAIY0lQOKscYbdl1WAFOUwxjtEEOTZmQnZWTSIIizZJ2
UFkCKHLtVIy+R+iRaTvsYju/KLqguc8EcaIyk90jFlTn3ryf2+9b9PnqoupnkeCN
lQecqAB7pzU4Fcy3u9jEq536NtmFqvNd6sYjh70TQ6KO63Dm6JYyZIO9Px7v0OwG
OOEyh0CstL4o8mjzzzNqjAxTRByojlrrVfTkJhnDe7koFeqeX4s8ABD0ZbR3RESI
Gwbk0cgxGBA8zneRIqF9rwjsAwY1V2kCERZxWuonZhx2rfIfQPZqPm46TZskBkeR
7TsuajMRQVfMQM2P8E7cw6txkqedIfWH23/m2dgYuK2gn+aBEno5DnPr06LWaJMD
7yKzu+vbAwOb19KGPSQJ1KSV8OpACcU/g81R5+AOOQwdZUMZoS3pv3cbkPA+axjM
UGr5bbyQZXYKpYjPj7HnJNeRbWsVu0UswQAZjj4T/RmKw+86NP9eF0fRg23i8Rdo
Luh/jWPEPzzEo1WP4ou0WwuOKVUGcCjmWQCXPZB3vyHoeXiSMo5TYK0sPD7wW/wM
IkNjBbZxhJ24pe7FT0b23baTJK4W4SgL4eDyME86mE3/e8tdqIU4278edteFwL1q
VHaJ+4HMTBgfNTtpmXQUbVuG7lOctDIEQBSPLHRdH/yq3mOQOX+5xjeBe8PiOjWA
w13KuLZjXq7/nXhcld901PbzLWZr2cPduxWrxWRzRzXZEdS/PGJPdjK/ZaS1zf2P
zU3QLZbiYykRdCB+Yzcqj+MeI1md+zGUMbvsDu6WSM0t2Tj6mzre8luefPKqZDop
RAjcIhJY1A/6SDU+JY/ZG1Y4Zkv9ov9EHJ9lBq0QhTfiwZ9FmVEFWjdSL+KJ+Bdh
Bn1Kwxtb597TvJAW+M5iHJAoIfojjfx2kU3z9lteJXqov/+W3a1mReND6pD+KIuJ
EEwL4epcmYyVtklyu5Bkuc6X6ry/foh1IqvggECNftVzv6S/NRj0Ztfvz7AGYjkO
vE3TS1ZhUz6GfgizMg6JYJIuZLkPdiauIIo4rWxIM2lAZjPZj3rvy2ixX6tIyqNs
GvT6SlMLetW7Axfp+XQu7eTw683hy08tLYOED8qu2JnRwRW01/oaosb+QRBIRIV2
kgFZgDbceqvD81F97Dht9Qs06XM7nCQYTnKKXI4eg9DChGWYVn1RBfMljT3QUBuL
BXneHRMsSnOiIjHebhmeyliCMxjU5V95/s9VETbJffRhDB20mOFvSCEvUJO7BIo4
hYFqaBQQL1KpPA6ZZMCtn3kwgqvbncZfDuTUDftnJXcVUMACnUmhfbtbdRBPE8fD
qP/1KNDV0Bz/5pm2zMKwOHy4JGpBeqmFPOtr+hjq3M1H8OX5jpoh1oA79za7w5fu
BJ47DuwCkmeIU1TJmL1manqFE0fuygY4soBqmfMxu/UN9c36oAvqcT26mwwciEkd
/C2tyvAojY85f93nmHVV18k8U4yGAI/CYwl1UzJdj9/76PAPVguXtks0nFdBkwZE
JI3PDMtxu48Q8XSR/56qYXQ/m7Afddrc8uExuvJQ5mCcFHtHtIZZOYb2C+WnJn8p
LSbnawiW5xL82b8jVTyszPsdI1wQei2nha3XqwVKG+a89Ljtk17IFp8LVgivajQn
6RQYJJdPccPaR0tZAkNmLouMs9M8ScibFm9Vr+8/t6xnpHcCqCTOXzWA/dsSpO0b
M6vtQrNf/9pzEJiSI9INtHniEyjiieUwgAcCYcUO5AEaQUSsF/7SLB//Og/4fPm8
R1sgMHpOH47k9X5kraRXB25DwLUBmNSlygF7hwMUUtiUm3eJTPP82RuwDx2v1/GR
061NwCzPq19F7ww00ZtZnn1Zz+cyyXzEJpOSSFwJazNjvTsV1c4M+6QqGNb2yy3q
ht//bYtWhR18jEVvZ1u9h+xI5yMcjCjjIRCepmEZpqcc5d2gAaWCNCwe6U3tBBMz
eyGMDg9EtRRwf/cXW3A5uXmicFccrm+XozKM9ILBLPry/v2VvnbQsX866G3nmP4V
ftfbJCS+L3cxoZ1G+Cjiu2EJi/pq4LQHE5/t4tgLOQ0hTGyw50/W3NeQ7aJ74JtM
K0DqnOgbfWXJHISqfEmiXbEiF2i1o2QDwYAl/UGZH//7mf+33Tzc/vhFtljsuYHL
xa2FcPRWRc484h9LnhgYTnlWKHKycwdo6WWd6+xbhGBy8FuarE1jpOy7U3zqOBsw
6zZTNojibNyX9WGCY2I44ki5sTZyTm2QbdqCbjTzOKQxVYfS39QXrHryx4bDO2cT
8Ey5xcwM20EcuiKhjeldqEUI+OzeGQkxo2RxoZy7WZXNWcdkWW6wgJtRTef1x+8p
Zaoww72OorRluDTpcYJMoE6ayUAJYOna4lJvu+4QLxFKEvTvl7bWW5rzbntWKVXq
ibh+YYCU5P4N+SExzrCdaQuRF0So7uXiz8LhaS/+zFEZ/s8TjMRSoiuO+2JFpGR2
Fka+MBG/uHT1UrelgQq8mhEuVTbQ7u9JCrLvuwXwgpzXnJo8k+Asl9FQxVsFt5aR
9DpMCg792vWLo6v0SsfwPpyR5c7Kfn7psH9QeNgiVZ/LbpQKqyAgKVvYyLOXsBj1
FoVfU0g+bN9K607XCvS0PEYehy2cil0F7UavQhAilYbLZWnz7u3h6JDLCR+5bvFi
21aqHTozeOsx5Yi9/I7nUo4Ef9OyrExCc4mmGeh5VdLMDqx8tHFTkdF7WUogaEHy
g9EDpx01KgMrJOS++QF5VRwkykt0DNXtLpoI4X5SwtWYLDBywq1LK/CeTkNqcfDo
yShRhoG6llx4d2oV3lhrcs86TDEzE5ArVxkzAwQIkfg7Igqlc7aGlnMveluUM3Ns
Fx4QPIBW2kkNflnZkbigt8VesnV7t2gzwa36Rs5fiCTVNkdLqL/JPAXlbPhY7iq9
twJTai3X9bJ1GzJtDQ13oNSdlb5GFA4l02zyG8tkADGKV7lckJu03tLik6avRIba
243hOyhoE0ZjZZhKoq7MsYud1LG/0UAOLRemFTiLHGaVEcE29o8ESK5lo2dEcVJ2
lhJuw+RinavXTG3bkGGYYM+o0j5MUXTQZcthKcYVMi0Qu+y8NDtQfrQgt0G2xmQr
4h/YtuY/wd1FC4mpvUBT0SezOFOG2lbDKDEVPlEF0pCEJnhz68tP4MjohKPyeDAz
VbgeqWadDUCtXIFMsv7ICu7iYaKdsVNkbBK1dd1luP2HyP/hkYKF4GQWySaKjj9r
vJejc9p/xQkI5FEoJ3U9oxor5+SNqrkw2J+lWV78IMoTkfcxgHzJi8I7otfyj5+J
I66A6gGVRRKylizqRqwxs/wYsGzTdpi+Qzf/pLEFcEgv/GrQ/B6HreR4DCOQcSYR
f1gfHQJEhzKo+qTNQCimtWJl3aAnyzDokNaUFN1dTTnD8E+HOxD1EhN0g2wDkGGa
38H79ksjozje16KTu9yn7k8+hh5jTUt54ns2RJcNp2mKrRfIuqZGge45X5OoEyAL
8aiuhsP5xqTRH/4nqAvuu1ACaeopy7j5XyaNEiERhIhsa0AquoMg0QCSPqH0nEkL
2y+orRCtnGJ/A/fmKJZYUDlFZcw2esMhiJHyd2rx0kUI9a7l9l2dw8S+TLawsDDC
XTa/vNnluav5G2YipEIJoA42K46yjN4o779SLXCMPj5/U7k0pozlPwS3W/noPj8/
HMWfUfWdS66QKWLA69/8DNg1M3gRJvfel0q/wTzjew6MAdVazFc4IWeXGfIYZ+ZU
R/PDxyAYLHHMN5mj+AzUExs2L9svFAili/88X9eVS4+3N8viFVI+7oNNf5Gnxqki
h7KZayYa8Ub1gTNG2SajYvVmiYTKRMnTFjAkhU29stYgQVMiJKIYFrN3M95fl9Od
Yk+6Oqhh/fbtxeTCaX7UxdpEOT8QUvnh7wOr0peKiLNMfxgXAxxtkSCJ1PfYEkW/
5SPrYXjWgfPe/b2/yLAb1g6qpzPRgqemc7ZIhu4uG2b1Jr+Y/SrZw840NGtnk/FP
bpH2XwsCexeQa5rvR5LrqvAdbvwFL41TGTflFIeWRoMfgxQ6vcW41IaLf58dMz2C
/clb2/wXAiza/51Xe1Jw2DX1Vv13f9wZX7P0Hn5F/PznoqBlzaEQGMhiHEsZD+ax
83VDKPSwz2BFbOsCvNQW6nVt1BaO2EXNRmWGZ4hlb1WKahOY9DwjOVZ2E21hIk87
oYdYmH8XWCcsoDUn2s6pCPd8Uk1NIPGJ6teCesQF+fMWbJrECsFW2cFPFkYd0iQ2
UI1svoqJ9d4HbuEMvTjmTU5nFHlcxHQmmpUm3g4jBVlpJf3Yu7FVfqnfWLBU4V1t
7qsw1eVqs97ani3QGNSjcD3Kxrt3qrPToR2y3XBBvH5BUgqbHxni/wL5N0ovbIUp
5RLis1AAXNPi9SQUDJad80HQrvjs9UiTFKtKATSNaVm8BIAfyJyCalU8xqv61KD5
mAvXIkQLfPdFQ6i1/s43VSo/J2VuKTFwkGa2QXSw/EatifAer9L1ypcwONhzlTk2
5X6cqNnwzLp3jCWmnACvyDSIffOtaiMDiIuYHhail+gyywRv+sjJKAoVh6lpqjhi
ZDFTs35a/MbptzBsnFx3WcHaSwUQfuASmCa254VEX6GEAlGYHLymdREtF1zCnOuT
akHbo5CRHn++AR4atASIcuMdT+t5OKWBuFNXiRt+rOWgwmuyMiFpVp4VrIBDt44Z
XFHl2M3Uaozs7BcTgkjbdYaV2oMlwzJa2XVWjJwBzRbps0iFhezNJWGPL44xmFEt
BiswQ7jJbfrkr3H+Kh6m/4uCtTPlMiF+f0mWyh7m/YFdfGJjuqofPkxUn9NrZhSO
Pa9CYNUXn2etBLqAyybqcwKXsuS/Gvd0S9AMX8mTXpnx1zIqGE2cVwrbIJ/QPSVs
w38q5r7cDrOQxjbvpkrVHetp0hGR4k4ICSfEGgXaKUdjOgrSizoYzUEFKKXess7Z
FWpZgRS68lw7hRalIxFfNl075RQ7QwonOWp0MWwPxrzfZmWFk48OK5dVmwUnihNR
e981qwT2Slm6SKUJk9jag47z2KLNpCL/4j0jxnq3OYymq5mxhhckHy07JSkp9Okv
PT8B3Cit9Ftm692s/WUG8bZpSGac+cyRi1yMmKv/mj5kBzuBkC9J64pzpiPpKOxW
pHEpevMnPFj5Kii515AfhZI7pEJbKJs3UPIDPc02sY42J8A/gvG9/6rKuoRI/qoZ
rPB5mCokXuAVBWbaJUpVGU/r2HF1xuDjQoBmh/qUknkvL+oOoEBdWdPTwv7VFOhD
q3AYdyiNWKR2/PiNid+7gp2TE6M4msHAylCQ+9NHvIF/nKeLdAEV36YXcbAfl2ND
a82uMxcB2o4Jlo89VIpsIYx+AfB8zzzHfzJ1ulwx44ORG++LvRCfq0jUttvKjZ6M
y25DEBEtZjhDVxd+sM/lZWss0+TprfELKBRBhfRPyZpH5eJdd4bJtpG/sIxaD0/K
wEJIVLcjzlFAdbSm7xtVouZ/K2evSmnuv6Z7Cbe8UBhPpF8jPDoPlZh/RE5Im5EX
T0iP1hAitH7/oe+RZo7+dyRKMK9rhlmCa6ET/ucRIVJWlchPX71eLcdgycaLRnxw
zg0X3cQVMflx+9JYaflSbVhIu3vzs7Zw9qp0VB/EPKd0TeZrhKnIfJUS3OO/hIRL
mDDyLKwuLGFjh1Cov6HOUH3QfW5j1WvHfEtoNzgfG2rhSC31qf+v/mEdUrqinyI3
hvEwGh4IGYflhMk9/K33CXtSAgNeOO0bm1mQCAwlNZyx1fVVxOKmCsdnfCLUKQd+
AR0U+nJkCTaXOz7D8oWPQpbZMFF+zuoj3qpFHXCPRMhqz56MixRg7tGdDE2BV8IU
fFeXDqoX10kCNcnJZNF6fW8zB+1O6fo4NJWNDQoy4BCvMDfuTk4+Cm8NOy/mRLAo
GmHkeU9cbg1S6HoNlqbiU//8P4LUXs9tVs2/04qY41N4WZT1PGXXfG5ysF3F/XlW
DWL2sRo+9kCb1aOVcZzaiLZbSaLdZ2ec9I+83ol7TA+tY8PcAOkAF72ZlfMbInkD
jMAUfuJgBPWsBYtZGq0tPo4GObJfQwMWvrXoL634o6x6Q54yxoTYQL1KPNYUSTC4
uy8+lokPcyMWSPjfabupAy8L/iaSRrSUwslWLrqYpnafDK3q4Ux94LH2cb5OFO8O
eC2nZh//UJS5cUOm9bnEhdkSoL8gh7F0VGWqPY5dCrkz4FjtbgoHVrH2eqIBnRfc
WSRKBNPbbRQIbX/8jbh9QvxuEDnrCb0X+SLJog5XmZ0KNeEOUc4U3HPHBMfF6FPk
5VKaX1EnyXZGODNCKZgYI8RqPG66YcQ+G4eMXighphiaNnyUMh5ZmLoLTHYlj8Fa
4QzfOHHNVdP3Z6N7wD4sZgX5h9xkwk/TsNmdlzOhqRrkGCuP55jOpE0h6Pbl2c49
qBQEXWwXDp4of1nDGOW1ed0jxd446k23EWyhFkIXeHwV/0tAapstQnXgUxalCbiH
7RcZHvDVyAoCJpD3POigkGK5msVmYg8JVQwa+BVyeRYaUEv6Z5fYVkqsf2cTBV/O
uUWOw3wslKojvpifNi0J5oL/n0a4GMVONHqvUfIYG8hPKVEZ9j7sXx9sOQCORAih
B88YmNsGXmTpj+PqdCz+sDkF+ftvyv0yw4NnYdZ8tlp0Hw4bZ5/t9/+E/j3YIoc/
lMCOrBAIAVuv+gQARvqus0snQ8m1c6PiITk5/elDEV2+lGzCButMIAiIWjeFIX88
MnWnJ8FJGIqFE29EVy9rqDGzJTln1g4ZUeANZB2EeoWhnL78Nyr+MEQ8Kmc7JtoP
czUixTmaFEmO9P6vQhVr+UMZkIo5CV/ctPhlP6kQ0IbcWwkIugd4XhRWWaIHQvW4
qJgQED/Eo+sI+MInNvjQcTmxz7bVzerkYloW7N/gb8aBem8hwW1KqZTzuZEy6noo
aHQR7gRgScy6NOEFasCjrdbisW9cK69TkbzaN28fnyjcboqIrFxCjpiQYUSZO0kl
KdZWJr4KbC8sda3kG3HLboHuGknw8Jm3GLw4wMC8lbCZPkjuq/4GtFVckvBXzCcC
+QNzrdl7MPSXkXxq7aaN6fK05LKhAvz78joeS+7j53GfpftqTwagdFtEMgv0xb/0
IsRDWUrCJrGii97fSQZMeSDjctUG3PLnHEjr2vf+OULMmo2IEScu2ic4RBgEB2UW
a/y5ycmXXRoEjceaJo6bNVYNhGjwuFktsEnRvNqkkFd//aZL6a6PpNLcqFT38AMo
1Hn0NIAl0busUk+hzLjOWEVKvhvYfoQ7c5aV2usNJhPxsBOxAJgdeiluuKYvfkpm
gQQ+ZZQf8Su54iMl9+74VCjVkXUquJutGHrNvbHAR5+kADZoBTxpVJ6HJzvQIGGF
mItfo1PMV4VF/LYUFVU+w5CtD8kwoMTqqPlNppW+j/mIy1Uqw3zD8HyxkKFnKqAi
m2TNy36OIkd7ZLxltXyc+nmgmTnDDHojiguOx09AVhBuY/8wpF4jGg8ORTk0zZGh
hIadcTs4f/YtkKtSq+IgauWebdHry9sN+FXpHSGxMA2Yld+n434+AQuBWrqiuQHy
E1OJUiHSb/F4xQ/GksgKr6fonLbuRoc6uQqgNIZvy2NJk0D/WUAuVY7IscKq/gKu
HDgaHPa15YdIArz4KHSxfI7iUgvJkgmF0badQyKQF1q6qE/Xf9QUaqGGVKOUCyQj
0bIKvubNKtlQj8NzjF4fMLvEju4E6oRNixxltxOms5TrY5JNLeuE0XIB7rFmBO3S
VtzoUO0+93Ly+ZMu+gjRDdnxwsVCVbnnQb9zafSkeOV+JiR7Bav+7PZUcShrFsdA
KfNi+QCyfhujFsXExntIWxTTYinF3RL912Bwf0XCpcNfEtkBiQHK4Ibe1dPVbYfE
Cb4VYGXUjkYgJVyZg4tS0c2TmMCOXAoKWz2TMK+1te+s+AmSgLFuw4p1ZXG5V/rM
M8Q1O0zU9Kwz/eWpGyjZzXESyUJgTbDRYkTBrM1K2PUzKn4MWMSuumLjNktV4Zkl
HKP32pI87Un/B6kwXAnFHBW7MVwvRvIP0AfCA6P5Ml8o4LtlR4jr+USlyLewje+A
a+HChBwp0MAMKMO2qIbbz5aQu7iSS7+mH8AWFgEDgmKaQp9LNuYnj5DNT1BosGdc
A2j2nABKq82izTCWzsxrnnCcvgLmbllk4UGh7Q4mKB/8qNIf0Xck160ttBWJ8UbQ
Z7MkjukW4l1H56GIs2R63q4QJWrzc6n9Fpe1JixdWS810wYHY30gk0mNhWdMjaIJ
zz6y4xxPhkWQYMviOaL3oT/GKWlA6/hVRyneKUOhtk4lWORa0OyPwk2p5DDwm+6E
N7OTUHJIbE3z46f62z2V1Ga0aF/6nA4+sS7UaPkCC2MxskdM1OunhD2cYrv2BJrv
WhFvlBIaHdryoZPuaQxxZJ2dPAf81uP04l2YiB4NXscB4SlB1+TdLiqXKwkl8Lze
L4GNZ69hZ4cMXP+RQ0FtcrWOeuFaIfDWrUHq9O7jo8BWJ1MwXfcUIeLTSNgHDIZu
8Fmpub2+UjXsWxgyuT5Hj/wOBmEbug4LhIKnU/39bHnN/1hZJ2g1ephQmLlQrrlR
MaHhzxxq1O47RBn8oKY/L/vxOiQ2hV/PWTCPofRJtn05BA+ZquIrc+xSHxQbb5gw
9nZbD8NvD0dXzLaNRREouJ/0jX+HB/5jfifz4t0a9v69oKxlyP8bCftW3v2bWJyi
FlNeigIzSIvQv0RHMm7I5cH9MOkdKOCBv1Y8IF0okMv5on97BOFu70XUdVV2HLCV
KW1wNLGlUW33HCe2lzFXpEiAg6XoS6PrZawpW0odYUYsf6VQUd5YIp/x19K1wG2/
VS7+/t4mKapjECvu486nKncZtcHSxH4YcLe3GlcVJWZKFQGLDVHErNEeqenKf1eD
y4RO60KNOxz+7uS3ezO9jd4mnavEWHVOmwHiioxTLZTmrLCPwVNoTUNX+/B4FvfY
4cPcwMeeDFvarPCBvRQH0upkYf1+axjVPakWXZURAu9P9VtUaZYHGd9MOT6Zmf/6
Wi+LtI7fTM5y/LFJCg68P7ETIomxEz2kDcE5zmUVat5G/YM2+cr+Ta2epJQA0TWC
3yay56yTfuhYedejGfw0rs8lpGgZWpW777l6y1b1+9Pl0WGZnV8cWZ3gzZWKM5zM
y1VrAVJSp29onjvaIUx86fuKewhpwolZV47scvu0vtQOgAo7/8pCE8Hzb82xAa5S
n6J6WBAQzhWOEQ/UDBlEMAgWJxuFLxaSVeUNKxkn1Bbs5WyRRHjrQT6NxCvO1wfk
DmOfDzT1GaU0Z1EpMzWujtmgYIcEf/khYKy1mD9sCbhgSSUftpUzwlZCn81w/44q
bsJS94For/5fPbeKf9GEDgpN3RYWo0I041LHE88efObwwiLwdeJ3e1X68kqFu3Yz
u5NcWzqHA+gO2zY3EKd0QONxVcskQ6N/l4icCgMU3+q6wMF1VhVwP7GPCcNt0Acv
02Ppe7k5mWiyhLp1pia2NOccKENPILbKgIAVbWv+XxSh85RyRbru5aQkCWdjzIgR
3JbIda+qJps5d+SlXf83PjFZ/csB/7WKO+duQ9vSUi5aED8CiAcWuwwPgsTZC7Lr
+2CP3DnRsvWwnXoWFc6bNTvYS/+sHZ/InUv5ar+hzVmQDGcLbrQqSnlBYZQvfzBS
REkv6UXgymAqgNiyqxHjt+nImv0MHveUFB93MREYdO3yLrhA0ENFftSLMPSoc3Xv
ab5ksXdOLTSO7JrvRAOi7Q6icKU0D0Hf1XmoukUfR40sCyNCpbKNUbeUT8dupb9E
EbCH2uar2QvtU0aS0Rzojeo8da5s3CqvS/XBPAZRlq6KrIyyfXT1Xg1CEK5q1OHG
WcyL8EeHJfsKUZkPhcx+z8Mh0P4Etl6vg//+eQKdzq/7F++uXptJe8dc2noZzlwW
J7spOfo1hq2oHaUkdAgID9TPuBHfgHx9bVsm61qBg+C3KRUTG2N3nj433NnJnOtr
ypIJFnLFxEBUith3Jb6gOMCfyMeCz6TbIRE2NJ44tch9bt3oAQNQiW20vKAHBa0a
ipaz0+/d40UxTaQa9b35U3lK3k7KPKnvnMLPC0uGFGoi9fH0shIOISz2jkZLM+Wi
zQKgmpojPN4tYhaRgXsWgeMmHjvM+xVIkJnw7G3pzJsjB9A/Pat8KxeX87r7cHf/
1X5ARmuXn5kwKpR0S7QUFB5z2PdhVH1pXUkUx8mH2FRaHQT0pchJVj+xLJHSxPG3
t7xBNbtTJZvMI6EoUvLN55CPysdE0PbJOsUSbZp1LGysWWzdYc0Zs3dhULLHzu9J
tp/OeXeFemZAh2DQrxyq8OvmsG7Dlz0KA7q35H8b8B1vbWo+ZwkSmYryH8X/m9jr
DchVT7xalpb0EYjD/hxARucp5C3Bu1w1C6zjL7cP6cG7Rf59ohNbtfBkq6yFrNou
8r6iHC82nN1a6xClY6aa179OdSzl1lEVaR7xtRMKidrgSvhGmulzaenHat7HTWnJ
GKEoaTu4xtPB8sMDgcs4QxOxyQ/WVyLP1HUqzibmrnseKhhFdKCs5fAuJ02XbCIT
h9jrxzjO0mZOSavlp9xilWqHxkHqm4FqS13nLCqmk3XROTemOLmpD+cJKs34uVKX
VTvDqItmUt73MQ9S5WcuFH9KCHOcdPYnfrG8jvcB4YofVAAWeGXGoQ/IHl5M14ys
gCaqvK5zYWNkCyNgtEAinTQGuWunhEBYTdfd27pVjTfXcRBYIUPoJv7UzCqq0sQC
bsoekSy8G5aNWcb4BAtQNBTESyKlgYOPVjiDLu0V9uOsSpKbE5a0DIBVo/tw/qLQ
qOKfyet/1X0tfES9n5dySZdBbNBZbay0NapkA19QRhSXh6ond39q4YESBFSG0o1L
O+j6LjHlmWRJsGNzSGx7Tce2z1jcdMzlLhxubZnas8ZRzjydr/k+taXfd9gQInrv
9275oIT6yynlwqEaIsgx3vX01R7Z/LltB6S6lUbWBPas2lYGFYCUsIi5vylpEMOj
j5AAp++t12wIePOiWQUeil20LcGhw0tgurWPPUpp/c0edxIYr2LKEuXIHQburtip
WfgS3Dtyl0U8BB/gUQoHA+8rifFwYmEFERNKIHIUrD4E4s5Djvpy1nybzYiBegRd
EZBpuRJqu/1iRYi+gkHqPZ8ahSnnNO3QwcgWLxy9zJBDaxDdVFAAtSebFWJ5MmwX
cnP3GK8TDK1XmuT4PPrPu6JLGR8a45Fv9hOhGRZaAmuBTFT3/M0CiU8fRs/M/kFJ
MfVO0HN0W8du4ZdRz9LZXwc2lCIvfufuOv98ZpygGHWSJcNrca7Knf7RtDaYwGd2
X10Cf3mUiSVqgqV7eYzoBNfzUTtW8A1s5UiIYpNe3UDioYNJHC91gI87L9KJUkwv
RBsM8F3+h9zMpNfMf/6fNbmirGfNIl70E4Ro6cLGIJgKJSH9+xbsKYZxMwM4Rxe9
Y8QaV14rNYb56ruaKDGqNb9nMwLmlR2Lt98JjXwy5d3RsVqVKP1LQ+U3AkChZshl
1DAoIsPAAGTul20wwrIS/qo58mtOAAiRu/inhY1FMXhDJVsKop1e6H2sWvLgQfea
B0vTFkpS/JxiABu24AohY0jgvsiTd+J9liAmTezDiMVpvj7tdmBgT/RTuv0HieMG
BbheW3MUjZ9Ih8VffmQO4hjH6hgO1g393bGHuUtc7OnWKTWuotMkQ63rc/UgSYTL
YXO5bq1r/+32rYTRsi37v2hKvFBiKOfthl7zNtpcNwJ+xKBlQiXZHLl3/kN+HaGh
FU4ydobUIxEmGuIHbpoENqUHnbwB51w7GKxjrqCSblgI1EU9JVQrOXdRzFzHXcrj
yfYpHwD1HAqMoVpAWQbZTlAI3uSss2aUG5XKVva6WX5+dX3QXULb8ySczTO+31kI
2E0nJwnNirl1ADgMwhP2UZSIpfWh6fnF2Ikjxn1uVFPPYjPe29RCzHlTVozMvTR6
9IywI8g/mU7xYBnX6+TJMiLP4QwwudJuU5XBSDN/D/7UE77eSU5Ji4P/kG4XHVm2
27CJp/zXCQssoONR71vImohH6YLCP3A/eB5AqSqQxLLbKeDLqR0BwJnUQcSSUttY
s5mycPWgEphVVFjtFtEE1mdpgXC5X9R9/OTJdOBm7Pu15ahDW/u8VIpml1QtBIuK
Tto27xDjVcYaoSHmTXMoDRK/2sLkwt5U08sNjhbWT7VzSNIHTwBvQmae2rSw98Th
EoPeRRfxpUhZWJCnLVVNACfVPhJ/8bYMkxS1eZDzxKOuFGTPSDm5uiTabPbPV9u/
ws1ScSN7CRIz9bpdmI5y8HsJIjsEbxoZ7jp+lEiYnCzssH74AHey7SVTdNOSNaTN
dGTVEoj/CvylC2h7oZWEKJbp/pZPd+g6NPNd4ztzM5NgBk8W07nbLdIwUMjSaLGD
RUd2Mm+vK3RLIUeJZ8LKR26FJ2DE/w2DQwMeL7rirgISOJTSLx7PEGN8wmvP1cp2
WALoWAkjpmrddV4pyMFlhodyVvR35mw2FdoF2FsILCSowU2s1DsCX+UJ9w3epv9f
4ZvJIA6hRnlj5jG/e4pEl9JB0t2BnCabNQH6Ebwpq6CsL5bcMywHPA76StGBfyyy
o/6ACeCRwinVgm10VjATBYfbb0y9pcLgrJ32UHXGradUuz3PGLcfcrais7T8Jfz8
I/8rKfcZQENmJ36QxvSBdPv1bhavhhKXD/0CrqeUrcwLJlJvvXdO6TOo/IO9G97e
HYISwrzYwRuO3BWM22ej4ACtFvk0ONG+tBnaBb6hhtBkPiclsL6ju49v5y47+GlY
NIC9hwfRezeYQvJLYLIduMUF58+C/xN+9+MNSLhuwz2gwxt+LmC5B8vPgQ+P+5vN
r5LLjSyTsgO9srInB0OmKyUuuIX5ZAFsYY26BGeNZaPN0faK7cOKPrRViVP1IVCc
x3RWmZZ7qU7kvUemPvZMl5WRFjybJcnkXVZZeyrqibGRo3hIaR6zWMFzH1tl8m7O
VksnxEibP1lKg0qaAmwSFIW9P7T/OQRn0/5k77/efja1c4Fb967ctFf1XS2zZ0xN
dtN67VY5t/0g6Ltp0DKLdlGSfbg5rJNAFyOUA02bz4WjoM1ZGEyuXb1mqYox/meI
fVnYTMHyEe5vmeGMeAvnMIkkq1/urT71KfWw5ClhcoeTOugnahaSauxrvDR1XzCY
uHi0s7oJdaLx0tUlxbCe8MgzUlsDqClQn74oUBQzXbPafKTv6ppopEnqr8FyEa+l
rme81SNLr39kTAi7yAiM77yrhqU87d13LbtTwCu04h0CvrQ8XJOnFABLeTSfATOg
TDtLqwowBzEa6p8kZ+amKfaOja4JWqmXb4co7s/rUCCzEvRu1DNR5ZNXf59s4d1m
HOvr/jF60pMLRvF94MprZ0AbzAeIS84FqtT73NkovGmOem+wzmPD2dXMxGaVjeFl
brItddqVWUQgM2HGK+CdVV31Ql7Mszj3AoO2/w5QwYdpPZ0Rr8Z97jlh37XAbeSS
6vxIEv+W5fQ77PXrmu0T4+vqUEIf4WHHvOq9u8IScyvBgXSJDbckr5yZWekKa2KR
Gcoly97SsvN54ycJUyky81q68IRLsV9GhGdrWeTcdoUM/M8gx3Amx+9RaerQW6cE
jkLkgTqF/FS0zrqTCV9slPkCeSL22maMH/IWp6EwvnMbM11xeChS5jATkhccVqGa
kCqW30d8V7yU7K7ZeAmp+CG0qowSqgg1q2XaNV/uBk6wwfhmLzNJ1j5/YyIzZx15
yR455RB4bPZ6HXh+PEHxPD4uRSAJnZlHWjxB4z1G7rE27JEYa1iLW+9IYyC/Osz5
FjN3BrbCqdUBqoBZeq53n+DFaahCbVgNEAMoQyRUNxcEYR3UnVfGHtHgS84Ol72i
xc8rDr4En08DrMnr50lRg4lQ8XU5G7+T0toQ73DnLfr4trq52XL8a8sX8ZKBug/8
OCf7oKXat+Lr5n2TN1/KGyG1dZFPfLuKS6n6WJwStR5MYD8DX2cRUo0sqpdY7mDE
OZWqJYhxkFSSqSKKDONnSpjX6IMltFdCklTc5eNl5Ph4Z2RqR/Ryj1BX3Fp4PTHx
bw3Bqzs6s4JpfGkNBdtn/c7iUv3YIZheCWgMcqtms77kA7nlnqwv+2XvXZH0pm7H
azns+e+V6cWAhDoRUj4f9hb8ZKAez7NsaB33cYiRPtxIYSLPO7Fl9ScZFOJ8EAVa
AhUgfX0yNKxTJr/a3ZHKOT1ooBpLBzjm3hrYHvjhOaaWb0419zrt543J/EpjpA7n
NzG7i9r6rpt833RO4iKlO91WiN7GDXRFRZsuA0hhnvhsLbb8lvlhwVqSgEYDP89r
MsH9LhMyM+Fwcx1V6+FeSjkxxcQ267oy0w/EMkafPVJIXVG2amJeQSA5LP8hrKVc
FfPrsCyUD/BFNVfCoPano7qdNEFfQlarR/+X0kIIpRkiTNMNmju4HV10lODGcbeP
kvxD3mS0QAOIb8VoChxTWNElidh+8sEV8rQq+5VJ6CmgrOGW7HWsNvBVTK0hUAYw
Q/YKL/n+dA6RVuru0ViF3HHauB695UoUSlCZfI1ZOZspcMczKGd+ahB+2eq4L3fy
5O6bJPNLrQdM+4CUmNUy0d6CZ6PY1uqMij2IKdEOK5sSgQTRDVheyjxctU1HVghN
B5QiKD6rO5lUNgFFMrXdtdRGC01UOLgTrk5Gkq28USvpLaCGiZposvFIzatFb6gw
1Op0GAyWfY9t31PQ2MvykLzVKR5tTyzY3MTP7EwJiG+MwhtN5T+jrfKest2TNfba
fltQWxRIIe6AyxSHduWo4hOA3FvENhPC8gnyo7mi2rzRetmSnQ1y4vnSpjAhLT+5
m6O9jPAJ3QncCjkDDg8kw6mL7vByZhuIjfhIbr++XVW6p4akmi1pfpezIvKwXKUb
LDt1/C6m4cSe9fxaVidu6wpc2qKbL+VUiBWOT87WC89If3ZFQTJF4u29CuPDxMJW
dcPkhwM2Y1W4rhrtXyxx+0gBWXhQUAOiC/fzpYOfricm1E0lGpA5qfUMiQHFUInB
HYt0/iH4DW8pyypnxPI/l/8ZWdoJEWQ5vMZSM78+v6FgVkuwKnd+zauIMupaUTiB
cGh8LmG9YQFcrtwlZxdTHHcWNX84lYfZZ4h+5CsFMlYFMdJ2HWluEEms0dUixe67
cCoTbmoCmGqFUevaArTOCh21rIr1FWmdQs+rQW9ijVc0aZdbFFIPoL4zbh0ENR6M
umKYzZPQV7xCoqllFjdvTGa6uOgJw9IZwy70WJh9WjU6qZ4SYVCH/kmxyL394kUC
2O/twOS0xhodPxtvjKGhTkBXCax4oKVpozmp/YlX11Tjyw7re2Dbx1pnJD4Ff+1x
DcqEAP4mrNd57MTWsWBBYj3jh+8FzhUwhjlpEdyalMFPTf+2qVhwwROR3SdtPS7g
cK6z4bS2VoXiwBYguMup3q0kJZ/W7Fy52cc+IFIVY2DRHD8Bb1v2nvq9M+l1gkPW
BICEbjQdBSk5ll0Zhn07bf4z9MAHgAeBaVkf2sm1j8SKUfy1cu6aWXKQLBSnxY9F
qK4d1FPyjelfj7LB76xRqEd+pxr/PvDshB2y8kcbs3d8XL+YxzGLnP1KFPhNWvs+
/UE/+c04P9WcQLJnAFBo7ribnXbH4FMZ2AjZFAfljJmE9CSnIO0oNosIj8oK5jUH
jw11x8daG91m7jn528+fJ3365ORGrAZcixBVLeFi87w9TLmyGae9RFg8pBwZ5FnK
DdU7fGIPcOS/bbBnxWDYvtUgkxxZH0zSfxSG2M+6ZnkbKyL15FI5ohh5L7TKdZbZ
vCMZfzFL7qFOHHnbOYwNh5x+ACHznJJnAXz2HQqKFOKAtHaXBKafkZaRS1fFfgYF
QuDima5zhFdB3HL2HqpyYeuSGtd3AHBIkuOyfaezVFlurLN2W5s1z3ojVT9wHnRM
a9l0ggZ7piWwf/b3v+KQLBSItQ4HEftOCPiVHQGvjzO0blXbNb9nj1O/uf6ovNxV
jTTpvw580fJdCh8iKtD0bFlZNcLM08DP/BRwov1CKy02mkKEZB/ukFd9EIsksloT
EZkuhxguPpm+KkgH1C+QptWqnyfK2AYkO1m7CCyw1DoJEgpsKWF9SxTzpKslRLZE
QD6ddF/w2NQv38zNsKD/Rz5z5LzrLiqSRXUJOP3kCF9o4RP6Yt9Zh7VLEuWHftDe
xgEIh2O769uCg9g3r44rJDatDwTPYFLbKLPGXn4f8QblWmKKPVdxSlGReqrvJ3nu
E/XYRgdVPzQcz9V5MXP5GfEeMJGizpByoQ9P57J87zHgRhGDaeK5o8g18deMkgQq
yhdRO4VK1D/u8bCG5N4oJReCsflmtAU8PZosW1qJXU69Gl0DT0IU2BM1DSnKeyYJ
ejUsOl3IQN6LdhvRvUgn82pN/wFSKpvo7jbvUjs/Kg8Kj7zLd0Of00iqqAwa1US7
ImuPj/eMvoM6DwJVVdZzMzP8FKBzRMtx2vzqfmfKSP38KIbBluJMRw9u42MrdacZ
gLTlwl2EXhMauctRTJqHqW8bxolvN7EY7ApcFlgpopEXo1dMUad0DyGBAoGEQ5ma
9j3yMpyDZ0qHzcrKc2wxuT8Uf0bVXfGl8LAYXWYI6JCwu8uPZkCJ+R1OtRzQA2qR
Na2osYZoOPXF57V/URwmNVdvd+WK3MgSJR1bCW9Whugi9dvuQxDK1GmRI8QCfqr1
i0uDi2mvV4BdXbi8YaaiH4FZvx8M55sJU+8sSeaiT4SISFOs/vXSDkiOP03EiF47
SKhIYR8IEjh/bPpnY7Ftz32XlEvxnlkAv1kTBikdShgwzm6KoSVzbjlId/yZ+Syy
lN1Q0jobPUZq/E1Km0J1Zo5h4ehei52KAfr18pMK8kZPOQkzJkk7N9F3rX9VgoUm
NysGMi6QJOHUw3RVrOjFhTb/OK98gNJPPbL4UxH48s90Kj7DRCp9vOdXmMpKajKB
TVV7ISNE5Iqxuasde5FAxFTuUz8Nz29lH78km04kJ0oJUjDIRbXej4DJb5DfU3h4
umIOL+Y3mpfjT6xbrfuAuL4E9eUqpjkK2+jZmZ/CURZyCnfZd1lQzm9YjCBQ5P0r
qljw6FEE97R7lYOiK0kSEHwWFusXp7hc2B06AUn893bJf6SSrtepHVIylapQZub6
0xUnNvRvBWYDUSiB4vGLkr7EAf1uZAPBz5/H6wg28Tfbkdh9jWZ9TfqHaBf+nDz+
d7c2gJEFymSXcYHCIvG22tlR/aTH2YY4vd1LB5XxtWFw/BOLVOHOl0MNhp86stID
K+wFEpqF9Yb8AAf6tDORdkKAG/GGtIhVGWDAOqVmI7yRh5WzHxOvfaKbpdBfHStB
hpJVe56tj9nV6Y9Av8GX76HHHMwrJ0mwAUmASyWOQ2l4HErOeUZaKUNt5W4MSte3
PrpirmfoaA9dwuOVXMPXUOm1G6Lphmus8xP9IrVB1NnJyeJO/2nBASmBm6ljIa/4
lY+dvK5OypSoniP9yOpQ/i268ymC5zUQwuta1TiDLGXZgiE4GOGqRskJCR2RbmSk
zLbpo3dZBz99Whf0QFfjOKYPnfGNM1/kk2OBVgBJZNtTiYSmRBDJkBL/PHTLQZv4
HxQpEZErmtpf1zo7Z0C0kVXXoj+BNS8qVcmb8iBHLCaewHfKI4veUi66wOAWOYF1
C3YJ/b38SxNx8k3M9HIlb8Ckt3nsJpgSRiypjkeou6XGWirJvTzoGYAQqHUNBFEc
USg2nxwRhPu+82ImkselZJLE8vJGoSlMzhTHdfrgQqLnt02vwetwqdcXoYP1IbpW
YI+o8uPlc0Pwr7dAGBEFDgXQ0NCjM1z47rdgy48D7SsciRcagEg0fVAR2NVvGBBT
ZqbaU5v6hd9DFew+xz0pfNRu1q08iGj6S6nLvT+q4zx2E0kEKjt4dLdjuR+tI9EA
bLJ69FkskI0x4iV56YP8Sgab+JBCEnlZFAXPbsmZ68SuvkLq5kHqbSLz55d6Pbip
kjeqaHP6XJu/5etyVRvYNtrtSFc0PM0gJIiyfRkB4b1/lv7KlLgY9DuYBm9jD8Xj
vb9wAJcXsxZBRgZjUDXBpRCokSShViGnOhl806IGSPEBd9sBL6GjX0H3sn3/PgW+
sAOLJpX2aKhSLFY0f0EVTD/Bl6kcruRcDi/aYTfYyC+aO3mJ0fW+I3kl4BtPIa6o
r8rITtvEk6wOlyNWCgPaUlt75buxFi/ghQkA8UkwhMfJ4SlLbVVEsGgd4L+PBK1x
UypalRUtpqks/HO6M+6G745D+58L2hwe2TD0Ku6sagtiC1MusLNCwyYDl6xnDkBZ
QDLZFXSVfud4NmTgV6/fCQIXJn0mPqJg9uPit+ao4OEjAfGmzWSgJGI8/e3q31G6
kGDzcprTFtXP4tYyWNS+RTZqgGXMqiuyj5ETa/7sTNov1mau3inPX3uwhWI43udO
muFmpTVdQPHqdjECspI5IYJ6Y60ssSGkjOBBqi8J6WdlSVKmIbJ9v8ixzl7WV3+H
tZFuWVkxKfh3Ya/VR3zSot3iz7c8oXKu5sNXMi7BcMHSjo2yjE4EhY29yzJ/88hV
OEd2PB7Fq7ldJwxFokQIWqPiQ6cHY96hxebbBpaCgK2/Jai8qJeC6Tm2uatc6BkE
2y0NmpUcC6UCV19juEHzr2tmFFOWgVE9YiQC8Qs7IlfLKW2egXjCWQu9Dw/20vJE
hR3vX82turtf5txnkGZtWA4ix7WAerHJXkrVM8wPr51aLSps9czR0VRjplhdcGOz
hm9bIH9apeLd2loRDBPecluceamJdLTRrlu2Jj9gnfpKezegzsf4a+5kYeSvCL7J
NGlEHogef1AApjsR+W988IF6LJa69YLUdIrlgn8aonZY2Orv/W7Nv4duwWGOZWjU
BVhLuk84kk95FT/14h4IqLhA+pZWyDm9zjzGk15/EL2NAyyLhJxZnSkeABl27BJR
unfXqs1WQnqtezdu8G2F6HeNYE/dDOKDBiQhKa+FyTcw+BOf1tsNW7k/dkR8dtc4
G/i/yodWWMe+XRWkmpE6Bh5YJgPPXzVe/SRAwl4o+lVp0v9pXPNellfCGeEITBcu
pYVZ7zlTzuaTsDVd/T1/rV892ODZx1GLZtNQnNGmgsETxRXcQ7YvXJy57ivSD1TE
RpOZakv6UED0Zq27Y1XACaIPJfgLUHr8j7ty/MfasqSR7A50vCIkdNXS36tqSoxG
kagMRrANnWdx7mQwK+8Vy7BuCGiS846g9B0arxTI+DRoP+nax+dNeGy36Spbh4zS
gxFrrAaFDX44Brd4fkj1jIjAwegIZVJ2kooJ4Ae5DusbuvHWZKZ8C4lMplcmDSjs
kBJXLU6jEKrvcT8Bmf6Pw6aVyl6LeXBMpALSRFPSfsL1w5iiG6YQ8bTPONXyv7Z9
BQBuUebuUZk6kHeFv59ZsiIA2Bc8tLkJV+jPOcVuZ0Lvk4vo68EpIkMsLrKJTlR7
wg0N/8B+Iuqv1mhWxGWiyke4gx1XqX4OfZQ284sTRRsWWy5h7n9PNcs/5r7XSTfe
vD+uhzJq6XBM7Xq/DubVkcL6td3ZIPJLDBNBPNkky1yV8VBIxUNsSSSWT1WzMpqf
tgAyVNyR3aQTSUFjJVd7RfnG/q1szeJfvI2PZbSPBH2lc839ubrPLssIoMoMP0P2
8icVJnerdJl8BcDVEpBR8tlKkdm9lSOhgI/juyIUbODioeL1+24xgURF7bWSFFpO
qNGpCUCnoDf8nBgPgBIj9fWLO+I4qggSizviVPOfeQ8MMXVZdGz/0/bi4cgVrxi+
VcDA3SbHjnRmWYpaIDdHNUP63ZU6Ped3ASuCqnwycBBy5DC0Boj3idc+po/BPH32
9z4OMFTvEykcrPskimARHKzC7ZO2r8ZGs4j7cCaQchKvMdDWGQrkdbn+U2GFTTXC
ij8D3ZVzJz5RDNQI9Mwvre88fDHfUm/JICnKjwTT7VN987qPPd2Mau7Z1RHQ7whn
eYs5DplbiOzHG0X/HQuIrkyuKwqD3o/2gDht3dRDk5UQeFREa0Ol97A1eiYGmRfC
et/aKubd/ZTdgoFmLX3pLHV7utTSAfFJ0DSngdiG/HIcIOlye6jHDZqbrcrDfpVq
567uLc/7nIgoOOaLfHwPd8qFCqNe9FkdQ6OTimMaVCej8xUwskY+SLIFjWfUxuQp
awJjEyJKX18oLAmieJpwQX7TU4RvZea2rwrYwl0UgNvjjqLKIy6cit0R6hhbiEIG
5wrAygYRKxBpQBlJiEgyIRLS8v96wQ4/45STgajHUzdguwECZQfE64ti9VKhqdkC
2bw7Gcg/9jOLuhALCwjiXRbtU3hflET2bz4O59jAUhfTanTy3ymfLoCiZpFZ/q/n
l0KWg4/bhOUyxBE4sVTtvW6VxCATvbVV7D1N4MeThllV2Hv9wCoDL/R/NvzEjQ40
aNgIcJrqMwpzwuQZm1FWrt10Ji/P5Sp+cJAZroLQlKe55xAQzWb3C77LVRzmeRdf
zProloWB7kvFVlMCoaYa2HhYcYXcUl4EqsFX3GGDJwdBouW/XJePfVXT7slYgpIY
fiuk0neX/o/Y4bOtsn/vEGnUwKZ9xDuqzyN69CmV2G7YCN6QsUJTriYQ2PqKBu2q
IW07YABxPxntEU31lDSLx2LsU9S88bhi8t2ZrZq1sW0LWDy0G+72UUgiNA7DAH3y
ZosFpufWs8yMbg83W/6swhkwxurYqIRj2TEjyQpnNDtZytGwiiaIPxBcEOyObZhi
eHsvTWqQJCbz+1QvVL1M0BctPBLM2q5sf3EdxGrTuBAQV0MP90TZLItRF6bYvUVm
PepkorccSWYkTC6gNxsnMxEdCerP4pW0rGSTE7KuKuWWqK38ngiEj9N0W1PmRV+R
ef0kI9R6R8oqcvNu5tUxbc+Z0x3orBqVeICnKjma305RvhUJ1++JBID7Aku7hdsF
YZs0vr3DJb+FhbfUU/NmlfnLFLwAkG14K0dYtC7pqFOfBF80cYdIuiKQwTDahJrB
vPKK+K3gR4J4AgqW4TBAw7wIEo+Jx/a7fPFjNveoOIfhqf9hXQt0yInSarSeSX69
rJiKtlHCTXcA9/9xy1bRMewJK6XfUQYRq/2k4uTNQc71XtW2AlWqCQ9WHDBTVvdD
wtYf5Ted+1GoWQMff6f4vqWrIhkhZfVnId+CG6/dkMzDQJVmeyYWDNV6I8hCKa3C
qKrwW8UKEHkQ9i66er8gMrwaBmX5FodNrtyfpr3qJQZH7o12d0kf7ZFvog5aTX5C
imiRt5lr7C7EdGANUtIKZbazAK/huv5ZSyCzEc6HVoiWMkVUWVPNqttRqZCMr+05
dYoto6pB/6XLEu9YNyX2LFC9In0V5fl43kSz5Ju2J8HIysdOPmxDSZhGKiP0RPYy
QIFcERiy87tbERMmrRT4CmL+ho2csHAAspjv1uw6DMuUQGJ9bgkrw8m6Fy3m5SSm
nyGMSHqtnWUZR0XU7MEvkEc5u0UPmjc1lugBCwIr9hTjzoTjC6DbTT3Dw/Hh/I2L
5my9xYE8kBmCsQdsx8UcgDZF0DQE26AaRnTNyQjQLFjP18bCzBu3xY7XRMIvDpOW
i35BdMAny1D2zA9m7lhygunrwsT2zC56eMP5oPIuvHuVT5GWyYBTDXmWJOEpElYj
yS2XGAVbpk6xAmiCgk2zxpfJGlBpimXv0LjHVtjtN9+Jzv6St4v0rZMJjJ1dEZRc
3mNULsBQInXZtkauZeOlBoAWJK6xZyKadZZf4xTMjN7XWw+j0xr1vc5y0M8u7lrS
kcORw6z3U51X+aRBV+bR3nQsmufND9k12JCceEzxXE7GB83VWkHh4ThIrRfWI9K1
T/dERzWIp4j2tSSrr8iMds0EvrJWHzhcTlsGcbqLaA/XDoJhGubQVGkGUnGaoxQb
UJHRPG2+ZexW8bAqzINMvRVXVhlmPmj/haYiKB81l1Fl2eeYYNzSDhZyp7Gv4fFb
w1UuqHn559ESk6bhE46wkgHEhG0/Z3QwI51lZKbkVPha4UcyT0TQpfOvfWR9XkP2
prp+agW+BD0bdQdCLurJ/kBOJpatoqF80MUqhz/DKXEic+5vUIpD/gXiJ/s4I8lp
qhdXxqoWBGyYPirlb7JBjnH7cvvmFjCGsbI5yYxrNo6IU35wTWCHhFxsWZdrOBiA
D4oBjWM6UeCDxDQo12+jq7qnLGCYk9MbZlbc3I9clYoNWnQGEbe/oV4jZ0V6ImJX
elvSD8obr7s50aj7IyXkY0MdkA5S/nVchvO8wwg5jKU+a8JkNJQElHCr6LktamSI
S6Rvvl1cHrmwx2A0ky0JzC778G4guZw+TJc15YMDq/SiYWnldjqfJvZm+9j8V7kj
h8N8JEsG9k3t4sA7Kbvi+k8A7k4e2oeXsh6KVQCZtdW/i/p9mvnNaVNQn02bi/kk
iSdGZA0zcm//jWg/F+/f3vHuLDXO6fcouRvBGAHKgzYId7KDbLmYULHOw01b8Jgz
zUIYAfjmwzPRRTKX0H5scPJVHzGcBYM0EW2+VecjGzShynb/SYp9eZ2QR1UhQvru
iibhsgP35I1PEHNFySocFhFAkqwZujMFnYI55G56Y3Yvp/ZIW/VnxRDoEVhit6p5
IBcZYmTl0ik4Dq//bU0HnpQuA8NYHHcv5KNsvnWW0U955RMNUajyuEpRaIpMVKks
5HufpRT4W8HiBdDpjupkm2xcEYkkbKSGaLB9SFFrTgK5t9UkgAw4vrZbgtpkjSfn
W0raM+EVIc2qpvDZKttfYNyxllBPCJSXPa4RdindTUDAFgzq4uyC+JfshXyTqQzq
OCiSSObxb2zf4oFR3ADukflMsBUz8k1qXe70UdqPhosSyRtn4FCudbUOW77ji3IU
y+eTfZox9G0X5jMoADtg08B4WN/Zk92OZiBtFsLIs9MA7Zl5fodK2IdMh1SxfqIy
hkUs2ghz0z9d6v285LrL3nIXzG13n1puETKDKHv6jQJGmkc9L1A+BTAuoAunOSbb
A2wb+xziDuRDEh3h43vIoYlEdnstZNHCXk+pdpmtRzpH2fN2kXoUWJv4fSWGy3mE
CWCABoFkmtG2RCmle3nUBNifP/74iClqhYtCRTPLaTBJHBi03DdZrREXHjIe27pS
dPzPw2LhagDxWXruh2rpIrKhX6K2cDGwwA6GOo6wFzlYUtxZReKcnJiZqHUaOhUE
9IqbXtO0RTnIhGVuy9U9E+zsAix5y0KdGtkbgH7aURj+YNKmUPbfiMkJkPg3Gujf
Ot6RUF7HuV7Uc+QhEeoz2AKun+4OToivNXxmUF92ERmLTI7gnZ+7hU0G7H6m7/XY
L4sGEvssiJdqOGIpFK2OzcM9d2F4KsJpjyYR+fR218X4f2svqpfCpGGgD2K/Z55P
UVmODjz6dQ/aZMARl6vR17gloDJvC8N8q8P2vsB2t1j6OnoMUG3q1olJZTbtklHJ
m3P1bKIzbaWXGeR4IzrOHmLBNLuu5uPoLFuWLxes0cy1YG6W3DIIdMLAY6Gcf4TW
dsdZtfwyAOw/KsqTrwdXVmW90eaTMJK5S/hlg0TKREcMLiRweiBR+SHp8zsgxtwq
zi3tvJQyvxt3eBG7mTZLZBBakXeS0HREQa3rA7HNfwUtau4XnNM+x/bSDkTKYZFg
dKkvH//OZYZ5KVLFCeL+GtX08dqDKLBTMPeU9W65fyejj7YqfrV7dUeUcpnSVx1c
u29t8Uo8opv2X0ITjxTgJdXrP1bDbiAyFIis1E+AglfDMKA2c4ykMjfOnjOlzEwB
qC41vCLEi8JEhylG+bg0RGFD9eY6SRsIgOsxXyRiNqmijaBMNUCvGOOVIn99niE7
AG0Yh6Q2bPGsXMtomY77lyCEPOnc/EAQO5L8lr+eJeoW2clYQiJpMH0AXPt0ZvxN
QPynY3TxWEEL6cZAadctE7x52MnVAl1ROzXDTV/N/0Ximr/NlKGzB06r7fSO2qZD
IT99b9DYSKNTeJ/kil71fEohrLL2UWUa1pMXftud0XSKlvzSeERWh5kQ9Lv9fbGz
XWbwEgHjYqOKH+45xHYG7Textws1BoYBadJspHo3upJ7FEx8f2g7LJOvlNl9RDWt
hZvsHutT8pI7soaCRY6OuRgty3YwWdTAMfTNCsu7v8RpyudW/kknPVcP7v4O0Z5J
lZdGrg6UGJqHvPKBKTG5oAikU8kWYCxDF8YVjavXZEt7y1DYT/bAADZlg1Dk3TBc
nyZV+TdYEag89vQx/+EbwtbxnsK2N10BpKuggdW/jBI+isS8Ce2RzgAjl157Ilx/
j9QurGHd18HVXbxMfCydAoRIT0I1xI+QmfiTvsV7CMvT3MCG9WbTsjdri7I3R3n0
zqZ8edjdMmEqNYzw8i0dGd5hsXkIWJoplznP+UtG9u9VUAlV8LdsNZrPY+KREzhV
NGGbBBT9+84GGOnVo3eH3qcaaQZlzEZiH4TpYE3B2WZJ3puI5nm4YR6ly+JfQ/a2
yvGT+0MtNSsQAl7+QND9KAaQyWk0Jo07zJFVF/kMKz4XzQmDpo7xZyUbu2Sdmyx9
QiBC15oZJHQb8rOWgK289rw+ZwGwiF1t4uwDUWKuztcswxBYtK9sxAmqifwhe4m4
U/LELZB1MgVLMecLwDhmbQpP1sPEI//ZAPo6aFzN+ELSwxGohlSYBMzd7IOLk6Lq
0c4pJBhzrjRcSqVbRSuTEUtSO3hN5geYq64mZUmPvI+Vu14wLHXRMhp+N5MEiC/W
Iepn1OEeVBRtTTsqvFqTBLNIuGn0gNObady0MHIzK9j4Dxe8TwYq2W4/P/oKboWO
B0ASBXsb+YFf9/iZk3mrUCdDAoL69jm2wMSOXodEJWxI+wMsl4bXnz9z2FoNek8s
7gS975JFF2r7CG7+e7gbIQ+7aLUiAbrhQ4ik+ww8AEH6Bd+ZnINJF1iVakCJtUVW
O8VhD1ryjHeR87kvB1UyZvBYPmSBDqjBxq6vndlhMlxc9iPAoY4XMvyGixSW4/tZ
u4sEl0C+q0KurGiOjOaWw+791auAzgpNw6tqyWNznG88iGeWA6VsUtkunH8MCIcr
ueVfvL6KR+0k/USjuQ5G5cmS+qpN01cJZJn5AfujKsY22eisBp63bMogGJVETz5a
IHr85QcaBeEqXKXauhlfHJFMfszyWUfyGOg8ZfF5M3AtLReHb3FSIp4p60Zq+0GS
Awt5nidYTUDA9Am3enUapCSJe0UAPsgfnlQtXdc6kZk9FoWtyEIwY2Fm+YEeseIn
Z+IQF6NvThDSaXlucaUbpojWXlnu69fYRKo75cDX6Xqgy5BekVkrdawYlds2RiL5
HlReOpAW4QuyDi4T2/D9kJq7sSeOUVzns7v/vEs5PM9Nj/MVH+y7o8R/HqjI1T0J
nIz92bVLGcxzCVT0r6GpXbrMMmoXu7bYb827V6B6XMDlf/cW6RFK0+pWjPKwYUSn
vrIjNFLD6HtvSquE4gnKnxWMgd8DJ+5n8m7fEe4AWPGb1Sm5pAUnwuDPrFUInv70
UVqT03gFe0yVk6qaypVQbYLLRHSw+sVVay3GLLi7lEM2I4Xy+N1v4zfxKFoKyPPa
YFcLL/Pf+k1MukD69V0DcMW2W8kfiIT7QyRAH5T3R+vEPmld0Pd9ZraeWc9mA5uV
BmuLiMkPHJPlQfuotJEPXF9ltumkwSNRWQ+mOC5V96pH+7uonv5utU1m8eByx/yy
0kbnJqOO5ivBZJYNmkedE9YY+px5989Z7+Xhqvx7gVNYO6/wHexevpDJK4dffzWW
aPVC8bsEHnLEzGOXHu7a1QT/uxjEMfo6w0/AM8E63eF7R8RxUR4n+j2V0wxbehME
Y1Lx8GYZ0T0TgergvKk7OBGcy7y7KFqbXzCoXSpKR1tC7ovb+0mwJBCpuZ5ZW13X
jSjhfFRFqMmOcG23nESK0aqy45yN/9ESnNqv4YgXzEhAKuVgheM4Z5UVhfeOqN3t
va8ASwqqdV8z0Vxoqz/6mgrmyMI2Fb6NaQNDE1lc3nXEtSs7SeLwVMkkVBfOIB1a
XUAFY/TnnvDO7wKp7DzCWFe5H92EsTMELkRoN86yxfzRH/xIJzVwoEaxK8Zbs/CM
A1M51tfrewtHM00cDtull4ne0iUnwVLx9Vm6i6GAhMN02G2DQVZ06paD2qk/Px4d
ICgBOh9NQJiL11cSBT+1iAthTMmkHeYTDhukI6qbVsrCpWGhou8hTk/885C1ZtvE
I9BBYzzqQbEr3osLogdHp50anzK1HkHw/2HXCM02S1A3sIGs73NaT9ZlLhXkyhvI
ZplmB7kfsiyfaSx4JGWLIul6BMICiGsaFXOEubCxo7KihTVIr0rzmRdvt1gWZeU2
BK4O8u9N2+uY8kCzgHkmmSxkHWx/y5rHT5Bt3xib4M7ZXpOfaRZ7Hof+6/ZGIjWc
ndACLu2jRY2K9Yne6RVl7jybaEEUzKL/gEDANlZs4IhgALLKDzy9KfZeeXUOSRlI
WZ9kF7Iwy8iBfSwdzmE25Z8CZOGThRhrPYx3f5LO2A1cT+xeRqk4ZCgqu0pTLhwV
z4HQPdZknymp0q+qHEfn0etncCWAHImXWQYkW0FgoBgpB/DwmxOyd2jHOwPf09nC
6vT2TC5msaeCgeCM//xRTnoLCHuClDZOlMqDpUsPisXkbe2rCRfmtFFTW0ZBGsTk
2EJA9ZcxgW8yGRGPFRDdGhLzsa4T8iYHapv+KULO1GMX6qsLUKKVr7W+KY/89hv/
OvFXySfj2gu9i+4NQ/htMg6tHS2zS3YIp3FPVu/TcxIWj/ntPlUBykStl2aqsYJr
o5TDA119F2D3o326oXukEyrW9uEomSVOlJS2RcRLGFhUEVZgiV1DTdwjx3ag0Rd1
yBZn44T/4pQqMGpPB9jiGx+zlxRn2Xy5jh9MzbNcea+SBqP0og3fhU8G1exk/kM4
SoPs6jCOlgFkZe1qc8lM6Wo4vZFi37LCCoZSR7aXrc7Ko0ZDqPYgZn2iDBjAV6JP
WGAlH2IQRmt7rwbPIDKynurlRbaP1AuDn2oirGV5k8SMv6QaioJyFXKMCgPOWEWf
E57Yj37PF70FX4XB5+1Qc+OxaBEbE9KWPxspcmwBmrrhJANzBPpvkXTAiuQaX81y
QfnQR2L6DvIh1Lr1Rt/2zhzwOdmQ2pL0cn4To+q9aU7wSc1h/B52icWUNcyYjp00
OUPNct9NfLtlw+6UR0VwJNt/DQac8NgwuAgUJAf2xQ4qntfYveD4tU2HOiOK9wa/
nyanQl/W30T16eaXDe0SvFyd5HFjB9BiAGbr44XQwuzFn84qnXEPp7xOy6Ru0ULm
PWA950Xn1qGplkav+VYQqj0mJkvZvy6Lcv1c4RYChZZtQnhlm+HnQ7rU/9WuKacZ
6Df1IU7qfWc/n+M+OTDjJvx7u6KUyP4CdcwYCILew2UPH8BIKefOIedxwI811TiS
D6h6yCjxoBjGJURe/ztX86+zIRaIDd8U3XZHoHLzLYtjOBWXWXug7T28hz0tS3dh
ywD7OyoQ/iwoDYceLkwn5ID8Io6uuvBDlkP9k7hSx3ySjsQ92SRQOdGj97CzDxd2
QLnNd5kBniA1J7ogWHS+EN1x+wHYaXEULsfsSaCnxdCo9P+fgCdslztRnFJKXSno
mWDquNKUzMbcyLVUkItYYnuGa8BImrutV0mX8YHCR2WlI2Ojh31FNgEorhJ1rfDg
FCGjSQBPk0nkluUZxSLhJai55z/f3sHDzBthHLONLWVEAeTRAWJrMe+Gd8g7gFkO
mfXS9GTdM2OQpDGxxjVv4i54bY+CL2co2EQ+DK+r6H1Rwtk3gUeF7rk1DGwhNOMn
IROtL/qYu3UgBnhVA1iRxGHjk49Krh+ccWGB89XUCczQlzxOKMUX23fo9M14WFZq
eVzYlgxXOSsIm3PRclE2Pzp67LXo/5v5hdgVVpnOdXqh7vTILv+ylVhCQo9IBcqq
b84dJJTuJpV450iP1ZUetIeba1Te98J3JSsYWyyqRfKzoZA+wOd7Qrz71FfssiTe
t5wjWlfUDdZ0uXUVQpMlqBUseyammjIVUm5kiScc8SQurRiNWRt0AAGZr0fALvH1
8acQjKSTmgDjOCxr+q8XWerHvmzJR5meueDnMERpryn31JgAoq7c627aRWLazck/
djEfqgVaUT4+DPMBg2MWQX3FcMNvqKp5VsezL27MDjFORjDFRJeXb8OGRaso6xbh
33M1cywdNM6jgOiJwdHxLkdne8SOBf+5afBQ86qxBale6+rjXz1QsLKu6Inafdla
HT04IGjxU6ZjZFk/zp3QXMgh+s12lYB8JVkZ6q4H22a9cr3ksp5wG+ltc9QIs+/N
Pt7JLXAIGFseMr2OG1J/U2uhChBlwtxvzBb9x5sB4UsARkgdohGZKPstEDOcduUH
Jl9l/tlFBvQ5uG8jp6tUriX2bVT6tP4ewDklrGYaC05bxJyyg1Nca5t3+DAeRaca
yRwlqqKXD2kguORGOVET7BjMUgaeVWf9J1GAbmXwdczgRnPYRKson18psbJnfYxU
yog0KA+motL0Ky7Khd3u5kOuSssoqRsGE62YUTEtKagTyFyoNig72pDBiXTd3YGG
cZ5DkVtnyf/DR6FyCXwlVcs6iCglDMsiRA9cpk0JQr1y4l4fH93aH6jXJJej5aHi
jYij51XaspOIjIpQu9yAskxfpATwtyOaZzqvLPDrLpEaQDbKuklWSFFC+JJhZOYS
/AabAtEYS+Iq5slLs7Ro0ZdVOAk50qwrUT5/hm14bcHApfrl3lcwc0dwXiwZBK8z
ik5N0wje/0+x2IcE+tgsCbFuZIn9pKe3aDg+ih8f8UDsnh0a0420EskHgm/OdqqI
ETqzCfn5LOEid3oK5vwh2c1LclBei/+/LogJLcbi24EDXY5ZiGt6JSO2EwPlmOS3
gkxI7gmmmwx7VgvTVXViY74Ypw7jxRekV/oJckhC5TOBvvbUL5stjPitO4ZShgjY
m5ZQU+zQzMCi8qCjL53kK56ELFe6vNaCYmzg8XBZQF3Pd8atd7VISERQhTJ3RoEo
HcLJejzh3FRpvoTVwxakt+G9CIOlIVRE5I+AeZeKfNPHJ2kyMdRBtVExkqT4BXiO
6shioDbhB++dRdjP/osMfGiLcc0hXfKe8t+rKKu70HP0ddPjy6XfbpvYXgEhi2o9
+lqGskIeTow1gOUpbeKeScLh3aMD4C2X2azb5F1GzP0kXrjZiRp7RnbJpzr+RWsV
eN5GCLdjKPRcB5oVikFLlaui1Ue/blIflfKNSGxQx3bkkapIfePbVgDSL3axKXUs
JZXdyWpADVxX/ng76zIgQlnWpNaK0nOY2Xnw0K6fATEkyJ5aj5GSDsvLiMd/5i5+
l/rOlCVXYfrjFjDFEPNS5bsaykk4yRRWKwqwf7DImFiVaCzV2FFpgJDW0yKCnmGf
kIrBcnxE4zMe0yzpTSosuHrkH+qqCVLANVvV2NZAPejSmPNThzO5LCcv+Kw9unbY
9MeUq28n3vZIIl8h92HvlubtiFQpnFReBB4SbFtPicbz9tWOmsjtVWF7HYhsp1LL
BF6UKOhv2k6V7BmYfaXJskd7Xu/OVoOM+VsUyhqWzKPn5fzM71PFD2a2A/O9h7sH
8uv4Q7yQ4Ucgz4Fl7Sbj/N6n7FF6b7sQy61J3BGTSKc0Mux6pJnJQU/XJZVsaOx+
t2eV0z/0JjkD/tVSVAype5mfdRfCLzJSbKnM1VG4kqX2JfpOxTW2hPexNQGPXt3i
qIvSTl6/H0z7r/D8w9lqaTkHMy7NF3NHvc8GisvHchkl0+zdne3BJBW9l4Wer19d
nA3i+pjahr7QpminEeRxir208tEn8OBrqe4IuBc+n6sPHdyAwhwyvR8TdTRS7q2A
wxWmJg2PEDSUGhs7sWKPuJkrkHvy8WI1JkhmEhx/VGauIkXIjO7wfoE4sHZUT8CQ
TUhJvCWvCqBb/6bUdh386t2ntQw9fXuTxVZODzIGNHnjnhodh3kS7ckYfOVqGrCO
H1wS422OabIE8Y+QIkpTZz+N2gD39dAiRYiCsgaJJ2YcGi14FzCoKlzwmqULoYfo
YLIAyL23a3IAXXd432aaYHcyIb8lE1y9M4FS26BLwtCnWXheMyM0yHuomlVLpL10
1y1ho/W1DrTTLXcpaPIIF3rgz7Wzl5SYgSkwOGFcVz4x+MXH0tYuc8Nq2h5QfcED
mT2qYRoPn47bv21i4mmsWjHfzzs3oexOt1imTJ3705bgc56qKDsj4Qb8VTTZaG4y
iBbXgENho3AtcezA1X48YW11WQSomcsZZmRnckuR/Vl+0vTMEXi+6VU5LSL1bif9
VAgskJgVwBxTAOIQoSbgEyjaxejv8Sw7ggv1DLFVMZKpmHX3zOF7xqwvNCNJ3qF5
teHmol+VFxpHEKgeHkUMGtH4Vkhft/PVTgUMvH0torUDDKxvayJugG49FEOOSdT0
iGYTZJl6ys4sSo3TdKoz8bCsMHbwdyESxnixKTZ8es6uwcJd2qWTYF71MUSAv5yO
jFikRTYFtzTH5YD0e8G552NekfCL0RrTfY1Czdbl33R/KCS2PbFLY/j5vousUCsa
xwnsqRGXhK1jKP6c6dthw9xIvSQLHrBrEk9YnhM0hksLoXHZrQFTiCeiupyU1Qoq
ALykE3ag2t3jscYnuFpmvLnZrBw8H7iCjc7vMOITTDrN7pI8iAPh4xASi+Ob5FAX
7rFtygxUyD0IC3b88sQKtV1IclpHGVRdzRjpuSZDTrtUfaz4ivPQovm62HCBYWPr
LpTjtoBVTRCJA1QgflqhhbaiAf4zGqwQWECYBQfqUUQp2Fx4y795CsDheF8AgMSX
93ZL8O/6+s1KffD70RwQmIazOXlYdNoRoBDGTta6B9JOwc2ZSoDvdm1entwX5+aS
j4q0GTQhsliOluoOPpX7abGw602G9o4l51v/U5BiOBvUWQzRMOL8JtO4DnF2Vx8R
hBv44LqIO+swfJexPr1/IKmckvk17W2esDplP4+Ju9GBTyz5q+nmMjPrRQ9PWaBr
/tx5N8+q+3vNfSlND4S8rL/BHrYbYMuV4ATjtwZgQAULa+s92ux0yrKzBFWI1piz
oECR9sUTnTxVj3ADmxObTzflije1YKIrWahOEiqd/AcOGrfsQ3zVyrt7mPfrp/3g
lpuc0m+CvjZhVwbV7x5ms9gsNU2hrN0+mKurZl2rKjBEdjtPo/0vy33iYPXr76i/
tKcLK9KqVt382Jk8UadQEySKbOGyBs9XnPTPnxt1afS1hKPw7h2oR2LyALZPeCdA
py7NpW64Vj93v0DJm+fRMVCSAqgjSef3bWRnl3g0NnO2XVl+nOc5ws08F4r8vMn9
FDciQ3RWsn1lygHugZCc/iX5DNjX3Zm9NizUwpF3ycgx5GwY9lbkJaQank7/3LWY
INLD0t5EkdQoYWiq5t+/FjI5Dax0WDb+P7yF9GN/HooGy6qZB4erj9bbndNvT0Ke
OwNLMDF+iLR3PbkTT5YalC9r+YYSq7Or6IgQ7O7M9BfzDf2RigmKyAqOikJticFk
lINEjopHp5W9SSJK200UoHhUd0fUw9Qxg2oZOGyYMgu5skF7nt2e5tZJ+dL6TmaN
PIi3E93NxsCkDoyAVl6Lnwh0IOSncK5nfGwUO3xNgxbFjLLuMPVXhogEKAfczvzt
PQkGN8Pei/Moy8S13aOe2dXd5jjxJlD5g2JsyKTujlaRLfaTc/PBgRO0iG2rpb2k
JsFUqBygXuTALDi4bxOK0maTMZc/VHS88MEph7yw3FY6J/o1AD/0yvH9M1BNb+Zn
m7DRfh2pr88Aoo1DyyV2uyc2O3gG87yPDPuBU/7zQ6odflNOeVYRNmsrED18GsEG
nJSvdroaYym+qe1NPe1NFc+vmrePKzP+8E2+tY5b18jOLrOopZQFYQ7AtKC/1Qdw
+KfrF4tCGiGY0VtAwNmorGe8u0scjLPvXA8ASM2zeZBfQzmVFznJ91wXzuhdfGef
11/2ewiSsp81jTmQfSqIfr3paSqvqZTmX1GL31HuXvC6Undqcc4j2XCSN32ArXmu
YhfFerwvmtxzVauVb3Oq1haKeOe9XQPlfEh2M80nAX2Ze+ih/eqJy8ucfi/PaZ/5
GAOI2zViu9t2YdWxiwhRsi9/zsD9Apatsh+8YPdmmZDnCJWCasORw8c9Bk0kq/rG
ZoIcQuX+YctSvNUbGl+q42OOBsJ0Kyr7CX6Tdbx0AWViH7QHprzQ+15OCz1nsjMg
wX670pDpf1a9SFjqZ5AvBZ8sVTggmcPaEmhQZahc2vaezIqdybr/3jyMfWlDGDja
Ap+Rke/ftLchdvG9IqQnqDXPueR/xK/ypsmLF0HOqIm69i01yRSwi9iLRDyXUpFy
SMFajnp9byOuGr7LHRbd3WUNPlI4n3eyCUEUAKHsGaoMsHnuPk3yQxdzic4PMja7
EeOAhYRpS+ADVYjdM+huU8+1DlhLdjg98fTYkt8K8E6g7GjNHlgsBIRAyGkiPGRi
9hWWAsdU/zSH3k9T0SzW3lESPY9vNNbjQDPBKgefdDCr+pt8aJelHYUonB7Lj/5b
TwqRR4t5BY/l2R23+qvt8kALn4zVuYGGZEWe8DxYDCtKlQiykeOKh4dhWRoiZnFv
wPS3+jzUPDCLdqUhvrXiEb+VTKm6gD5ahkuK7UI/1c6O5pjMAZZommdd/qU+bw47
ZLnl+YW2+DUqhiTyfNdYm9GDRC0vOljk/7vWYg4NRrHAFBdvele8vQsaxTEh0IxU
dX6tLDA97K6VflnWQSMVPbYMvtz40mq3TD3YJ5sV21QfRhw+UbTfJZGXY3cOUNCR
Ji8QxeKG5/YgrP5KXH+FyANW8iFa2Iy20SbtbV9M9oexTT8xrefrAIluFjA+Kd17
+gzGRuTSgZrXAxjH8E1Sm0zIEo0i8kaaBQM/coXyu99MoeNKcXUiXmCKuS1qFRVI
d8n2gW3ohP7CyND2UxVjPoGwgoR0m+8ZpN6jxKp/9t7xBpfSHbBoH62cKZzv+CsK
3ujJoLQ7mQERfKI7tZ7DdPAqCm52LdA5cnxvSWw8G6XLdISHDBKAXXUFWSgxz2ZB
KRuKR/8YnOR+NhMzaHNXJDb7AoBwGQdhboveH6CURwPfzp5R5L5cA78cE8x4jldZ
SBdluoTmKvylJ9S1tui4/je5cFIeuFv5ex6p+OI+2nZorA0dqpePyWu1iUGbZ0nX
O9DeJgRJC2ij6K/T4Cfh8lOXlOAqoYrZHtQJRtnsiuX9SRBVyWEyunI4BhudAsHk
WugZ/eHyr73Va6Fw5Qz7EX75HxUwq4SDrrCub1uYs/CexHHHuzVwVvtLf6NCORdr
guVJ7lbZaNuoKMrho/h9mU0MdXdt58PzOnQ+fReY9yAfQgrhdN3Ocal4tijyuc/n
ZCc8urrJgh6lnE3r3OFokVUxxTNj++7MWpOI94scBCDKeKjkCAA0vYucGaXZRDto
HTl7XRRl0HfVGUATvAIcXy7EylvgSqQJPV3ZACcT8xTQ+oZsbEtmqsf8UmsLRUc+
WHaRmfX51c8+pn0DztmnLF0hXtjkoOlMuThxhXtWijUY2AY0UEMgraitX9jMHbP4
mY+sTme6ie95CS1NFNtZKLZhvV4wm4KfVZEnCG8TuhZDci1tlJC+XpAViRZM2/1q
0hril443+oCXnFl2Lva9lsaSebw7b1KN2ueqrI+O5N2sMFDnAR5OKq8Pi/kb02Av
4FBmEw9TvKvaDqqeXkfo4XmsCjAIiFyB9spJNcmx5CYxbYVFSCyeDhOxVuLaG2Kg
vNSra6B71+Xp7Dr9a/nfVtRVuAxELaZjvKZCz8CPPwE0HLnxCsNkKOlcwp0LzupB
ofcBlMxEBYegvglLxqFRoIrH7yQEXa/CIGWfmNYsGgF3NOtzhw9egjztk+55qRaa
2bWgeCVSNYDWRT6KerS4+71NhVaIOgEnzhI7ffdr7iOHijvuh1ixr7kPYrvHPb8Y
zAwf6r5iQNeRPuhR5R7GoLGwqpGzcdG+wmCi4siLlnEgeIcqPG6lukI871F3o6t2
PsGdc/7l/ED9rTxzT9OKMi5czip5mss9AmJTwD5Ka4Z1zzigldwHFTptrCprojcs
DpTfZMechk3w8mYFvqIhYzATRHUtutoT9QSPztT1A7PNi7g2gdPJbtfATVSRO1HO
eiSlyJtUzRoLTrOxSU1q9kxVUymxqyy6xHu7fJzzlE5IHgnMLQQdWVbQEkWT7IhW
ajCUd1YZ3ZePCUnuYcOzix2USNUVJD+WTxw2EAvdT9dBnt5nV9NZSI4uCihZO+iQ
yf5Z+cCHNhpUJIyQryHVeZsFdonfPPlOOxHzcnBq7sI1x1DpvPmzVR1Mnw7gTKRj
MEa/2+oyh/hp6GfvPf17wnkLibwotU93FiYMz8w4PAR+ausakDC0fECx8815APON
Z2XzlfypRYfVhjQHPxMnm+WM25l9SYf1fPZFSYPXbKl0AoWwigPmYlNC6xU7ftjx
WYMdmUFxyJ4ifpIpaoHdq7lnDJiV4XNaYTp6CbtkTgL+wSnyIdE7rGALa9eYmZ+h
l6h8/klWmH3xpjCf5ISAofwAmQjY/jDo3UXAXOWATqAIIfZlWC9isaB3AA+kBg4b
fJcEu1kQf5OEpF7ZH0AgLSl+Vqm5qgNx88HOfkbRB3+EhalKgcwINw/Z86pEV4E+
We/WAtfJLsbqwtevMVYZSxGFPxZOW4A36DxOlk4eIhJuX3XIEJpWRsF+AZbSyUqf
581BeG2EQBf+mgumCXBKKY4sYRjA/zqz1fTlwGvD2+/QAhD69bei9rWSHXSzl8A4
LtwCmOkBoxsq8GExu2BVI1WuUt9ROPwMqf1XyQhViwrZRp+HbvG4A1lst0svYVfC
/wvuJutF3dGgmk717v5WWWTygygGcuq6s5yzkfdwRHsK7qhaDODqdYRfQv8u6jGz
1e2KuHPinMiUaNZGvReb5jmLgvk669+Kbp9y1a/9Wop7zx02+YEu4bxOZwfOVSug
V5B9Pcr6NWr+6FegXVzJlFVdWnpzUMomW8o1whSeE0n5SNd9E+/GKFM0EV+T56yW
GAem+jdQ8HFex503CJ8stOr49CSvzt5umQhd9Z0IieStJbavy2xnxyKppwAAuof9
sh+Aqm8sW+uyt/M7VW46IDtOsibVMAUo4bLp7uAY1vZU1rBRgFqvwjhPX5ngqq9e
RQOUkrKcDsY65sEyNeveDhNmcy4wOeJVjQ7fZAPIIMeQ9C8oUCPgwig/Mh5itmjW
QJPRfKjKwJLt+9zmi/YbJETD9XAXTNsbKphx6wk9bMDykD33jKxjb1gCH+nlJDqt
Juu5i7nLYxx6ddoHrEHIuvr85VZzbAHaFHpvw1otiWZo5hhJYgk93KJiGwzTU5zs
nfqMWQo4I4NlJaXAu9s0I2Bp1vBm0hmjmP52nREQfcUT5z4xPoW1nV2m5an6RZ0E
ZXBMKRd0CBNvafEp+baLddrItQKrMH3+WVP552gxXnuAgTZhEMrDP62wsBWeRmuL
ah7QllyO2H2iVxrsVkvblVJlqKzOenvF2jw8pFCZp/J+ntEnVCqh+CjGq54SQEZT
0ega1PiJjOK4Mv0bUEYMkK8imtTBDRTiZMbiYflLKhN59sR/Fa7d79Poqb42Bdm9
kRgqyqsKfx+14YG6IvenB+yrNqWUOXSqukpLPF49vTQUvyONd6+B5RS7xXNc1IAv
l466pxHuWBVWxD+uEYtBnbpd8L18+Pe1Qp4+/2PbxhL6A2/Jv3jUWAO7JelyoXfe
ShXgi0GnDwYhw2Fu2xwVMYcZMQz7PDZqKJSzWGwlRG2jxP/I4DmlOe/HNO4tCaCI
WNlsbavGkDftrHYDu3y1A8s7k/synBL8/6Fbi+rsDaWQd9nSTOz1SLnISJtkqpWk
b1SIKLA8/fnmu5r7Mlp7K3C5p7oBOzJmv9vRAx2bce09qK66mdTAzvj160uB+Mf2
vp2O4jMEBdhpYnSznrPZbuwejRs6Ld/v2IjXj5c49q1IC4JzXHYDPSxK6Tk2YPIo
u85eTnxTlCeeiowsHJJ/XJJsAyy9ZkvvGPCzrjpPwrf/3JPqw9BjpLxYFNM7zbWY
AMHcY2f5pwJX0l5wHyvTO7CimwlE1zmkd3Uq54k9I1YA0cZ4HLq4gHAQEa0q16Yg
4ysru7xoaUOdPUpLHivM85vILRsgN5Dh4nvulkAmfiHSoscObxAQkcpscAUHHlf6
e9jWDWgHWawVGQ68fb8uxyN0FOvqaBNCXrctm3tR20LAc7Wevb8Dtxfc7l+rTvyQ
L3J9ufyWxbtSec9HMslkZl/LBT5JHyOjNBpWRHa/UYRtspw0JButMmTp+faMBSiC
6MFpAKOMDt6AILtU9GcIbEUFkApMPt/BDRVV/zLYnKYqdJL8VNNYexf3nBmQvJoV
0oA+YpPnrG3hxfkC2vhryJqwxIyom6gCB12uY+i+r85jDNoZmOBw5u2qrw9nVO0s
lPi9/Sw+hg2r1PQADb01S7QmmMcpuJRSE4/u2esXP/WIZjUonEf1g/F/efX613jp
hNoDoYfY3PSgheze+HjfSRQ3mWJIMJjhKAhop3+q42HGg3GT0KqhJWIL9PR8PL57
itleaeD3C2O+q+bYapZoIPvVQe1WCw1xcTrqIsReQjZqs8Yn6VKZC0Ju0l1tz6WG
XjjH31PbbcUtncSbYRWTVDEHhnd1FhohySeC7jeDq2JujAUvo3xPywaKPblMq+eN
OPAZx0NMmocBKvL23iglwJjAdVSyTAw9ACt4lAqPLFhVjLZQyvDweTjboCE589Cm
YUwdE4gMu4ojFpJopqHy9lomiVBkuXFzO7o6fLtlFW5BDabTQHxEHt/FrCuG8hBc
BrSOsPz0dWuz7Hgm5N0M/qaGMYxhYwYX1+AZdezOOYxpO8YVNiuWwkeWTLVbBPni
oynObYMiZ79d4mZmhxdI/qu/1npRC2af8htxJ2hpw2Ir0dmvHKO1KB3RJl8KYAPo
Y5QruCaP9p+1nED/f+YZKZalggwVbw+wQoOyEl4mCnirjM3Hu8XENiAQBHaKF4rK
mDut/bxfFYLLTeL9HgF4sk5ba5/P6StUlGoTR15q0vw2nK1foEO9fnO0pdiDp26/
uL+oW+fn+hkI0DNUaelAftvFu/V6Ai6o+EpQEyo/PJZSCNZYRO+ZY4H7QtpJ5/Xf
pYSa+TVD9uKluGNRhZpAhHdbgLWrZkvCic91bfdTwnOPMv5hpZTu/zZWqfajzhCF
QeU4ENzX0VXIHcvN4di5l2f/kwKah1vQg1V+ZqzOdNAsbTnYIXqyYIAku8bqIeTi
7QZncqHCV5qKXkLQivZUUDwm83bkzzMFVNzIP5q6F7I1cl+JvAZGnm79bfryivSe
DPCMgYTrntCsdH6DnUb3i89suZP+VQzM6NAczuyUaivFW906fhsB8eLw/BVK64Rs
fwoO2ERC7/YfxB0MQBtUb1NBlJ+fd/oZkdl3vEdHT4FSN05Ls8qS+l2SzAklOOv3
bGRH59hGYOYG1IGkM4AlBEMeU+eCcfbvdjSzN5nAK/b8fsKpMNRQRKtcAm8YXCPx
4CHWnNnzeD3dn4wKBpLonDdK4me8wicncJ6mhCAswXreZD5E4GWzNdf1bNazoaIo
aWHuiIc3FaIxK475ynNSYdBG2ueDTNrEFImkcQPe9McC7Z6AUzTcL4tQUC7YzU/D
UNrYm7oOr7ORwsk6iBajClqgtaj4W5dcuN2fdPGqyxaZOwV0skvjgJSEZ6t+OM7r
Kt2tT/2+uXZQsbp8AXKKe1V5CyBereDrfWDZTACohZrd5VHLx3WINMlXK6hZhKK5
J3cAIJpcRr7OuWz1YS+j0jlFRgrjoExvpgcvObuVRk7A5lKgxpMnmmuLGLZLRrvQ
ircV7DAmu/2qpMXWCKExSsFcVjORUS/Od4Z0j8IW5Oww+cvm4QsnvzgRLP1GxIdK
IJFNp4u61KN8Qk3OSgmKjRecdv4hD5tKL2WwGz9hqmekxrMstZVCNvSnpJx7i1ro
/CW87Nj8gJl8uYp+fpMeTkkWupvNkm+sO80fmnu+uqsjgy1F2VVxSBrQa9fAWepC
ZFfF8Yb0i4ig8hZdmOOdxHtyJ7GPE4+EhlFx854JYsOjbAyUoj5VcXfKkC2Nz803
onqQJbUR/j6/nnrWMnIwgjRqG13yEiZESVZj9cHOCeSZ4JW3ENUpH5qIUl3kW9MB
8eRWIAvPhwsbHaGr/15fHWq0jaE9e45e1G3+0Mucyi3vFYSUJokf9NUCqsk9hZmW
MY5AmjKRP9io1M4N15MmmvGC+qaavdAOmyXp5I2oeA9Q8V6leuJ5epVZwPpXEDYR
/gsLmejXPPnM0RALraq/uHghZqMEivHmINmWySjFPY2f/obSnZPFoOoxSCjn7osF
/eJuvQyFzfLsVEDMZoJlKH6OfIor3LQSOpItLcOOp7D1wafpkwk5nXtZvpJ7gJ7y
iSRb6WbgvEri2uyz71GB5F7lkVAjPkGVtMfewjI93SifJYV1Snp6wmUrCftMQCjL
JHmSYXgluHwSsbFrhw2Ics2ipfHRLK326+ppk1O4CpP9CgCnndanf8LdZN9lexG1
625MnxKXVCo51RzrUL4EpIFdmzIpiM+N2lTOFOru2srMySJsl3IbufMykdC0dpBk
iD4CGJq6BGTrvztUWXZZwt6x/rWZUD9NA+ZmtbeTbeBLCPZUjz2/uNWr8VvnJpmA
ONGhaZlyRQgpDQaQB2O2TKMlVJGIlp2Toz/DNkgzQO6NLjWoFsRa02970Skoqn37
c13nSes5rV43qMrZ6omvzsi0x8NVzmaVW/srD9R2QjhJP0s7+bzYTNc1uAfdqRRd
gecDZFjJqiLy5vtrCuPU0Sd2z5+GALDjr3jO4mBQKRn7aXt/Drc/+PS1vwQTMqD4
EaVG9P0tMgs9azywT3P1kanaplAG6HUhLobOgjxvJUqLpFjqUcPj79NL9Gk4kXpC
ajtNPD9meyujPACaGRte3KsFwpyxY1PRGMR5LfTcLKaDBAOO/9z7B/oWqxYfgCnZ
cFofNWSII+koY7x8mtYBfu1y1vTYWq2dSCi6cwOmEO/aCgf/9Djed9c/bTBmbXH6
odg5PsVlbrff83flfTkfzdAORYlG52ZtIdF/Z6JuvUoDM0LAJ6h9aUZCiUaqr1QS
jaTBkLGzTr70UoX+97wRsUx3SDjbDLCZqe/EyneRNqR1h0WuqqLhRfguzQ8MXElv
/aF+G7rNaTwTtf8hvvuv4cTuGXhu9DcmG1OOoMqg4ovsB+Wb131XijEaYXchucV7
3AyOvm5etVhr7/KlCc05WK/mF9RQyGZsd855GApFNO6QdlLO6UY2nzzRIL2smM+K
OI+PTuLch+9AiwQ+77utNAEYT7cqsSNeklqIt1YN34z2zo007qTFRXGQdFYUpohy
PWvO4BKLBkPP35LvVg2z5zjbyStUWfNXNXj+RlrXfWXTc23cVwgOrW2Wb3vKy7VH
/ANCrPzo5rmKQFho1ib/LK+OyqGxq/e1vz0jEhrhvc4BvgRrPdPeyD4GbUqTBdAb
pzEX9u2QtSsfUEgSNoJavosQl+rPDa4YnvSWo7V0qrPfA+Sqp3mbmz4cYMDkOqt/
idyg8NRmmqnvuASIHKZsliPDm6TOtdEfGm2TvJfzHNDunzqDBr08ya66jcHSrkXF
ZhtvlUhWcTQvBKmvmJ/bECsdUNr1JBQD0f7w5KFHj6ioZmflkIIGxP2GR5ysBGP6
jEgHQSVmE8MnLxEMtZeqzWedW/qIYxQqIaCKFs3OZGrr64tMjEZLF/1Api8wpOS4
taDmTMzqMXkSlzNIqz/4bU6E9O9SRPYcy3PfoGkUJ9Tf6kpF0nJeTPsNF3ITGLdN
rfg22zK/V2tJONV3TkMUZDXSuIoQqMqH4RWzwZFg4fD00sAnDQRVgQa/qmDEjYhn
u+vDJKDCt2z22IzhQXMV+isMzhq62yUiBUdLwdgCsiQiRysNcqrBcyIssRrCqU0D
ZI5p1NzdQl/YpbuCZz3aYNvsloCLObd5nnonblRhtQctF5gbd8ioaoZPXiCx0WoS
A1Pgw4f3bs+8wV31jdopfEq0JUjXsUxJqB6ee8DUaaYscOxHDEEMxlH8SP++9+3v
WIbFbXjs4HqSqwsRGUft+UECGl81b3JN756EGy7yC8DEpSKn9v/M/9ej6776R5+y
CPgrgYxq9fDyGaIG+GHZ1N3lQJ5BkbwBam7Qb7yp6NGB1N3HdjSE3spxr0HOzf3p
`protect END_PROTECTED
