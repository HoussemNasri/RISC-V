`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
avsBCjIBSRSEEnM3PakgC1JJh7j6z8ih2iedIFx3ZjULEnt1Y4lZ2fd0FCkZngSC
NxFN8LQdTpyQG9mMSut7P5Brb5yQXsjx7/YF4Qbdc5Yh4hIzkyGhlfOlpwzgrMRs
+YzMeclddhwytQZLQVCdn+QO7MQ5w/lH7Cl7VBbRkHo=
`protect END_PROTECTED
