`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WDVLZ6+4hPNvWbjVKIeQPjeUQjxIXRoR/xGhIWHyb/MrxtWluIrEsv2d7zZvyoqX
ysZzX8Lm5WxqVBx+4zdu1m1H3jakP0VOBko+R91Vt3yDQPC2dOzqifbOrdTme4bu
fGpk5LJtJOZZi8VD5BsQiq2bsV4GEc+T4/Lo1hlEKVyykMqlIosZPJdnpjEZnOwG
`protect END_PROTECTED
