`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bdBRqXMyFxWNgiiSdqiMlvyTsJQ+J/10LQA/A77Rk6g+wR5iTiYBQrxieZkbjzny
H+8TD17dAfOTxBA3TdEjkZn07ltRrhpuWomx3Xa8HiVLdl5i0jKkzqTCTuZ5WgpF
yOyZ6ZXk5HUZPKs+WAZKfSxnaQiSEVsYBxguJmQ9RGXzyC4+1gxVgQRLiveaHkcj
ns6WfK+vknYwUURFc3+/BzfkvKYCHp8uZ2EceAXnL5S8D77jjWRl11rPxdb0N/Da
ptU4Bm0Y6ivVidYrsipVnKME4Pd7qEfEDGh8aaSOTeGci2CAsLE8rmXyBxIKI2ym
oudMSM1smNjKzC2UImwrBU/rT5hsebrWi+SV33n9tZ3uPZQpMIZDTFhPwOI/mOxY
IVYAevFaJZFCDVtGap3Ds7rYRFsKukbvK9e2re9Yo+/FdUNirRIdF68mBWn2owzE
soUtrPddGV0zX//1+5Tlz906WU89FAxeLLx2+48s0lgqah6n6g6DTYqPnTvnQQ7m
gGru2pbd5j08k75BqQPtM+nrnBxa5kbf59EnWt4xvV9UFBi3wQepOFcfXVARD6yQ
TKi+BFG9GSJhYrXBlbty2ZBG5elg6LdjHDVjFE/ndRdrS9CcrOQn6lkQC5UuKh1W
5KCHr11EJczd8qPiRJz3FSnbOdf2ISe6x+as5GsCBcRZLwv1pF7KC42GFiJ8XKG+
RipdR1Wjaj9wdsnPWHD7MHezqXYXpZsRurTzx7WHEWMqcgA0WHGy7CzUg1kMjtZe
MKshvpRsCyLvZ+S+1i5hsePzm14RkwCQ9VQh1YesIQ46Lr2wuadIKhCXgYJUrpKd
hj4TIvU8qGL7fTgzIcT8iYNTsu097LmrA4rPGKNPYU1hVtnVzZN1RrVo0ho3W/tB
Nlf35JKoHNbcegKFqUS3D3siZnrl1XqBd7i6RnbiDpU80OM1sO4Cr7/JfRtfYHm/
C2BkRyuLDa6mhXBR8Kn5oKyaR3tUl32TXFsML2GI6nf0o+k1wwdjPX5/SBupNhyc
3XRxMRr/L7OI+yympHa39SACdW+ubjJeo0TPz6UaIWQxB6czCRhyMM56Yye22WHs
Tk54XOQhACwZZ5khFzgjJ6PPLX39L4UpXSsoYI84B9ZJPT36mfN2kBcFDGRRfiPn
DUYkUT5zsmmuW755SdGKFxPNXx5vqKFJckxlMwoyftZQ7+gYIqWOlB8DdQGS5xEI
DYg/Kh+TqtbJDiGdyCdQEexvSQeLEnrjRbXqnMdHTDhxpufiJ2iKuRy4b8MNowWR
DvgQh7mTFUUENzq+heeMguKZSQeT+Ggaucgq8yePtTk5Z0cb7rz4aCkECKgDgvPo
zGShgI6Bl+tuDeM5urHNKu6crEja1gwUcsEmP5vT9mKKyN5uNpw9gtyaXgTJfMUB
QrUrw5IgAGzsDDCsCVMJY8PWRxSpCgk+iQ/E9g0ftd/GVrJNew2OzCrWOtKxxOOk
UGx9RjXFO5ta64nlM1t8slw1oY/frVrlJ9WnkGpnSKokw4ieS/i6MLbW2FudoS3H
FWcVW/d/EiUrj5AGOPh+6hNarY6UP4SBi8LklvN3hiRuJS2enZd3W5CmAdTNhp+d
cCClq/jOqAcEi0EUbHnZ3YE+4f94litABXtymvrswL8XXiq1WgV4mfnnZnN5r+RU
ULWrX/lJQm5Hf66cl88Dj2jIzdYVjWj9qPmR8JD/M1epl52ZKplrSIVT+nSs4xkG
3KL9zcGE4SRdtYB6bfe0a66kJf8+Vh3I2mHvyKBIoofe/vsGWgRROycveTjHNG8Q
nHoxFojyvy5Qofl3M9OKb3nUea9sZ05KMnyh6X7K+j729vX6Ku6BK/otCCzu19Dr
RHzMmlbkrNOZVt7Xi9MkPz8ukg40M0hW0wr+pIrul1SFF835s4V90FJAYL9P+jtr
Z7FlAT9TwOKVaBPIEJq0aCW3l+8dbdogwfc/pbY9P6G1s+npkb2BPdkngGFOVCP7
CW9LwlmiuM1Qsdq/0kSOnnUOnd9rGvp/+hop+as3kLb3qtrQY/6vhzpqZhvamA/E
A7Ka9PJBT5wouADtEFlVUAfLj1TQsOo7VYe/Df0jFDkBpquOCI4PpT03J9BMtL04
WTpw1eaddrPw7nf+4FPQQQUi3SZ8rXzRwWKc9TCjVB8f97WNdqqC3GOmhsYy6gGT
B7FxLyDJ2fLvyFhTFkIzxW3vDNz3/ayF60b1+7gqd7F4ZcSCHBsXrmdn8G7mWQhT
LLEwIyG1hRurjXNMbDhryndXXSafDqMKCPtEHcJNamYVfC1xxBndTgGVRM045an0
8jqQLHtzBg7lyZ9nLTML/cmoB1cLegkyusMkAckIR/Jl4StcZ2bsA5yKFiBfatj0
CS9X1nFUcTFo7tJFhnl1WNiSqPj+9KVQp56VeKAOV+fUYKFTk5CZjYc6+fIiyzLs
PrSeaqbIhigVOpGjETQqbWHudo6hxQpahNAUGeyvGhLnu3pCGB6JVjmoB7HLNWKs
HazTIhhCv2UPKO0ah/hUTi37PRW+3a6U947Mqw16gMmOgOt478MSwtkpYvOfTwuE
5ZLlDLASqJVo7CtjIGMuf7jgNWpv1+P+1plNzvG/PxtJNzeP07tA53vMmzT2vkVi
KdX9pfV6LASl1sMCdkZpEwf4qPTGMoxEXsrXw9Z3TW+WIEnci7Xg3y+aTI8C/nDy
YovBg+Zem3++0rSLCPv5sMEOMDztdN24rSoiZmB+9e/pQQJN17bGuR3l375lFkIQ
IX+AsjnckdeesZKjBq/cf9VKBsecOqgTjXEcfR0uXOSJiVb65RriMDBBwABV46V2
JQRkPbc+sLkyR3ddNNsXn7TPWZKWYI/yS9lgtBQNn2DAh6VUH3+ScxHLYtIzLSyv
ApfHi6Lc8A1lhrFTJCjtB7kMcVQECfzzZjyxHVU1+JBHhon0d0SE8Mu9Z9LDkTnu
V7Z77QrWIKQhgW6MDzHC/g2GOiq4tH2bf9lE6FfCnbEVxhfNm4TbUYrpuaGfwZTy
G66TyMdVzMo5BuVxUIdba11w5aAUBdUAFj2zSdyuoLbcJxpvYheltA6FZWq3gJVY
BHi3MRTuJMT7I1BUjUFhmVCejZNMdKagP9UscKjOVxc6ud8tP6sW5kTn1juOb+jr
73iophm8D6ZDcZ+sr9h6yX7dr5aCuwE1XJ5phsCiGiWlCBoCNbG8tSIJIAvW5Sqf
1feDoukV2nk8kX4f2sAAZxoZb/QQDyaf87JL1/912VJPc6xQXbrctllYoStozw1N
IjO7mSlwjeXOZa5ERb1DNNBAxAzfFCzl+yi+iRk3eGOrz3nnssv+6mR6hR/D+U4k
RMzaCxDCytLiYXdp9qSpwn9vsMwAFbjtZ+or0fDCQK44y6qqqLaA60LIx7Yg8ycS
QmrKJ3gRPeTZYf/M1zFPsUeQmuF49lMgDg/xR378BleN275CYQj2P1Ei+uMT0W0N
TFqKJEvguwLIRkespJ4DboWriamXaxpduX0os56nXKI+5F7g/uQxH6c4nYUoEnmu
co7UIpvpgO7PzDGdjdnNr2HZpQ97HEiFciOEXe6JYsul+sLvcib3jvYuIOTB1CPx
abkvUFLzCcYXcDt+YIOxlcKLZJXpJpwUWE4ol/LvNgtHgFqsiaPH13wB5eZA+ZyF
VIN/XpXXsvYxpoIMC5/RuG1x++y2FPJi3YxtVe41YkyGQUXHX5dMS9dkqz2HyFEG
Rsbx+m+qw5frYj03oLltOijmNwHHvpwMOP6VTDRanLvbgZgDlowqyAqdcBx30Law
tbLD7yzh6UnSCPFq+0/URUqwUDtrE9j8uVwhomIEXBaDbYJ722nac3biUcsPcWBl
0KIRm4dn/QbTYhX3kwAWLyII3aWbJL17g5WsI3eGmBr9cTh4N8sDO2qAvzb0mE5o
ZbHcYsNmvud56UEiXqo96JyU4u5jbUN7p0KF8FXNr+DBvNjlwIZLgI7QOqZd8cSv
dRDfcKb4IhwIw08N8fofgQ9ZeFoNYxsXXjuvI5qjWTB42qjrN3vpvRJxpRV58wLp
OX6Zw7QJUo0MRgR+wAeNlBZ9sszGcKorD9AS5eVP3OhoWWkiU9wFnv5MfnaY24Ay
P/KHMX3r9KBPHovnrhyC0hAilLb0//Hi5jcAvRQm5kgts71HcUUPSFdbniWKs76T
VYzFtmk2JrOycrrTUwgVV+vFFCokAqmtOTpt1sNlvClUm8Xe1TMz5i2MPORNKgfI
8jYPrwl/xCbTh+d7u5/HKVZ2JGeTT9FLmjXbIkIMs8dtp3T0X7nlDKvc9yUNgjjZ
LJcabQptj/KehoJKCN3l6Nnpg1UVMBE6rpHJ36UCkdSGp2ObwIpToSdnuVHXmWPZ
BSBlJZ9UFr8WgVS9J059rSytUy50FpPgENS8GB4BuHfr68nDQyzWx8W1aeP2RgHj
F1c7hL5WNgeDSb7TV4E4IoSPfLGmcSLhXLEky4OZlyNO9mM16UEuhK4FvS4D7fn3
iySRYi/i62SztJORWhX6HB+wNkyKFtpBtkjDHsp3BYD3QbzRSBl60t3AY3xhyKBw
KFwuBlcePF0TPEzjYKiOYkqAO6rtWGbm1Jk8YR7i1fZa1ONwHNKQKHwvAuvQD5MT
XQuybj7FaD2I/Rzyx6/Q5SD78o6sTGzvNRKkEOgEh00IhMsbyPBBR8BMiMUWSBwO
quVo2HsM/uaeOZHdtS4gD2xTwqHDQ66SzIRjVMHy5ospXpirXJjV7+6c0Tr+7721
28kR1yQYfKrBCLV7tXc0IcJbk9Gbvw6rEpGT6qHoLvt+E+PvSqKUbg/ZDcM6sFfy
7nlp+t2OU99B2ECKqh5tn9nT7Nceg2dNM6MOAOwEC3RWA+2HkLvMlsZV3B9z8ytI
axVPQn/picuFspjMzdIv5Y67bCaCcflG+UIPZ+FRI4Q6GShHilVxIeBGy3DwljDN
7QpLDhYQ11M+IYWCjjS6EI/8YvxzCtLYescJWJiQXLP+ZBGff9oUKsJP97Tz0NuJ
DvxRHD+liJI2f8x78f8blbUu8A6V140dLlwTHwRIRjSZ72yPRFtjqIui+7sdzv7+
w5Kbr1kOceIDZ6PQPtNRNv8RQG+BtcrmpDOxgmS27y+Y5o9I98blMNCuq3JNJ5qS
JW+A/INlT/gDMLh0Rdw0ond2SQyklUDUNkPto0nV3Fr3w+DeFYNnXgHICCivKDT0
p0/PwAK2pIxrfw31qGHlR3Zt0T1tI6tF/ljruKsNsiOX8mnigUIArV9+oWqxUlYL
40nMfRG/e0+AkLXzD9s/YQ==
`protect END_PROTECTED
