`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yirT/0qTODS8sas6BJVbrxkazr1jzvKWb7U1TsnfEHGxdGFq1snJHQX4NYTdjM+r
YYDIiAd5Lb1B+nRa4IB0tQHMFeLG90UssXSBf8XjI/BPkCnpq1Cw42fduVGD0GVl
V8R7Z0dX5q0/G1inkrj0nP0BLIc2sc3PiUB6qzXA7LSeU/eGXQojBkaBlI6CFXX1
u6PvRl7uxomb8kWkYglg5O/nqFDYwcfiK979CQbOAgIAVzNJKDgDA6UcmHAdyE/G
hkTnjR3XqxQIuyQcpC+/HHIlMcEq5yWywtORgF/1oM7DsHa+28Yy1RbMoKjUL4sB
87xWAMTPoz//QhLfPEXCTr+eaS8NDalz2BAdAyont3cy/uQ2NIMAk2ptbJtGnATG
ym8405QvcnyU6u+GY2eeVjblNFwLBIM8ZaARa+bOsDDbE8Qm/IEqVQKNXs+wZ00K
3KcbfTwAvMStpH7sn9+xH4oJmDjh+814/jf+SuFR9FvTqAhBX4Lei2rSYwNsNRkO
2ERNQJ4O7+9AtscDPhK4UILpQJNktdOpC/PPjmPDi1GltQAC+6JEwoHL353nx9Pm
xEC8kyHqnrBwiJWM+GxbdQkW3hiwCS92M08xGSWdMKmXo8twZL8H5kr2/3bZcFFx
vEh4s0claw5D6c+n3OGr70F+YNg9nRxByqYMSTzZHmrMvaSYKd4BpPV9qRQcUEWC
5k9rCTChf/0GHfa8zu7cAw/MBF2j/xYkv4n+FJMDiu7Oh5Eog/Rv0K7qxmdKOj9l
m57YoN+Xom6GpxQ09K01NBDHVN53jHQYmADmWlk4eERpGfIP3BFkvdQ0aNGweVQ/
Ls6TSTFU8gt1hAvZHGuUn2FSyJqgMMc2ifJ+iFiLKXD3Vs93v0JStOPI0K1tM6/D
R098bHW9J29uIIhrYmvuVzKDhtrH1NJqqIUBRP6OnqzxFx+J92rslOP7tu8oRW+C
gxVIpJvTcj7I0b8MVxb/4aqoLAZZK+hk3mdaa7n3ApJk9sf87V/CBi6MzfSEC9F3
SiOfCkP76/mbac8h9Yr6tMM1IoupW3nsovwoL5cJoEVipX4a0/L7CjB5ix9hOPXc
CAQFWKvHVpFGHGtvmVVGMDodLfB1tjmCPtYmQES0ykfCe9WYicY+JHtUfEDifX8f
G8RGZR2yGUesWSBvWK1GUo1FUUyhGU5fi7aDl/rCQNIJLiCDMyhIOtYbZSjludGT
sOMStADxOq90wPVjd9k++htVfPN7k7WOnHGDWsyXs2Fs7Lin+aBBq9+W8/kFYzNH
koX78Y0KH5T0CyG9xd1kgwze7L0wT1lRXfS2wMQ4r8tqREsiUoCjrzWhQZWzHHto
lFjPb/xMes+co8d/nA67AyI2oeO0ZF10FM6eRRqIAxJI5hlWeJZ2+clFs1fDh7wx
QCFRqBPUi/Jg1J3xGKXtRwDBABvlEEUrapO0u7RwEoDJbxW10uJ8/lIjdSL3Wfhb
llZTyKjpIy4BdbVi5Z68Qc2lxDVRmZrNOXYhvz5TwtI=
`protect END_PROTECTED
