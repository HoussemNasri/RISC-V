`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p7/Hnf+cFCZaLzrksHofEbRLJdh6Zd8whnE2gDN4wxs89ILp7avuINioDndKc+RZ
JjDs6LL9UKDjC+V4dYqzT11lgDIrQNhWI6DJVmlM+bQwQFPmRs+ILbsn+T9PL/Sa
alBwz2An/3+uzA9E4FlQx4yLgjxYmGCTeclYSeBJTnfzhHPKVnzbKOfA+cSd4sKZ
OEpfVrS56gsa5Ww+fVicL5TyYMlw3jZIVtSsijU7c2BYwwDpjeboH1YZP1tjKlyY
6YoMR9UYbrBkeYXpYPR38GYHDgHzy/4xPxkssrIlZ2CfK1dOCCqS8Oji1XeyCbgZ
Ss16RL7X4OqmNLF+haJjOE5m/LNebQHNZV2Bip7a+2IieoNYVy7BVI/hCW+/AQUa
1NR8E9FkNVX1cecIJQXodXF46Jy2Mg0NPHDKpNH5iApEEKLynpICw2m3uCGjqxAF
3CJqt5rX94NMOT7xTcgYFAaBH/tScKgk3YK/ba+C2Igf8XXkNGy96SsypAkXUwn9
eSZ4oDyG/kFNaEpCU9PwG2ePibuGpsstwrgsva9oe7/tpDFAqLhTIM/6BxlMEwz+
2wOCLPHqcknxRU7Dz4pAsFBsUlHRjTvNoGHlCG5G25Ghn1fvlHAc1DeSYjiuaM9x
WeZY2KAR7PVfHDy72p/uwsr19eTD26Is3USju5sLi9YxqBC290d/4qsIyCg/2oPH
vOBh4YaxZG194ND/ZomAgeC/v8Xw/0WRnushHRTbVzHX2g9H0q/LWKvPqXMkIiD7
eLMSpSZJ0a3ghEqpE4ZuZ+rNNatBOK2gAVVDRuu57lM+YJ2bsE4C0p7KL5yaOra7
JDXJ7mpB/bKxcejKcFAYfXeCaIeuBDt6+yS76eMB1yAfq4QHIRRvoxkc5FIvb2H1
5brr7nv38RiCtJBS+jq/segSlKINx5//iLUjSQXdY2S3QPF+3LWlcDBB3Z6H7gxR
jlVVQtnqv/SLGTYSPBm+nJ21gSD+uYEzQ8g5BSHuVtdDEh7yn/OS9yCnKTMZqPeR
ln1SePQB2TqSCImoYImDukgxHW2t8307d+rBIYqMF5k87TIYx3HY+hjX6DIAml0r
shlX7BhtGXgSsBYGNg8SbYmdPUE42g3jXsgvXhE++XA9F1HCSPbvvl2mP9anF30w
3VEp1pdZCd+GWp+7r+Hb9VKa1zb0VWjdPkINugUoR7npZV2YL4rXu9bLVWjiZe6k
LVdiPnLf2596nyXYPewr8pH0bi+qzdN0HyzcRY91UHpwjtlvMjVOufAAjK8X/mol
cgxC96cDZStz0MvjnWbrC/pKxfQtXMDR61YgE4Zn0IYOoQuY65IfZohUbUB3brij
nclxiy1YUFchDJtqhfKvT1nzfxXsoszqeIG2HuVb3OVLBy4Xow9ReeUPB6g1RK//
pyXT4vALvFrqof3xX1l/q0glFTSW9rabpmHWlJOBnoo4zHy1xYTtG/0gPQXVFEwu
p+uYy1wuPp8kOUIk/gAJC0Ri4sB1JKi0BLFccYT9eLoz6rJFoAs285R9cXTPaoI1
Jb15/EyhGaDuN12aTjgeIPWk+763QFQYsWDhv0ZKbxd+U1aDoNWRfpsDvV2eLoSt
1uqJlfwqGefZTtybl2I8cCyWw4l3AgE0q1EQtyXM/73FBf0piE0GOrMEHEhxHsGz
RQCqVDgdYLriDfk9JC1pwwwOjg8/VsFg+dAdK9m7FCoOJWMS7oirWz1d3knZm8jK
wpsKU7Bb71MInaBc0F35rtKbotOgzIaOrez/65pa1pcMA0108B7PrKKMrWhNl0/G
yN/ru9ka6skVnxEMq5zXBNxThN55pIm32y3ddPHNtCh6/vbb6gLafbrCkrGF5zOu
DbcMFdQ+mv0hhdMFh/wSWmC/Qy5lYkISt246d+KArE8f8RvjLNkFhGWiN0T3CSuj
Jk7uL696XFs+ESCS+PeEmTYGGFJ0msrE5DcWO+adpq8xJGPgtkLSXJXK+aKPDOCV
yzykwNkJIgkBPOwe3JUhgPFqr62iGq9y2FyWiXFolaUXOPTd1I5KxjyFL0Lu2IOX
hjXMI++ZRE4BG/grWAirc2z/OqnovCO0yDjzsEK6PwAUJNpzGYlGhdZacYkXwKTU
zHT0q1mwbEmo80jiaDaZ4u3jxprYoYp8T9RrYXpytX5A31WjrChXm9JIFlqCjegF
RsWYo66Mn1s2eAAswnmgJN4Q+BFYK/Mmzi3/jDdVd/gI6oY/i7boNQh0NLh5O92q
tM7RDrGvljR0JWsQHy238GKXpgjnY7KbjvttugZytlza2H8sZy5sDLOWJyN5HkT2
H0/vqqs1svJUGFyCEAZpeXBhuHJbuTpczABRJrW38SKdYM3iTBPiFZhBeAF474XE
Semh7jfLuEbrbVEnGYprSkXUrU8j59DP66Gy28OrsTd2WnM5F81J7G3ngC0oFEiI
QWjutYh873iyCC1DhXjGLWUyYcwMtL7cARu2XkKnQZvdZWGEIDkyyx5ZBoK04ro4
+JgT6rVIBBLj4YJSlkpa5FbS1WEHA06S26JKTkHi8ROSuAvtOJII7jbINqdUbgpW
OiWf02U+KNrILyf2OK3l9/WERVFwEMgRAq4HlkmTNyek6DlQg+BLff2m5qS9ujdv
a5HCvfRw7siYM3+JGGyLyAOy5SWpKuEEp4+alf+/NyELW5bfI+bbDWhQ2r7TuodP
a0IWR4rfWCd5hJmb1XyyVaaqQHomJ33lLTSVLE+cCFwaqcl0pztGOjtOKKozbILp
1JYIvwJc/qq4uLvBq3YlsRuyLVojdv3+0TZOLtLX6/h719ke3s7rPP6iWjzHwr2T
kNPJfJfdgsOU4SP7k/EDezTAu2+VPXS+XVUdy83RItshUDxI02c6o+aOUIhHe3lQ
UYsmB2Yq96egutZqLVo/wq751jWUIGd9BkbdHPJ6S2IN+dHZoajrUbYv8GC3510v
ParFKKnrgkyPfYarkHnWM4zVPpOJbEekDlo4S7Qju2szfmvSKe6DsnQxPj2WSRlv
yZ1I+/Kl8zyQc6rcufaECwHjfVz3QrcwtEMPM7tZLuHuNyhyinQUCZGIuIWEJ2Mv
VJYgPfnDTNUpKIYy9rs4rZz2Koe9rTVfmVINk4hx0Qdw8NSUskZZalYIcJNAnr5x
JRWPwfg5Z3cAcBxf9RBgArinXr/dd3tBhkYPVwiN+xd7p2b8AXApPYE36i4pHX6A
qTQtMu4UQYyE2RIIpxuXUq6W5NJXgcRPoZ6/QvQXnY/gjAcMu7YlUpppWyyUrzjA
UEhJP/uLvfzKf1A+Y+Hc6fKSI2JEFCc20ul0udT6Wa7KZnVWHlTd5Ty8YSK2d8mr
lK4SmsN7abAJbWIxX9EikT8KjMldca193ks3WUP0Uv1nY8e/5OTZ2WqygaCtnTW9
yM1Sgo1ck8Bgpy3Vx0Z3eLMxD2zqFF9PPoF1fJH15dLIep75ieJFZ6SAoyLP2407
EsqNOTipofTFcg3XeHBcPxd/QOU+9esoq2sgYr90fm/qp0XFXkdr2it1oJUWhiMS
ejo9gRPI4uFGskRvj+dnZweidtX/9WguEwMfmr737UExQTkJzUmFIdiW3uNcvEMN
B33J0QzOpuqVpgUIzNtVbwI90aRGjiPFat4j/0IANt2ZCjTYX3oB7B4+RyA5w7Rq
xIvNBJRaUE0tRaWuHkCnWR3AJrV1sb36vf1H8L02dKnH3KJxPsokgzRJy4gZZ4js
V4pmozb8DFOeeltyEzVGCBiDXq9ZGhoIN9j6Ur9gzg8RyfW0XdqF7QgXsVbcUSlX
wgo7AV7CuSbXUXxw9LmA0W5T/IdZuWWszSCUWN5JDZHrRHyFFq3E510OGGnSp/6J
z9WP9B8eLKo9pTYODQS+h/EiQmIERT24Re3mEhX3uNODyWVOVjKj8sD77LioX9Li
v3azHiXabvp5VzVD0Y0zsn+9+Lq1kYi4jOKviPcS5+v5hMqhBf6OqejRiPmzRzBO
0o2ikZhYvGMTuSpaGPfsDkFCtVqUVgIa//qV9OBkXjLOBeYlKxkw8ji2d0DJS4O/
j3M/ueJNfDA453MxmKddah9QaGOES4aBAqhKJ2yVdxqRAzKYUkFXXejAJkB2xR2/
/Aue7rqZovX6M/3GLTPqXG4gfR3HePfjc1QmGQHNuKB2ot0baL5MsVfzOvi1ZlZX
dgsROqIClYj103vsB5OL0X0ywGctSQKm+Y/0p6E0C/j8j/gNRFp77iXJx8/cwpnA
E785aPtGvBNbSdju67f8kPV6RqyMSUbyqGS7GnbD99fp9HJFRjZI9JV/eK5Ox4fG
IONWl9NTAh27PQ/zqynY/RWcB8PcO5OMoU6eB7NmEHMQtksL6RcQS+/J2eFppqJg
KjLwDmTsKU1a0bgUAav8B5JPH8YM0LANacIkhGRitKT9r5iwH/LdO19HjWDURa3w
JQRSimApZrHSSQEMM7wT27GLZEYp+/+TlYWM5cYaTnVC9JBMf22GP7ZE5jwsvP/o
qmoUSVhwQsPtJhNPYCk4FpuhLBdVPLJbLBEwj70Ku5kK7szXaIIB5X3gi4voBgQ4
2RUtQJgvL43JffIpi7sx8DCrQibLh+x2XZ8WIPi6GRs1Hg/fi4eu5jr8mxh04fo0
S6RiGyEL40TdgQRt06cIgXpCnsaXUeTGbxgbxJadFWBdzHS0ahurwVrBatoxZUuV
hbWr0k4xKQFQI2UgAHHp3kaw0UC9nFSTJERBLmyZPDyNfs2l7TVirAakSVUSNs3k
X/GRvP3RBJz6BXYAGHbxbB2dvjrr0HpbWBQo/MSWYcrVjO1QxamM9MEpSfyxPJJe
0JnjrAr9WzlP8WQc4DhzKkilx1CLFpnraSpT7kr1Ks3+c69zcog+y7ZNI1qBJI5j
ygqTwwLfm9C6MbLiCC4+l8X9O3T/uwzJIYyXul4Nip9AjBdXSxZ94mwbOdLdTrOP
E3edByPkPf83qVe2Nu+eCm7ICxVLjmrhySohkGrT2rPhJFcr6K7947oTNywdbLey
J4VzowujzcWTyy1kBJhkuv4K5k2cRJcRNyHdHP3ocREbuikxV9menSa8mwax6CXv
e6u3xCK3l0VduORJlPFPrrRRvubeLylhmcCbFz6f3Z8aAUfYd4Hg8m9l+AbdhHW2
tMUJGYaK95qv9ch+y+MoKUCl8rr2DAZJSv2/2jGjG3REbCzZXwR/LxhY0p/jsET3
Y/zoFsxAD0nHumfkAzC9CVBq73FgAEvhnlSekRGtGmQWimyKNEBDx6nwdAeporDv
xOMiMBmN93NFWSgdyTZWlJOnFvIxf9XwzmnUUoVc2HtZYizU1gzeeu2G8Sjsezsh
tiKtVQQJm/Xs+cBQQRTd+q49wrRRoeZUziK7Rmv4YPG2ER5H8YuoTeAhzkjE/t7q
5BPHFZd4a4Zy6yAso1MgjD9zAqiLZdiBP3dW6JHXdRtTzfjSWcDgdVanHaM1ysVs
tcW1mQblV+uhBR1Up4v4+swyHK2/82QtooQhAb82D+KVma6tvztlyzNkKs8oOryc
kbygZ5LnVY4/3aiT+Xmu64vBm2zUIOxjT2NMyaIJzrp6sZonYKg1vas7ZQ0N0nmi
BIN6N4iFcrvPE+lhI4SUbkJaM7BK3Rm2oshpvYJHIn78DEwbFDnguDS9Zd4NrNas
UpO8uLPP25iFEmIHc4ePuRCJ3u73h0X8La7cmPHZMXbXgKeLTLp21Sz+5mjRZxF1
b0lRiB7AwKBFiDGsK9LC+BAQdWgFoi6u2VcU2A3j6l0N8mJ3EEnNa3+rIoZJpvgb
55GZQOikH462/WuXcGqf2neFxtqR/lAuUuHCzDmov0cMl/8KwvF1pwi23sHjjseE
LwrBR/sFAo883CZM5BzvurA2o9VOvRarGJJ8d29MwRKZG12uNLnI5dNB3zOdpgy2
a/vPqQNqFyd1DpoQ/jZEV7mIiNv8D18zDsD2VHOslM8XU/ykRhVV7Sm4l68fky1k
GtEEZAtsu8yyv2wxTqh0BnazyFuUfMXlOSxIDzCM4Dr/PSNABc5LkKx8oNwVQpEG
vxf9TdjNHBm42gYQTWgSyDwPErR9IFh0Fr5YfY8my2EwRzFG1i1o4SQjHRGnlIS1
LevIEXDYk4ekdqwZhWxSoQbKqVFEXixYNs5xwjrA9u6gvA/eum4jd5j6RBgfxJ/O
XoT9tN5I9VDa0iCi4mu7uyqHoGS974WXyXQOsxROzAxBZCgfqksV0mE9DXTJCoaK
9jUUJiJrInPKhUJCCoZINPuUgAaPz1AfFDBGt5GXyzilE9HuX3W3B8pzKkuHZKFS
S9q7dkS3DZXdP5ztsT3OMLgDHrqv4UIfdQbmAoH2JC1K0PRUiw+NvYIq4uW0Gg+v
MFiWc6SQA9ulEgmxrJpW5KOFsQeDY3qFlm6stwDyxMcBXvftQysXLMTmseDtJ9g2
jTgog+YiL+RAvCRqqOS2DZzHhhGGl8Q/dr//ZlsydsUv3IYxTfTy5bf89XKnZSF1
lrgDf21tYZ0Gr3RRX1lG1UNjgK5UYflh0II+Tv8ASnwhsrnu9/YIewF/DTafH1XM
i2Nmha60vY5Py4+lbJHj/wEvJNSbdU1UDKgb/0cwez1nt9slJuoRt/2AdOqNmo4U
qX2jrZtwyh6bX0pb/HOKCQkN3EpK/M8VHe+/FwSEx2/DPAX5lVs6a36TPDSyyMil
wqT4s55M4Ic2/lH2ocCv2GjV9f+XhrXLleG231SrWVNf6rWMU6xE8SPHUP81xLxG
nA8qIma9M7q/B1kRYfAgUIEDUCj+Zmj9OJLG5YtU/+9yjBJM41ZTXQ9gKssKt7pr
un+56ok7bna0s4IclDokztGFwiFdSRL7/rHeYfWzSbDawt4JJHyC5LsteXPJ6UU+
pWzcYfN7NTNXjT4kor5WcZXbnUt6tCcY3qzkmQmmiwQvd6ig9IVmn6Dqa05M+si1
C805csZdFfc/riCtW8m9O5s3yvHX3RTmZxPOnxns/VmpHxI60IWa40y43u/CEN9a
raXWqcgemVuxObsc9mF3oqIVIX2b81cE/KPRU8XIFxjmLuDi/Fku7JTbr3vfo3Wh
XuxQWr0n/r3b0wrDaNUe6/H0CItE78WmndyPxMJ+g4m807ndJzBT/R7vW1AhIw/a
poPE49b8wWhCRIGqNMR9U705HqEXbgSloIv4Wkmik6VNO3XrPlLa3fZUra1LNqha
fSDoye2jssH0vLk+tNPn59lXGIx8z4Z6nVO2axw/gJKVusm59ez52Bq2r0pvfsTE
FWHasF+/MtkClvVgn14xXmcr+xq2DxzTH4ze3o3UiVezQgKwTZSdgIVMKRUu2GsK
Q970vO4O/ugRIOFug+jNSi7kzofstiTAluzqRitWoZBNHqjpWqPO6d7vwVS8SaJs
auS2VlN/OAVn8eD5jG3JF76z031QAlZORkVB+UQBPgSAMiRA0weKN6/tn69Z1N9r
dB3WYiOcZqFpoQx3zq3ov5gg/rS2hPjixQ5bcu7RiU7xdvCzEkPhyYzNkUCkqY+5
u3YoinFxW6DH6PkfgVzyWXVOihhBqgrTLkgbLmFUya1AQa75n24FaomSei5tv5zO
Wo4uyVjU+0lE045kbO+Z9cZcQFBT/EdszfMwDbneYFW15qwKnCo8MHqL43vpzfHK
K8lEKaElZHOxVNbxpFxr5HixDA0TSCpC8beo8Ru3bGgDLjyOQWd5WjwXG8w6ulzq
Ci5sgjFQKlSAvBRe3gSJ32h0C1P4KWJgm5kxDOztpmJP9ICw1YhxFBTiMjF1WI2X
9jguLgr9mxVrC/C09SU28EiEdR/ldwDkHclwIHX/XqrolRjeyq9xErojNfhorSLg
2yAE2UqKhD270VL5JUXd+nQNC/WHhO+nkzNz2Dlp4aH6v4YKHVuzotaguxZ8l9ds
DtVf6mcD5XmxMhuCIM9VJgGlHrXAI1yFrDtYyAfjEPQz0Yy8x5qA3AABlBmZ5u8d
/BSGSjY5RQwKF2h3sn4eILo8RjjEmCH0W5RbV4FoVUMdFoHuVHlvxkzhwBaXJRcF
32Nh2rPSQTvN0wf/xlHgQybTH6143p+02SwVZzwfdaGUuUB81dNDC100O7vOq6Sc
1lJqLNT5Q7RysbqL6DrAmoqUr46Azj7DQ34jc9f99KA+WopYmQ5VsZrttqBpcwSw
hrj+yyLlAjbchD6DOf3nQ4Xi/5NdKRjlNrBspuPWTBYX/AFKenVLGsxDx/M+cPV1
/5xXq85no/rrHCLZ1l2ShHRP4ZGPXLYT77M7L0Cot/umKLv7u5+7Rcx1m5Ihaf6P
6tv7HL2BZ7fgTlr90mqMEhwZO6KWlpugceUrfJWzVUOO+vh0IUDS7AqJFyqT+1LQ
ZJkL7jHY7DmGX5e+kQU4AHHXCSgR77ypQxVo2rkzuC13WgI5LP68gjTHqgYAGgdu
/HASDXaUCGaYGssugm2ZIJDXCWhI40pumEUKQZzNmTPJ7nL1aDvOrGYTL3sSjPas
S+uQ/zGA+Et0tixNwhmPopERJfSNdOoLzguSWOs4jwvD6Dz+zWz0KAUzuEhL5Agz
V3GEC9/kVqahlYPzzwIX70v+H/TNTieFbj4EeX2ZFM7p6h7RJF1Ol/aF/hVnu4Ca
Cgh3u4694Azcq6RjvOlaghe7f4DPR4QNTg/66BH5GyFx8xNdGYU96jVJ4asX8t55
kcTfkoihNR3XiO74W3l8A8zIccPZK0KTNb2RMi56ZonwcX5yGvLl3zokgfBduVFR
3m6HQ/VUetjAPit+rsPTdehEHhgl1jY/diohfx4N65cgjstLMSc3DIptjEfbTnUf
0kwy6n9Z9J0/tMRyB7VnEP1PiUsWsW9mhbMa5aZ9GYovudegn2d4AFwi0AT+sFbL
lm8y+kJatfyJp9QPVE+WuqiDJSuDPREFz4MiL3LtTgWZlviOwJXn5j9gmqDBArB0
M+jEoab0I/dW+KXTx0X/3Sibr+nwgOio+Y96UZmbxADJ7vOgkhif+Htlc6N5GJm3
9L/YA5usyu4UyoJCsO/J7AeVXkV4OrgYGYqaCAeECTvAJfm1gLawZOOgx5+PMn/X
qvQ23FAPZXy+O+yYrVw0a4O6UR7kIIiMxwljAQ2iuNigkuGQ42Nt6SbHAfYvAys1
Gx1o8wa8/ahU8L5sOfULJgLOLOmeJhzakQVigZSZf9+aeCk6V/RTzNK8GfOTZZHG
MCoTqUx7Kpm9xufjT0gYrYrxIBHa94bb8Ywt9pGk0kSzedi2lUmb1JuMFdMQcKI5
NA6qyrOK20z6NxyqZfqO6myvwC3Zi8JskJbWlO+r3fNk03ZzKMvZK2sXDDQCKTvD
lkWka3HFJtIAIrKfv2Q1O8jA3DCSZMbtwhi894FMS+Sv9YwQcuuQK0oxMpY3v4Yg
0BT4VxUTwqMSsY2fJ3+oR2OCGETxbOb8Zl7MfunbVi2E/O7NAc2Z7QKfX7wzZhNP
MtYYx25wogFm1LS9zMC+qpoZM7iMtCTDPj8Gc4Yt9o3/WRqj1Ki3cro4/ORxDx54
Ji7H89GcE6H3OHgxzKb0/m5H5hxRTGtfy8XK84DicLhSc2zHNgNKuhHuHa54i7BR
hYfJiwe8wH6DB4QM9GGtpgpftSA723roTwAYIq0jTtgRfwFo4hbt9yL9ThSfF6rY
hTw+/AJLN4w2PdGtC04RhjS2VStFEENBoVdVLA3vWw1AeXKdOS41KeHfJcg5KmUd
zyxkqqwOJo9k6MwN7M9ygHSeWytXxa/Aufh8VrnlsneyhPGSL4SK5o9tNCY34OMs
5BPDFQ9cWTD4wtkGBnfzrhX9GBbg4SS/ndEjzWIUKSM7HyLCptGexnif8z6VtrsK
p0q5ZEO0ysLp9c+dUn9NhN+2Vo45vUnlBwSAkdwCTaKDZgb90BZdBMXay1ycUYr5
7wsDsZDVjMJwJobR6boZpJwFV+PD3w2XnMvmA1TnnmZcGtV1g6iGqAaEm1YA+ENd
vNeF32AGVQUO7HymeZSMogqCeIVPIQbldnDHZjtiZWZn+d3Y1JnqhfRDp59kGNqE
Nd28iN7z9Y7iAKLTZAo7T/O7gQcv6uNS5BdtxWnP5uodzNLUumxcU66SgLrxFx6d
LnurWTe65Fwq6r3AhKsBXHlTh/rkbf5cE32IwNl2SGswaQ0MSjeXgX0yNEmN1JCJ
SiEMgm1FXfuzGyF/nN1Gkrt+3AkvCXx5+GTbSMus/RuW1Vr/PgJ1j9x/xvR3sL2U
MVJSxUrRa1EZrsav/sq0QQqCM1oH1bCL2mgEnHPj8gRHEhuqzVs3avNFytqFHxfh
QW6u78SRy7T3b7gt1OGeKyMokQ3nOeC2n5INAqhzPLwMZ7+q8VG9IUtpydrDrxB1
Ll5qLe3UvyeRFed7pj+v+xjCZcvsfGU82Iy6te503vKMoCpXtkS1nCfonl5HpqXp
kqcYK9xUZ8N2VyuQyflomnCiSlcsdxAZDwSkeWHNXM82L0PhZrRjE/TYodjd0zeJ
F4XWJLaA0GFcHJm704BqEujGaySCXXSMRjFFX36Ir7aLLp9L4H/oo8AY56TJl6BS
gsmlkycEAxjhQCmwuGJbc/RntLuMezUiK+OTxH5Jz2I873vPKW/N4L/h1pyfN/Wp
/3jE+zZOvXqU5u9zqLAuMGGkdRLeTcoGJQlbizsDLL8YqjYPgsIelfQz+at4Sy+D
BS4ArlIOoWBIliy7QD7bc3iaod/HIjk522hzNmSYkGaak8SADmSuHjuLERhJ3Jwy
LGaC51PQbJvm8lhjvqMGsKzksFwQeFonBiPxi5nsCkDd1rogZgyKE+osSS5xnl25
07KQFoz6PkWs3D25csdRvhgHAFkzuGMnPTzqufxkn0YpNXZ/wKnoIBQ5CpDbBtSI
ClsvfBJZ1FHL5V280R/E7ByeNs8RtBm/dfLxQlR1fmI=
`protect END_PROTECTED
