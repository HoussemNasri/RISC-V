`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
miT41LNzcLf4RYlEhhemHiDCH+v32w1qBCO6RtgloAfYdqdg8/s15lKVbAyTsnxi
Qx3UK5RwPVVcQZZ4B9DtD13U802gK0P1kdzbCVr5sbD7l5vcSWgRJzfmPP6QnhMy
fWtK0plk7V3cwVtiAD6HutFX3kxtsTSRtF8fMzq3/tfqQFjVi9J9g2U7g6MaZoFE
8zJs6Jkv5PS3jnjVFi+aaeHYRf3sZWX8s2b9Iiy6DQ2D25pbjda41w0urseEDO5f
o7+Ye9BsiRBOyrKXDRWedYhG9kL1vOUPozwSdkXbhw9g6qudhAYzGuoOiyMEExy+
Ohg2qbpCRV0lapEOvHUgFNLMoCCS+zgRV85zfckiyRHxfUd1DASoGvOl5Vo+q99O
MRptieIbTzKlapAh1iMAGaZt09TIWohFrsGDy9OCvUom8KLCYp5l422vBTR2+Cv/
OV/ATIl3sjyu2Yl9iXW5rb+GiO8HReXTVec1/xGTpoSHdHNmKPSOjtaFFiCCt1cp
UfdCQQ+mBCqNKomWc/zIMPMAhzi0AMDRJFs8b4AhklupClQI0juB5f/ASGOnhaEN
GY1SUchA7WBpt8ybYSmGbeX4SGYx0ydF1IwnDIyNne2xvoZJuSQRWwsfeor8rfcp
0iXMBozeBnbCWBjtkQwk/N4gDMv+XYt0m3tH8hTBHKCNODmfnDn1lTJeO3HNdaH1
NYkIwKqKJzvsmv3nybgvtSSXgB0tZbkWIsVgoezavlTVqYvGHt3GhPTxjcLzXzWo
Wog2zqNlxIrGlCVM5JcAF1DCU5xOCJEFVR16yAKltWnECndTUs1yVLGcFMyZxIyg
kVNt8wQqDlp30v5GgLz2X6Z9nW4ZtUDncISSDDpD7RUXlVKPrQ5h6Ydub7+j4vav
iKsxRdIoJXQKPuTnsIM9i/up3VS4e/PXkaYw0iVcP8+nPb9iyvsTvo+eBWLyOIrU
FcUG7k6qvPmBN4OXO/UbRbrFkSECpwAxVtHbMa/kngivSW20To4NwV04LiPg33u7
dZIRVuC8ux2gORPK8yzfRbSV8U7PaWnUAecs6eM9PK7HKM2vnBcTnbMq/L6Vdwwe
dnL8e+rq8rZHvnZY5SAlwwM0GUiw75rkbP45Beljc4/QxhqdtrUOUGWa6BN0WXgn
ltDu4q6TfEbtEqn1NzC0f/Hsi2zE4CAKGCD3ObPzIxTloQoundO01G0WGENPx8tj
RSyHwyWG/m120RXpEGZuV1VjiTMBOCgCCd2tmTQnpriJPrOgVXG+KKXqXzPyp3Gr
hD+VJyZz7z7hJfc0q4ywgcMbJ/m/Vq7NqzIm8sO8YmJ30eHNvHuUShGbxX47kbeD
Gbf0+B1LZRoDQW611BjOkIxr+U6MkHmG2IgcIbDWcc9cIbNiXorkbNVYkQFvfLLi
w+fMItgir9zzkmtLEruArPGQmXV6/pcaGKQVI+m70dkj8o1p7+Jgw3A/8dlsUL1J
sD3CgDJ5GS5TR5jX9HgfYbPBNBWlWvsf8kiKQ0EW2WfU7R1lqe49JmpwMoBLV1Fu
EkYHPbsQHYG3WMYJ3RJSUq9PGQxTajsB7lLGgr17Wmr8E3mPw1bJCiWxTMnP6Uo3
WMpnfOeNNqM5fFfDZB8gHy/IGXZTrapwCrrQal1Nj0YhN9WHVG3rXQQJ5Ql711qT
DxA0RH7mpFROJ1NWp4FUIIBar3yLMauPumNRegugnY/+WfiKx3vuNj9O3uZozua+
vISFKgTGpmgPjpagU0MQlqhzcK7IYFWTdwZCelS0vHGf/mMrxUVTyN8zIL32y8ec
GeHjtT03wAeBqpwghV82FTL/b99p9bk5dNt1b7JsNdktj5tl9gecgC/NBT6OdI6g
MBnen4UpwZyn/lkBB618UHG9OwesmcpT74Wa+iaG7mn27Ne3HRa/sunUFEeAIC0P
6DMuqwbFNT4qdVKwaV+e4Q+wRBGygY7NZqrVtsl3Lq6XNzybbBKESjkRSo6DrHit
Rpl2I1IqLS/kMCGVdt/NuTnmkr3Zag6CvhhdKxx68eII0YyQ7wtZCieZoltLUCos
hvzKWhNJIO6z7MvnZ1oVBIbE51luTBwnBzMBw4lMNvdWvc+2GUP+J3sWV4BXr/O5
ZN7kXxahyg3/aIXch+A+NHvcHfVFs/SzrtDmIHoHxF5ORgQSt3yevwUjWQ9U/cJ0
4d8AoWKVUhtS1IC3cHSYB6MU+kqvDJVEGDeW2aTqdhzrhLa7HD+l2LU7EoXcWiJX
PaqwZyLOY0OimdAZ03N/uTpCJ/bQjTgAai4YdGaikJowWPyJXxVBEKRx5vtQmZuq
A9DXJDp5bQ6r3kZwDZ+Wct9/WjybLql2W0crbrHaFQh0/Whugl4cKhTHz35qh5Bh
`protect END_PROTECTED
