`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yI1QgIWiYz+pQ+mY6rb0GffRnjfdEwA5mhJLONwr3KbLuhfPKMhF1IqrsW8McAIC
wFPXOu4hKaPFpNam60boLJewd4sDnq0EHrXZkSE/KebNaM+cGDFsGjXeLosMYrNw
56rPsr7bB3wdLHFg35EuEzwtAgg+pzlv/mAwQxNuMQTy4CYR4wuQmwfVAqdu7Vqj
AOWmLbWKZzr2V706mARCHuGyG8ffRjeYRGIUZFyna0joEq81CcKNjrs3WjJQYP8Q
tQelSiInctlFfdZZVZvR3Qs2sSPNshkv0Ll1+KQQoVoSyPx4mvtnQXgJSnYK7mC3
vllJu+9wM/amBVdY2sNZ4EAInllUMxlABSnU/FYRoQemcUWziOugUqIoNcxPi6gh
w9eMYJvBdyJZqhS8eS1XlNZNJ0p5Ts2GtYp7HFSuHFZ2rd5DfHv55Jz33gYSBe74
1aIztTRn5w8xx+jVyAThp8n+lfahhduaQaZ/6q843yVkG+GrdvAbrTzTBmw37U6d
B66HyWDiDVUhZYV36VUPFoJPJp0dknH3uQnhuaA8L6zzwnr/YAbt1SbvpuIdB/b6
C3RHefpgBNWyalyllTjbj64JFY/DDChiV4GZ/GJNSMDNccsWWqLbbf13F8nYFm6v
aqp6mFJoVkoYQKQZZeFh7NhhcUN1PIQj20RdxuKf7FXtXh/ZaGJOW01yzCPGKWzu
TNijFLOC+pi3R3nw7OZ2/Q4O1aGx7YtK/d8qpBWVtXKfMeg0S1d/LGrWiqrMKzFh
L7xJIwLVGlcKBy42u55G/0ni5dLdMEzElzxsvM+41yDbBNDMCyfTfMTRt3+aqdme
hg+lfSIVA01HjW3zm8+g5D5y06CcAdLRNc2Lh06Kt8SZW7I6djeD01BOmcULdMOr
+GB5otqjq9YZg/3Z33fxRplJBeUn7CHxGzq5hAV6frDxoqgBBrYxAyvQj1SsVrJL
qvXTWECg65jr4+F8O8NkCHJxIjake9oiva3KA/ikWRZY9EmooqNSNUXvN4w13hg9
mwuLvHcopWYQqjNuHSieZJ5rCIakmCIwDw87RPj7VmoUn6c+5fxMX/3K+gmpVwkb
7MWWKO9ycHzKVWYtCIz1hVluZ0lyc9RUbZS9msuG4u6zzV30us3hVWOq8l8o/4P4
fsAXH0NCoZsN6NPTZWMf/z1QLUsWri+4Suka86AYsugO537vVVTYTFiFmL9lmBFd
BWMuAD+FdIBPy0QVEF73WnrOc8dTu/+8KbJCMfDXBtpgef7Znyh+CN3mz52uaIv1
HVyFhqjybDHHHSmUT9CxxxWkzzahhKIQKPfSeZpOnrMixBITaCe5bgLzebnmTmM9
oWm6E28ftcePgLax1SoLmtlEFm+nISU+Vv6odKdezb/MHPfeHM+o9NMSVOusaUfj
Ye1HTqVfEHczxd9+aU/zmP+pj16hdweNUtRZsI6MFmv/Zo4LuuaWNK4SByjhPHBj
6Sx8dx6IyLFM1d0mWtExveMqvOryRcr4Vz9p5NvNS0HmlWHau3itu5qAQvgmaK5y
mFT/kG96udBaTPx3sWqkiBQxdPSpI11CHCgq8Arl1ga3KjjhA/vQyY743x3FyPQZ
WLpkjRsG84HGVcccpIIHKDBMYvmrdbe13M1PoMng4f5wFIXpmRZWkyiA5CegC3hz
QB7/ULWTScd3oc9FlF1CmyL+NQE3UdKJ9djcHfiA1CrMzo+5HjqKNV0ddErgm1Ll
jtjqe8XTeJ4/MeOUDjRLX8FrzqNFUUT3XHo2Dvvrr6VWE3acMX4E1djnczWl+HsI
rjxjOSpOIf+qb0NnKGstqoCcSWFEewPQFsPwF6aRHoNzqNdF4ulPL8GKsZuaNUp+
1nPXGoGDXmP8WVV7wbufhAs+y7MVHQUy7IVbanUdMDhi0awenW82JsAOH1xrsbsU
UTBi8F7YWixIJpo0g1RAlLkaOQDDhUqKaTy1sLExWD0IO9mQlQnh8NoVgWWKOwea
QT8OZOKW8VnIMgan+g5pPbGCLcrcjgSlIeX2I6OLXPRlX0MYPGTNsyH6pWKeL7sv
neU9FOc7Ar7nbEFzKVf2jyzJlZ0CYcn1ql4fmx07AZFlDDcxdnf1XL0xVwFLno/Y
nd4/DXwCvek/mUBDljVAsNYdOEUaL6fEksEPrwu2dWoUHZj3hMqfoN8GuFLiitec
0RT8dIZZcjDsXR9LQ3ACsJmDU6y4POlCUK0Qo2pF8wXk+bu2cPBmrmur+nuY5N5v
/bqAw5iHDN+TnRU5PHcmw0RwSjf0T1FWXSH6wOrVT2e8dhW6i85hQZG3jYS7rqwm
sRzDo2M/64EfZVE9WWpBKXmD6LsyX/gxjdFqNloywsu8ozi1WhUUmiimR8IRTyvS
rOby9wIPvzq7yYmq6dyjgyINj8sLxJUvCK6mCxhGmrCmcY6O7+cwc0M54VH2DP41
86hZpRlopoKjjn7AcWKmU2rXYYPAC0X5C/1nU+Fq1L/rrnp/b7M8nS3Npv+K7nJr
JEgI2c+LM7trlVY4z5suCatdjhtf/78NpcO9YguoKvRXFenEDnxnDcclu26YrULG
RkzErV6yizjUmQHBGJDJhP6GPMJQtlxP3f+FJIlj3dvhwW0sJwxUcS2MeFR+7VxO
sTRTwF5+RWt0yMYDS/pKt4hYLaB7wQdajvks4rPtUdehF9NT27mB4Yf7fTqhfSXH
5MWWD7xwpGnpdtW5jGIlqiRdR1KOUeqxW+TJcb/3eVweTtivH09iXpSkI7Ug0UIk
BZYfnhiid6Ik3A+Y3qaEmUXc5c8SQoj7RG8ngj2J0Ii0VTeq84rF9vpni0iDEtgo
f7xxeLZqZRBYoH6901VnOIw0rPjjj8xE+M3HxfCaDbZZotZyLAAN5ftgen/YnHhb
k3oPgV/n7n1rvzATwD+hrQKlI2rgFpBV9uYqo5CBTuNAHDvGcrf7trvpCsqTQZY8
isqtodS/dugGE4RB0L1esBqvtM6AiVjBlyTjuqa4/PHr39XtRcxd1u9GL2Pe7oID
3B3lsAPKYvfqYhHJzRwsSn+EgrZPHSXFVyyxHzxFGhIKg18Ux0ikewWAM9hAAJgc
RGAkfH/PP+JwhRNUT/PhiRmd80jJr9SbqxYvSIsbsD8OdSAwYZqiYFlnqZ+1iSKm
XxBEYbVTkHv5It1NoAkE66ZEbCR/33+Aych2aVTtdQBgYYbpGk7zm6uspS2jJJpu
B9zEe/k02ddnrN/rgJvVfCOq9YSMtSBHK25Fy8krb8zU1oNfP1+E4ugVvVS9fUvl
qQTMtZ/bDNVzV+4UbbB7uH5aYmK5Oxd90kvTvwRNeLxmj+uCO7E1U8OXSaW9SFuR
Y6q0misM2GsE0pSMC48wyGlufvU8SZGidJf9gy15rEbETiKFfEJXplq7WHV9iqM+
2fy1xjP8H+VUiKX9dsUQ6Wep+e/3wLrb9QnpgRX/difSUZzmTeWd0k9rIvjSmjGp
oHhAhSRvLRWKHOhXCquDIxOHtpVMLpOyy5eog7wm+h/luyziJT3HozNjoEAE8fkL
YOMwzbhJfqqPwLcwAAT3ab8XQvvSxq4bg5Ex/kSy2+YpqQ4KWcB+YPU1WSDzyu7R
sb0qlhhd2mogO+azvKWwha29tyOIspV6MFwXn6rypb/q1kXEW7JEhc+ipaKmluv8
hX1kZx1R9lHid7UQM7jrY2N0eePJmCoSNjWDpQqwRg3dcFcrZKY1Qo/4Sl4MACJ4
CuanscQffsWK8nxHpme65ojrJV8CvlX6tRR6kaTfaI6u1fyNdCylvLNgUAtG2ot3
iR8gneCG0wgMnOqJHM8kZ1CmnJrVYjSa0hWfAy/FVvZXxjNQIElwz0OMnUGckV/E
KXQmb+Flb40iF7CO2bMlGOIiJyD2JmOfUiOuLHDNrAhJcxQpvMqjhLsOrE71WG4W
Wxjc6sbIMX2711Nn7Pi7D9Q2H72ZZW4vJm74v0GoSibT2QX/YQRNJkgfeq3g/FA7
8AybcgXvcnjP9dGC0oAQElrjpWeYCXn0zr3xThSwcKZ4CxIaaFXuedwOAgGfy+Vy
jPq0zD2UMwZv/+pQHyWozjtw7Wf9FJDrJ2UNn/XUI4a5djT7eSkhie7bHjST/IBw
IPGmGMVsaJQhS6DOn9B3sLnKJf0CJ7xHRudOeQmwAYUdRjPQ6r0oic/BF6iEIe8X
2f4zsNedJZoKMkbFemM6y7tvWh3pxiDN/WRx3KhIbJoGra5s75z6swN5mR3gc+gr
zCSLX2xSP01UBa1YIAS698ILfqe+uLJ5lMzJJJMLo95E1IC4eOKxZMW09MLswvfe
j+osFXzwk00J/ucVTLcxcJ3zHcOkEyD1dMG/H+LekqbkUOpsvY1eiGFcCl+ygSlg
ZvVV0s4sAZkoLuzxWMjpNQRNC653Gl0EaffTdNwCAftUTqJjN6YpmoLDCirG4O/3
zDUyxjwnmVl/AHXrLvtPG+6Xd1c1jGSYRk4jd/qYkHgxmmQsLnor1icfsqP5iaLb
Q6W4iMh+rxBsxmjBo6JoD2FzoMcqHFmILJ9Fj+uWQXZx6qGh25KdX22xB9DhbUdj
sYMm0WOBbAUyxfNijjMTk0piGQ2WkUn9RRgfHtHC8u1xf2JjYUfmHjmtOmNhLDTK
8Sz8OU5mem+Sihf6RGTmNo2QJRPQODBZUNiQEUamTtaR+9NxRV+FXzVh0aiaH8cI
I4woxbfWoj88ou/aPchaQPoFLhLacVF/ePQVWygYu+FH1zqDh48p5Z1F/yPegZPm
3AcskaDeG6beXsNYZCG0C/z2wsI2D2QszcDGE8NNdWTQYSwAegngoX7qWZ7T1Edf
ZmivOAIJye6X50N9wS3M0qe/yiQI/0tRksNjaIDvNxF864LQ9EqrJgPfq0cXqSuE
kBVUu1EkHVEL0tRTV2M/qZ3u64bQaJOehvssuHSHK74NU5Smq7WPSUKHgW61sIal
TW3ypFKJh6JvFDXtSXh8dk3sJ5tNOnXsuUw+/bFta9YbwTy9g3NKQRHSaGmtjJC3
iTstkoNjNp2q8Jn+uIC3KU7GMqYkkb8VwI1sPw8P/yVeekWuqKM9i9lXP7Qr9hr5
l7iL4z/PnghZXXeexLji+91dCK109ShrMGOiDpkzyTbDRt6flNDVGaGL1JDYDem4
7x9Dhw0Xk/xoAopbepNErcksvy1wHaNwJVaSUK2CDqx/+wq2cXB7EGKkh86jL4OB
Md6b6MsIGEKNsi1qkugPvUgOFwVAVz8Ld0ukWxBelSCS02XBjSIHDh1Ukz5n5XWk
c7cqyxdwD7klXXvS5u+ek0YB6vV15wNMSSspNGQQgIsoxFg6peqxHo22wT/0RY1N
TYNm4FZ1tQuUlynHeEHl25CzjiyGHuRWoXFtuOBYO9q0F2yQ74yhfBssGrOxjuOy
cSExzPGw0/BD16uMq3tAgBTTcmgT5LxpHU7AFa/FhlUtME+EdHHiTw0URNkZ/mrT
UFkkFxZY6Q8x52L8F4nhjMOvPf+hNrqyzsVe6A3LVWihEkIovZh1V30sCGbxxVNf
I5yY6bqbOUhVdpcZwn7c9PDMQ2EHzIk+nedzEL2MXzjHt4kYm5KMtK/v5d1z1lt4
FSM4SL93T7qoZleyINDHtH0Et73FiRuYUioXmK/qahdnJiFuIP8Am2i0xHXNSgcF
LfHNrhADpuiN4pyA/FcnDcuTm6nrfJ1FiulGxA5vOUw2pYixmfgpMd2yrsbM92XW
HfMDTEtMd8+VdIZlsw3ORzRejF5OUrjQGDjY3Fnw6YmlHkj5Rd+iLZe9ZNuS2EZe
49XzJaW2/mW75Fdw/y0bTEIm+LKNTgCnGarEthsfikYAg+n+ZHIXdj9X1T8w+Mtq
k+8q9nasEuhgAl6XSpacsm+C6V9P9X95KYA3NPaJh71Je374JbasBa2i3x2jSptC
AMe8cd+3604vj7VJuyJ0FCPMaojbZdY0ZxoUtjXT7UOU0Lh9k3IxYQdv8dV3CHOY
Dy/7FtPlTXrDbqn/uKirYS7/SP7avg0A5WY7CQKiBg189ZIgZ918lLWkRs4VLhxV
Fl4OWVVpAsSCVTmDmyvX9faKjYTb/+2YJMoq7Hzp2UwxJrjJKrDf2eslajvNf2sO
3cVUSE76OMLJ33BZ45BPplTGbwhTCIzVOBioJeD7rp1Zjit3S79UVBFDUGvN/vxK
HSq2YwQ0bRHrT8EsgximylXTv2pLawsZ9w2rUa0j0rNreHlwtWQTEz7ic3UJFHR3
344vZjvABxUqSYDvZ7zExXltoRphZ78stbrPuezzIqfkBWkTo8DiDyRlBFUhSv67
od1PkNvz/Z8kF82RGLffh3Z4wHEpPqohUwaUjWkyjOKIhRdu12q0MbdtmEjkzqQw
vQFNON+P69AxB1Ol/pZRBRPhlsff5TUXDdkPkWEEWXCAC7r4097eQFSE09bmvS40
pxkdFd66hGs/qP3+5Y5ezJ/ziTcZJDutZVNaHKF09Y9Ym/3hv7QD5hk8Qal7qn2b
Wau3c2NPBBLuafciGtd8QvSKHFnH3vfELIFC+uu4L/8ptZI+omB/Kg7fa/yVHDZk
vrmBM1eS3B49RPyas9nON9uYqcaIWJJNJDKdpkECQ/EVG3MU3z5cmponGEgx3Wje
RBP69MiEFKe2r/oKUj8uq4jeXCdf9HhbC96TeUFmwEES4z+eNOSxt7SsgzRUPNfb
iTuQjWlLsjrWLrO6okOEiRa87Vokc9UZImNn90u2i0weAj9X3Ndgq3cq4SzLac/u
71ZTAiMwFiuAZ/7B24tcFpooXFEx1wHy0tfBMDd8R/2QPXmaJhGcQG9pfwjDF3fu
9q6DzPMWjgYtcvxRya3I6L++PWxj+Z9JPxzjZU+s48ynTj7XeV+O4TSTteUjmqwx
d2azzt1WNw16StvBDK/ye/NVas0Fz8xZFiyGyg7oVifmQQhHYKH2a+9baBaYBFA7
JdMPJIPo5uVjv0d18CQ8UHc0GrSgIMpIu+aXvSYTPw8sDL9+bDY3hhwZSMBieMHo
KL10EjsyMjzs13WHnUx9xfMiDSR6lAXF/5o56Hj4WjDDnz0vjFzMOgggy7iEK1SV
Uv949/n8rGagkuoxB+KAOtWK3az3qD9pO6CSJUtpsrcZGLA6EVHlwVBMRNx7SrPR
fij9WPJxJbWGwQP70m7DdZ92QpEIO0yx4tFLgsfkfpVA8WNa53fFCCxyoLVm+diK
FnJAIJ71GHH+Owdjxlr0NCBEhVUlhCurz6mNMY7JSbk0guQftsfHSjS7XMdFTrgk
wa52KBWUHbkvq4IBb1A8wHEBl8bYpKN4rkpCn8nopEVh0IK7/taHdcKq+PNH8OXu
EQTj0ytED2wWEzkudeMzwGnxPa1fNiBLPATUfoQe5R8ikYFk1GYIVbS2bBjqr4Je
UAXo7WOEfG9Pigs4vY9zZHSLUcA9uRFA/L0wAuGZw7bn0Z4vpSCFM70G6OKOPrLy
8JAp5/zYBCGktQu0q09RutYzPYtvUJJ9EBSav2IPw02u0T+/F5ub1+SLzbzNz1oA
AnJWGusBW11m8DSNc7T/h85vtp1MDZIUqwlr34/gSa0HvxaHkyo/qKa0xM1WXXWx
auDHLnZKEILlOgrDjJhIeA9pugAs8EBXVaTY0TLXWU6oYQvvfUVY1vFFChlTM7q1
+lImJ2hPG1ZDirKJlrj3zqbw3PzzpJRKCpXMc2cQum42PUPMeul6VvHusyuSABLP
uow7E1vvfwc2p6LbtYvtOZDDGDC2GpuekbPxzhAHvXZV9HhbsMOjLJYBv8qogW/3
EWHIkVtY2WUkWerPPTpbVY2PrYW+3f642/phjgCosgQBnHZLcGm1hmYVEvtp4BMC
xFgdFjpf9J86tM3qpr/vqSPQK1eN8W9lUMXYoWja2ytq7xVBLvIQpB9DgfispjNx
uVhHuCTa0IqGtUoOFMnu16J4ru/amFu2Be/nrzuHv7uXtXrkhadQYIVlx97gAz8h
40/13++D+t4uhKgiY15BBAdAhQOc4r2QvrvsbRkFyQj/yU4gkM6+uPcCY2x92sy5
NKp02GnTgRizJAEhjRYADx0oYtk7pd8w4qDwSKPTSfx66ipnjYMJLn/d3vIM3EYO
O8DdQBIxoHEL1y19RFtALmVfE1H9LQiWMPqPna60oN6MiAr3SQ0CQ7Vs1QIyL73y
Y/yNs10XhJWu3GSiq2+OLo4OiJDLGtMibdtr1rxPghlORtGlazeJddBIFI4mwxgu
nQtuCugsvfFhCb3Lp/iiC0/5u4RRdJPAc28jdKNYy9b788ibm4Tvfc2QCUsOSG6r
Ewm15AWvwPhZ9mcsa1zBJF+Br1SDiP5te+fgO4yLz7BF/njaA1OwniajXlBlfbWj
1a4ychfZ6oj91h4R/Veka+FUlhLxYeaMKu//c9fW1OUSxZwlsZHNQ/JjDpJ9DCGP
El7o1984/T6KV+2rw4bvmsCpWx/3fhgQDTRYRmqRhtlD97iRPuJ1rwPnyEXyO/8R
DSTK6p3h7qAfCOV9R5q7+3VheJrMHl2lkINdIk+zLGavA6/vAI1i5CBzOkhCEQqo
3FGQJ/ERSJAMeQuIHQHHT1W5qS+ZV3XPSvh+jshMXSCBhnfVq5PVHgAVLSp6BOI3
iUVxal2KLbqy9n/QoWouYvvojC+7bG48Xr1OnOx8zDqIN6ihlVvZddW7yBbIfaIz
QeogjDuU2b8D3Cn4diNFiP6IefM+BCEj7Z/OGbjdjkPWrol8KYfPD+pVH4CuBrB6
+VcYrmO5O0ksoLyeEzhbFgkhfFFQrPWMjQ/ojg2on62aRaoW8bphE4L98X7zI+Ct
/1YHdcv3Yko/IQOU2D1HmoK9ZEli2dSiOT0+1Nt3bMuc25N5W8GETFMhfagUozDk
vRfxtYNW2NmkD4AiskiZSRLBYY3xY2VngxedFPlNHfGblIybQd7zfzFA06HzbM7b
KACAhQZqSXOEZTabXM2/lm3PeGi/VHxumyFZ7YCQCqPhrKqVOsFkVwiFRsw+Qqor
+bi/m6YP3mZrRXp/eAEgmNuLPxGwYcubF9eIX9znSjZUDzdx2m0Kzjy75bjGXzAX
rrEjCt1UOS1VBT5mRREaPymoWEERfHQSAVwPBNV+qcZcTVSoQALwCC5wFt9pQ2hK
F3fGBJszUADntOPu7Y4OLq/C/NwQItR/6njGlaFqeOKR9ALB65JmAnP1+HkN341K
yNKKai/p0/wInYcpi/FwBIXn5D+ej3qOXMT7HK8I6G3HFP2777NQQnOqBUZ6WviV
f6vqdyxTdVfLg0qRbGbdk/W1N1YxrAuvtaKa0/hkteA/2yVTO7wmeghplNeFyUbA
CrGmuYhyZPclh3OhBb4CJ1dq/pekdrpzQNxEeEiVF193tkl7aSqw5tcrelTiPz/5
PYO+/mhlxpnvHedobjQSwrChYPM7RKRLFI7jQYVZo8boQjunXD6THEy1ds7dtUp1
5tHy7Q0ALYvs/+H9TNsytbOPSdtPVl5OaAXa1wcl6XQcGNg/h/bFoN6KrWx0opvP
0Q9xyArMBFtYNnCWMtPIH6h9f6Ocs3a4Lafoez5LXnwW5KJc06ANKGuSJYF9Z0pA
CpJ695OU4I9r9634SqD47zwHANJRBrNtycl6G9yDmfm4QT3k9X3MHx2NgAi2CL3I
d7Wx3x8XW9/8XDnLXouCAR1kAne3iiOJqgC8ORUlPWTe4cbvxumR6Fk+Hjr4wEMz
+JYlM3PmefbgKHeR9jqLHjBDFR25ZE49hqVaNm/Ac2GkcOcXm8zPyuIKkclp5EdA
V0wo22YjwqcFWxlN/KLr5lWkKvRt3x8PVY+vPygxQalkHrRLXnRzPvAM4kWoH2Kp
N+zEx68CPYky5nYRthuSG4iwxevqr5dnO81JugyUMhZ1Sye4yPxVARCs052zypzs
RXLASGxyVkbtoAakwt2jye7YU7Rq7dp0zke160gcb2sNCT8FVRdbuRsxoYP8kds8
aUEUR/TNnOIF1u1yH+A7Ts1zpP3uEBLBaKTcPtaUKgz+SvyFV8mfS6jlc1UooTnq
PETgBykls9vwFlMdTlagDkAR6EYBhFnf+UeJ2x3lRrLW97rmmtmYMJ/c5itEGcGn
xAID5IvwSdkLmmpBEADMpwRAQ0jiQkRNrqi26rCxbiWrdlEc2bCSV5sezNKaJDvn
gTkZ2uHY6iOFC0sSAq1QsCvEbQ75oRdacNuegmq3dBb9xF6DOMU6ug1/zCHZNIZR
HdKdpC7fSvosqX2DrAHR7FK0mK/CTO0jWt0p2VFCvvhRN8L+HswwRTnHVDVkh6sZ
U90VdleGTd57mCNuLFdt2pVaUU9O5yp5vx85ejEZNS5WfOHi9eoOzFxQax3lN4ff
WO6wvJ8VuLc4UfkggaIinKWCzk2dBLN1dI7aGZuG2nrTacMlKXsDhwbf9qjG8GcT
MnF/LckbVWP5KJJ2DRxI8T9rjAzh8vjAJndFu5qZR+TmTqZ6/JF6ictcs5W/IkMN
G+61512TXtiks+02Dpm1FT2x6yIfYa8idPAkdc0NWdFzGcwbJT6XS3dBilcNbB7F
RLqFP4KzLzGaUZAe0L2sKtabnOocG1RB2yG8+D3ugUT2Up1YO2KbhfCLEwZ74Ywc
s90gMOPzW7doUsAAQwMUYf4z2o86I9zT/szf4CpMhHSdGuxVv9CAca4y5+ZXfRKs
aqGoLj7CgNMK2NCpgPbRhzzRpNCfrQxr0stdqtF9X22WYGSdYiiZ/yDyJuu/sGId
T2BrzksWlSedk2nOhsU3Sn2Hs8kiEE0c1DAMCSi/vLL0YBUdK9Msvs/a90PauCsT
SJclg2qIgxeQcQ2ajlGG98vJo+qEv7qOT0OJgojUOOXsHPcXXumjBGcKs5MhTj2n
dUSpGgRMq8qSO+FrJ/zCyfkdE0q7sU+AfO5t+hdCLVEloW4Th58Y0LDYMFby7SEq
KjXS3rZspY59GPy3G97TPUAw0QwouvlAERqcoylAyb2lUii+HzjNA3g2nC8Trbz/
qHJVgdvuTVf6OEkWwVfQaUSOVCKH+d600Vofvo7/40EZxvhPeXzs3xjRqlOIlcLP
zwPCqJD7NS8K0VQ3Uy+iffkSEzj++OwFLGCuJqzn/t0iag2P94ML4XA6LanGAD8J
eNpnZA9jaexsNrV3zXNtUCaNeE6kgSLG/Lg3i0ioi7aquoPSz7E1FE/XKJnpfZHY
lrozSSbTp3deN/GQWuOdejnppf4fuPDQFG0Ah3Uqnls3AnuBILnyrzQrFS10lu5m
D6q/Sr9BVTWHNecP/AzdkMXOrF9mkxWOxmSU5MTIYtGNR4z9+44isskMW1pl/Voy
beFYl9CP+jEksXCfnpu9Nv95D7cUKhjhpC+5B/SlCvqdECUHxfH7l1XGttg/UjB7
FWSJsyQIuSg0vys7SnTubw1ElVEBNbNGufrxUuQVoUwyCQF8AhxTL+7W89GbtB+8
ebEw5C7g/4d+am4HKIKSaizPqhOYhlwIIIIjAGeq4SjbYeipX8Qj7yuFAjyfsrbx
D+7E8ba+19Xrh80Eo15ddIfFloZFy8QIWtFuhd+FRF4w70o4EGLlqdA51UT6mMoW
5CVlIlwEwlg0v7m5NERnBaXxFOvjkH5NWv1bAM6WO1znkJk/hw7g0quxjvlp2ZLx
Q9tjBlZR470HKypYwwnUQkCkqjkz02hNceR+USqvdocUsTjD3Q2SNrmReKkShamx
HPemkqaleWMp8TEEIZClnHtpzy9xkhpb3x6+XpRDXCg7pHeUelHH92e5xsyiIX3q
JlIRMEoYrFRKtBb9NB9UpE6e6moNxQMTQH1/P5M6NXf8gFb09+jNsx5fC6RSyG4R
tqjy4lQBXwePuH4PehwCpjR0G81USMNG8r59j3lOrJVwPjHqsZ0lr2lEE+oubuLH
6Pru8HcPT48UA+5ap1+5ILbayTPg8BSGUwNPs9NlUnrEItpQd8PG0O0scWQpvNXq
3jdljdFeNtc03J0R4hyHb4K42hB1CWfjSEBFh8Su/Bs5ngtUMnLQyQt3rAHprIi5
5JONuKzkCsqnNCFL4Cl4diD21U07jTyFLYaX3GJytA4TiwcQs0Z9SXfrMLXRzKQr
u5+vOzmU6mzHOkTYa0nT02MADVxxgJ1V+RKjBugtjnUaK4pQ+gLFhJcZk6Bu2M57
dSacMAQJ1sf/P1S1rlVU0uPQL2G7ETc90ShCnpismnlckAsrEb/Cp2fTdOCvzw0p
fSJTy6qzjG9htyDiYIxfTNAFenlfN8tVmmk1VJHgvzV19CyovI6vAtnPNcs1aAy9
bsCerR99Nm6l8DUvF0ijjYPodDxRKaEmsgQn4UNUYwVJoak8fMsJCwxhmkgyMa1M
jlVOu4TDxzGybGKXCY6xIbyL42Ko5MXh4PWOQXrNKKn9siyjOQ7/yAfJPEsqCtyf
uo9dtWLQDo3eWdgNbCGy/PhLW/kOjVvi4UhRCFsXHoGXKNXjhBomt28hrO/YGpN1
FoWjCOya3Rt76AJUk3hTN49rbGub4PDp37RSOCVcPn7qs36xSw2htOFq2cdaK4n2
b1fc1TwlqOv9q9VCWpaqYOAO0xvu5MEOI7IvRQXu8kQSXELRI98PCH8O2yghHqBy
vRS5nNq2yH3hSZdPidsMxgKzCjqVJGxcrN2CxfN31GaYXeOzsHSEsCOrasr3t99+
x+dV/Pn8VaB9lLA/Rn9TWCszjRwGJHcdhz/ILBwRQkDv1eNo8BSaE8I973XyHgV2
vcw7+WrNikJuvM5V+VSwHsT+H61mn5IC5Anqbcv9RTJecoCLr06BMl6i7+evd9Dn
WHROjmHDjhJcdK1NohioQ8US+s6sHx8Cn6Sq33BLWpF2WOjZwyvObNHjOXCINNjE
mgzWmLzNDsEg64JXZWJHVkSId03yG0H/DiPcKPZ5pMClpYac959aKHZV5eS/QhQK
hfJfjKTSeiuZALFJHh9E2a7Rakq04p/qd2JYG6AAHu0G+qg8yMwHJQTvNtAN31XI
giTyxoG10Tgs4jltodJxwu+NzsLKdB7whiP65ErIhEsILHbpXjq8CSjZBFRs7bcA
QHR+chXWn/4Ta7ydMbKj8p93uJ+sdaKZ4ryzqYXk6k7ZEQDwjfHwy/U6F5al3OEl
g5hlajnZFRpKdkZuv+Kc4xvM6qR+f8TGb9XYgx+qeaX8iLc/uwXEtA+KVSeuM9Oc
QhpDd33jRr5z+zV9ljfQc+6530iBSWCx/eBh1FUJlxuWwmrkcrs5qqaxp1Rot8O5
UImmbS7kGRk8h8oVVwIxgaUEC4AAu7GWTGGb5kABCEY6IgTPNafXwcfLQ8n/9Pxy
zO+THgKLveOKkU3Mj5X33Dt1acXDXCm6SGek37ukY5QwsoIyKOf8rsZjdcxtTaWU
M+FO4kEbLY1mTarY7aukOKrBWgaPz8Nl5EsqOflb/CobWZetJFcVvoOc2/k2Zl64
tlUW2QaWX01WlIkiE7k0ws9qT2azLO4TDcVK83zTGEeU6p6DUwBlu9Jg/9J8Vw4B
6S+WpN0G8CjPcD7andghuKD2uH2SkptB0YzlZVu6AoRKOekrVQo5Qrz0Kg+4u+5Y
Q5gbAI0G/VsazuT+M8hdc3Yw91004BqmlU+ElWs7x58xxHA02wwPnUvkzXZU3DaX
4aXrFIfmb54awr5MO3tr+9uAm+7fI/lWfX+mAUV6p0cYybZciQGtE6+c+vNMIXl2
BTDzrSLwoodxLwK7s3lt/iGQaTCb1sJ4/V6sGAbTZKlYou+Jvv9O1ndKdjdKXs0Q
9laP+1Qjvy+wuHORzJffLZlUFwQyD3VL/0ufcM3E3Y896RTYOOhAwgomLLsDNwVQ
o23jfZlLWDvHJ0u6VXHOZPXSLYJwNsjF2dChlVe2UrRo1sE209mG6Jm2+5wGr0/A
A94I4NzZMP2zJZHovIc5a2JWm7w+sGSolYBZe+ClV2dSC5lNHLPdWVvOQpIBaCit
CdFGte6okbpuelZcK1JLUs4IVc/JBy80UrPC1WQvf6OIY3nvHyam6T/pYmpubMni
J/tvA5bMhrmMkeEI1tFGGDKVOxy81p7Hk9Lh1okIJD7Rd8+suWnw1QL8twke8lw6
B0s7CQehaBC8TL8xDx8LzmCNSuMS+dF0a9lx+q2Hszd7GEbqimRfeXMZriGOdtyN
lNU+o3MEVzP6YhMKOtfmnCCSSpoGWzF9WcHd5dDHK8B2fEDNDGSG4/AF+xNM0nur
acEzgqcxPwbMfuKW6IvDsRkzwLemC4kD78wzYmZuJRzpF5U2e+6miU1R3NXMr7yx
N0A9P1qYLl1oqxpmW/o6SusBTwxOFUMGp+AQiHhblyxvpu3RTDGCk7JgCQvRmtbh
9X+MyKQRQKmWU8mVFSAqlbmKu83QDXpUwXQ7w2HVXzMHw4/gdqhDP9s+Y3L1U4mc
gjSBXY7moNlxCkViVx2BLOvw8PehsAbynAT+wau/2mDBEuD1VrYyyjIlnQeWXM7O
Qb2CmfoneXCtA5ecAXjXwOgElrhqV5qSLlsb7KDSLCsDMZFSRcLQ0vBVsAiaQ61L
gVc5IpQwhisyxE0ompjsobzrtJHGWNsDljHZmKpTFKm4ZqMb+UtyTDW0K8iosVdf
mKTxkfScXfFJ6qTLvwRhHoXCTofiNP4NlZ0PBcGx53oOARm8h4FTKdMolNeX0PLb
kxjkqYGwhZFVTcEwBTikUOZNwercy0wEUbINUIlwbyxIBQ9y0/H8P6TIy8ijzYFG
d0R0ulr9xFD/yqkPy9e53INgZZxO0/3nGqBvpZTqqc8VNAGmL7I3vKngJx8dnIpT
0ygYwlT2ngDfKn5FzSiK/9T/iwVtclQblOcfZCze/sDR5MCgQE9hOOBQqRvd/2rq
+AVraj6eL6sHbfY3REDA0mfZZYPo0+A80blH2+/qUp1rJDndMGuuxc11+1TBgdqk
InMlQTJ62ARQYJ+piie2gVsStaKP5vYzmxsG4GhAZpnL6L24CQ7QeSSu0yiABIvR
xY2PM0bMsgCpBbFa787xq4X2oNT8WjW6UbVUmBdugVmm7HsyIYk/9OJRPM25cy9x
vxKraw4RchyLy4ULGfD7vCUVY++bRkHbIAP0rLGE721flWb2tIQwLUMDn/Ja3bpm
OV0YP75aBOg47RF0mtPmQxg13mf+kWYH/KOlBD1ZHJiqSCbmATobeWD0IcF/UJFT
/HdRzOs99JI9/iKuD0d8O5AQHtb8UfS9FeFuTA8NjDy87LHAHdpBN9UkjqoB1Wk+
Fzivxtgqz5NLuWvoVta0WjVTsxeDuJzUpZJSp/rj2RK9vZXmY1XeLxPh4n8B2+X5
YnKW6z7kzLoccBqi4qX8jrUbYlhjIfhqQWrdcvIWJBaVSbmHoJy/2xoSpJJwEVtg
pglVfgNMgpW8Tkpq5A3dkzHU5woTkfESAi3UzzRTL1sp+zxdm2l59TbILslj623X
qBgmgLvFzKpRMUPdtgL5n/aWVXDx0Pjnf0nbbD65AeBHu46Y4pecLLc9S3Oxgj/p
2DxqsH38NUF5JF3gWHjcLuoJBFNc4llKe6wDTDzeOfu/3HSwjicU9IRsl8J2/xoC
O96jGb0ED/s+VT9MAuHFNs/3m95y62zNTAF8lVt8B0ruEfotsSrfhCAgrlt/cry8
/wMECjjjUnzvzhoacDXI0D8p7UYD2J4nUAjxxZuggMl+CpftqboZR8cGrqPMLAGB
l1bVzcGNXGv3giNs9uGJr8Qd04dMwYEab2fm/w35OcptMnaC7ns+bRp/nKEiaQuB
4/4dcQ8RTWRAYx6/hdq66PQEOdOMqP5xdlenNq3Iqew1QeBEwjmXgRAS08+cMlG5
ICks7WAUt8kbjI983kADaNKXrB08ZO9HXdagYDfig/FZK12OiOJ/+90fyB/fuLvF
u1ax7kGn2X4wGpTGVQxmaDCNe6CVhxJZ5Ls67M1CBM8Zk86AG/VZabSBW3HuqaxN
pKYzFYANWCoiV1uE1cj+sBbbfCpP4J4EUqzPM8E8qQ0cCHspju5vXzMuQ8uez6J/
FM5ddIgFXp000rYARJdxxsvPb9fGDaivDWa+gggC5474H6jFsPKwibmHyFbBNXwV
pS99+meLhujHrC+mThuBk5yPqigudRR1LIwp2iK1FDFmU/e7HCKCPkHaegq6Ngfd
lYooTaTWWR/Adcnjkm6AwhCp+zFdTifcxnI/aIjniUrC6km0H55BM3heP0ZDtewI
ROGcOeGbU8gkUqxDdsf9TLDYeALfWI7kR3+M97FX6mDn1NFNR0xaJineg1ScIGLo
wjkvVIPAyNMLlUupa68JXdeDkwqY/jbcI3H7AOfrFK91t8vyMpD6NjgPQUS90XqX
TVfJIunGh+3LyYevUaiEMG2UU9WpbzJ/AfG4XduJzqfrma1Szk6vzRpiaqI6c1Si
SZC1DqhjQOUyGunKEh2CeXQwOpbFX2g+mCR5I9cdDzmB0KTU7CckBYa6Q9PBpnfD
D7Zg1Tf2+jrJUxsrfy4rYDQ4BSxaG66r5uKj/hSxI/wdtLrQtztVsRSO02VBxIHd
fzWV7S2JGBai3vqevivmvexfTCsjlcKjUMTWioRcRvIeWP4AK04HvgqsLzKvKZiA
0ymbZNxXlhJ22Rs7xCMX5YbViroEBKzsgE5wcrQwtuIHlUro2FinBJMhVxZNT4Kw
kH2E/ZaFTa66OpQl1tKST2RWKnyW5oBH3L/2ApRhJezdY9llWcsOXHsfV0MWqYV+
9/VKN7nrM4MOzvsRUkQEB85Fi6YrCelxzlk1O6IboRMW/m8saEOl5kV/u7jEvUYq
BwwRKYOsLvBW5GhdhgHXiAHZDAPkMzO17YTdiP1ohv7YiMvy5Bd8H6Rxk1b/YWxo
Zw3Aexz9VtAgrJg+NGz88JVTwomi1krrA+S0aOS2yGhFow7l78Cq0V6RYAVrDaTn
wSkeLLGODlDCy7KRk5naRtjokRh2s9TnyMHi3JJlqmXL/nMOrpsdM7GySyzldAAS
caqdEL3hZlE+CZvBJ54IRH7AzJX3qfaEpa0dq3PBQHjsF1nTWmMPfDU8xnbCJUkj
sH8/aXqQ71Zv7+e5QS4mcL4BfRno+q4uJbiZQB1bshuyET+3NdcKndtx+hJ5p4On
FTc2cGtqK9Ekt5aFGD/9cNtAtfbKss2ymVhp9iGhhL0E6Ny4Gk1CCpBWKpOZiO/4
wL7Yq6vDlgfqNSsjn/RejM8n4dK7LhAtx6FxqKwIIdbT8ydgvXigW5PCQPo+p22Y
/tHdfL3/7/qSixAMV4bh5KYYoeunovq5ymTfKqgUP1mZVh12TuENJxNrp4AvvgpZ
4+VilEmZZuEvSXf5/7CendQhtZgAddnENac+SthuYDIZTxt82Owu0LNKlQ486p6F
zAKGs1xN9gRfKFl+LTDBbNH80amcyT4zJ2QivRacFDv9I6jV61iSCG5rXal9Q5+I
/KJHo24R3S8VeNz2nR0ccnM7UDie78t9tnpBD8+EVHyjf2fnq1BdPi9G8SNN9Tla
rxT/tpP54gPP0Pk0dvOE80jifrjmzQgywYA+QIpWV1JVeYg6AHmwhpUPKSw6a1cL
4blp1UmXvAmpk5REHoZCGZn+eJTpIWVHjCYSEce4lX2aznWZnhxBfqJMEPz9g2Kf
QdPZnd/CjOyYFzDDef/BpDXN9uODWcVTQG/N7s/XaF3vOAoVy96x+3VfzzLzeEPa
B3P+K88dbOLYEsGSVdAEDoPC6YGt1kNOEiXnXkC0Qw5wk2w49IMvfGXdalDAg+gY
F6TWWup8KJF6Xc4PhVx9i4/2pE5dM50hsikYJxMFcFGqzuDFgv5o5op54JCQ0DMa
fy6/4m8qXeP/GH1vWCbYAySQwYXDc7GoabT85tD+OlBnTITZYy/JjymyHl1VSsXS
fDurCVhy5QhpH3baTP5af44Zb2gv9Hd7X9eRkio/w66OzITU37ttduwLb1xg/+my
3YcgwzFkn2/tbLP9pE/A0I/Snc0nS3uuSOl3N5xcF40WtPP9mee3tTpdiwN6o0I8
di0FRnbBf9R2Im12wmh5CAD0UcSe+QJhIOGAPwoAs794Auumc1Y6cq4/qm+wRJaM
rWJjjvyzoMk5l91oJUexWEHwgCJaqzkkiXZhaMNLJK5pmnip4ix6kv6IecErfFnS
lTw73KGbX9QNPYn2eicFXQfH3HGbv41LcYNvrt/US2cPRJKAq25kDNdhYYNiSCiH
3Sb5Qgr1RXLAq6VAA6psdK1LkOuKf1bmInwP2ZVQhZXKwZL8XfTzyZtJQ6O+EiV9
RAqSnA+13J6G9ZP07b8QLgZCGVKZfaxzzGw+csxDcV3nbPXW/pES8vZD3scpJ0rq
Z1FvzLijSciw4+BCjv7pWzSjtyteI9KqqoS30t1BH6kVGlzVzH8bNbko4ibKtrrD
1Q5Ik7yGJ5MvoLCS4Z53Q4N8FfqyKflF+dS1NphcGoK15jAvhyfIieK+J8FBnuWb
MNkQHZT+SbA6w5qK9SGhrfOWDYRzhVuipJWgbQ6LNiDCNa4UXBWL7afuAAEA2KmV
vPRCpnUM9UxJF3tNTP0TjbC/yysOyHOp6CWuoXgLE42xcZInc4xCyriGI0KdZIv3
fYF6JUhweqOHvMEokyTJZpqpRfQgi1C5GLCpTN1RxxwgI+OzATkWR6qXb1JZTDUF
Li8Z+REP8C3TtjH3RaiJdWFL0uBFNiRLR8l3xoSzcvQ765xkBJ4UM603Y0JbtGVO
7TMm6zX3FXas0X4gZWDHemyUhBdUWL3RWUTp2429sES9qKp8vHaxKgJjGRAadwbp
BSQlpK4Fdyh74b8rMazTr27hFHywEKaA51z3xRXO6jdCuOoZFArNLE4+GfN9OV0v
HLQuLDxFFeVwcMQv84MBRCXmzWcYzS91rdDiR+wAazw3LOUF0lfaR0oHBD8wYnd6
VaNb9LnFMYBGCxUHhb6IarqX6zvVqxDEKnPVA5f59POa496TKaNtS5iETl+8eoEa
hUl2YMu0cwp+bT2WBm6ZW2zjVEFWBiQjJyHtmBtUXz7lLHC1KvyWqJ3b8nIxD7Xx
Ne+AIyINfuuX9mebF2wxkFEgv/Svj/8rtG4eWCe3RzmoG+b9jO/os9eBkng8xpch
wOXJA7QzLdGUuPuEr785LMjJWwkFIqE+zm6qzJ0Nj6528XztF5OH/r9nwI5+NFoc
iY1CrOdYVNQsgyMB0fVXVLa5+61PGg6l8RF/URj9F1PKqj8zPmS0mnic01pidMeC
pENwmWmuERYGv+zpa4LxoHoJcGiqW7N17DhXffHWp62pJskvEhO5rgfMpNoiseAd
mNw6qQ9UJQOYQeMm00kxanSeE2bsPeDaunqtvRPioZIF6hDBnKcJIpyCx2W5X9oH
lPxd7kL5D9Zlqs5gkGmZfhxqmSyfVMpXOzcn9aet30U/+0qkHT0XC5b6FHhLj87B
46EvuEPn3zKANJKdzcQM2pe3pUFOP4hxoJXhCakqgmJS7POtkBAKciXded4bInJZ
5reXaXYrwJlPKp7n2C+j7e1ZotY8IY76S72Xahv6KxW87EXA2ZDItkm6EVrOHqIi
DsNdUfq2sGgUFmODZDDxXyUpbVb5eRExdV6/VLVaOLi0lGoUrOk/eGq8u5CU0pM/
wCFf30JK1gBzM3jgkaNGZYXcCxw+76sitoMAZ4ubpN2uY/sUbhF01NspxQ9S7rwN
exM4/n8rjkEUrOProIItwRpGaZW/edbbV4m7dQrk2PikMkpho4xOTS0r/WiD87N3
4RWuTLRhupQzBkjeNXYf9F5r852OGBT26B9RauXFc8Vu92NXwsmlhUGEQbKIHB6r
rS7XL8z7O+vlQd+b0KNdLAqTgQU4P/CxS3Tw0GyT1z3y6JJvcr5NjcMzKjqUY/rS
/Q9daMH3aRLrVSoVJUNOHJMcMztEHpNP4TczYP1cdQIZFeIJT46BE17hEqJELgD1
qC+uFlMQ4GReaej98MlHFRSscpuPAbus4UxZ/nDf5lehMaPSPRrYSTI9e+hOcW52
Ea5ybRUOJadfnxZopteFImS/5uTOeLeKqfEGZnWdKO97y9AXwXFWSOtHkPuEdbjD
UrFzpWPiNgyHiEKPGyS0KN9ZKWi+I1Z3T5WMcnkcTKGhvwWLiJFewJWwlxiNR6vd
CVzmyv0q9YzOKuCIRUIa3GA2ZHW4sisOt8V5MI2hToeigFzTdL2t4/8TgXzgfITm
17105++8e2kCoMn3tasXh/6jlEXctILHnvjWIye1wjCVibpz+mwdoTqxfa1bFKpB
1PeAZKnkLKG/4G0lwzfyKZ3m3/BSD1pgyW/vH1AFso79p864R82eSWA4DiXtg1Jb
TEBVYYPTpq06uFVlYmX83fcuq0grzy5t3mOVfNKUUQbr+t1leQZ1Ap7yH/fpKmm+
EFLF0FAEDFHi187S8D+vZ+AadTNgudPr/OhDG3fZPPznlsAxfbrrMTI+iXFSFgxi
ZLaJREHJNUFE322eQ65xqWh70eaYScYAs/ivvnRk+bVHn47z5aJkgGVWUoNuCVSl
AWiqircD7LavbK0e7zyanGke9yJcc6zuhCwIhe36qFL/801gYx2yKACn6X7fblQp
b43eBy2RJCNG9OlWDKLhqTN3OQhow7MXS21TL5MKv7T+LFcjmDED06jCs/fP5BIc
xFocZMo/zmiki/l+oN6ks6NdkO/t+7zJ8L3zRRmTdWSKzVBYGvAazEcAjmDJ92vH
lYDSPkT3GGn/Ro1Aeq8ZOiLR9eHVWj7NXeeep0rGq7a/xJPlvn2QfCbtO7oaP3k4
olyYYZdZxucYVxbPnbBSjOn1gmQzhdeJRqPCbbTRziEVmDFQW6rxH7XXDYr40zxB
Ik3yZhcVwjuXzYB1hk7ylC6h/YYMcEkTqY0rSa2ypgp1BIRR/wreoTg8EsRyTfpO
f2fGL3amnMkFSXkehtsnJG1LZufAYfkLj3AlbOTLl5LouRHh6OmA4kWWxvcmkmx0
nPh/a3uyXEO9NwB96BMKq9p5A8JvoN/A3nAtCtjJzfKcA4/Z84uyFmbxza7Q6H79
ymRnSkkEulA8guLEJPEkwgNRsqL8oIrRs1Ji0R4o0SGBJCmGdOw0G+QnibGauDuN
wUTVngyH0UStmX4GX2RI+T2RriFTw0bwxHnZ2pnTZZZU2/p9VShQTad8EpFxpuHg
oesgbz1mjYsSs1WhG4DSJuIzI49LbYH/5lUHYyl+5dECC8Tj3+NhIYEYBzQpivIN
PAl2wIY/cH5fbLChH31m3/SYZB5XAtXS30YOv3ud72EeGgm13+E2wfCeHn9C5hcA
z11dPhUsSh4AOkGZK9I9VZc09eVG8dbcwFbjrl0JlcB1gKyFtdiN7YIOb55+pPrP
qIMsumlVR2VcszGa+qa1Vz/Ppw1ReXeD+G8thJyE8HkiCf4QDlAApQNxfEL34Nyu
u9N0hb1XNvc87aZNp9e9SkhKo8WTkrgHgnc9iNtD3sQW1YGMD5rPqOqqQG0LFbMj
nMrhR+YL4AReUOODELCqIvb7KGvVVDJNaOG9iYRwX6ohSV6MaX2J98LLIyn2+MPP
nKtY88Ha4/YiW+SBSMdbxBdeDIzq1VJbp7orALqGv8HrVsBdV236u+buMlFcc71J
RnNBKlqCOga6vrtJYuupEq6fJJHQgbEWOcwtYsImtCgWFKz7Yajr5v8sCeRypugk
dAMuMqEpseLtf/aCf0m3TzJda6gmXiu6/azx8O9Mau7BkwEP2Er7di6KYYqyhEB9
XnaY32WPUhzl5BZIZyJZwdC5Sc9IJ+YT00+9S+fHppoa8o1EryDRNcDwIqmSMFNN
NkU9NRiqZvTH7NbIfXWltxFKdG0s3h39JFAd5qodSWEoz1QXkgf/C/HvLauX2JkF
zGr+/17vMsLIb5qPzMDmN+efN4/Xm40vQJO29yJq97oz19yS3opEsA4vtupZ5U44
+WZcJEc5OvZTJrmtazqB6bTMEmjPwq4fsLIapDoPyI/Z20Nbl66YXr7N7LEvUW9b
eHwYWi2xxlVldre6zq/8J+QEf4ByVNCCUuIs5SdvcXqyWzJRjrQRAtrZrU1QbrRC
Bmv0FEQyrdWy46LDk0SjkCsp5xR6qY9mw8gGsoxQuiUJ0VQcQVcwy/zFAh/w/MEx
vXa1HLIZa/4u1sf+hf+Kok+zFy3BxmDQbbYKLo4CiWHpzMf+iGukD7S3lb0srBbI
2GODrF10PvUGtD7pNLtRY4LG9cf89SW8hWsHVph/EG4Kk6HzRUtNUN5HQTysSsuU
583UutFEyEb0Sl0sPolE+GA5+pRsKjuHwsB6UfETQL/+HV+JqpB9mQ+J/G+hiKpv
bqOpmXzF40EP/+WOWfdWtJn6bisopqmag1QFF3XR83d3P5PMFPzRW6G8m5qZ8TSj
tzA2BsjtSlwpVNifiqf6K9AbhkWnEPsrmZkWaGuqGoGSnamhi+IPUqus5djEHgRF
lJaJE89jk4zQsBReWlDyACZkasSrql8/T+VHydkV8+5sYoOD3tB6PWv5vM+2P7Ij
LnvsX9lWqWJNLIAWXdQq5DQakIWsjAxFKygphWjbd9tiOIq70KbJSiitzesXx6Sc
uXlgB3BjT/pK5mSI4M6XQjUmuqaahBqq3xljSvfFc6Yx4XbmjLsW+gN1vGhxWKnr
W0PMu9WGi2FPDtzeBPKg0TnT0QcVBuXHcXrGTvzOMoZZKRL7Nq1C02k6WYxuy/fK
Q6ReM4O8tsXMExGa3A+vYJ8vhqNHcpFFWbzr5SDEwQG38IRisuP+KES2T1ROESqY
d2fr9w7OtHkBQCX7mXy+GJGfMfCHIYnakT9EkVyfM0bYS5qeA2hGIxVINrpOTzTu
BUaj0fvHFGNQJI/bdUkKpWUn0uF1R0paUdcuRUahw7rA5sbuc4yKzhEYOzqZkGYM
E9/ZjFElw3RIpHEIB1ejRey3d2xXDxKZcrNyEj7P+GtNBjP/7lHVBCwvK759lpTy
cpoO8KACQFIl6dFTKs+qsFa8+5q36Wm80BDbREv+SvH7QfELwkDth11Y3RffSLmz
OfUYV0dnnhXmLK8yw8gDgqlHHB2phdhDApuaPnAxMvjRQqdZum4snJZX4cLKG9v0
NpGTuc4HXLBiN8ICJDv2SDWUCKUzXdRO0MF2ssTEpWZ0DrJYWbxZMfU4hKnjGvmc
tT5fWhlz8Wl5fPjMWV6IxYnbpRAG8HtfZlSlIqvpLDXfy2fA1QabcFwT7a5xpFxI
VFEy+oNK8gpLjLC9Sd6XbsVPKUvmT1GRMsT019TOm5Phh0sBun/EqAd6MX+8O6kk
Lx8DbWNjJ0qfqKu/33Muq1Q29uueZAew84NPiYEmvffZcoWqpK/yaOG5Ma57bitJ
ZvFbCPs644mltBHgZ2piKhqAX8E7RMkbctckcg+PPVw7ROhK+VYuGL1iAhOHmw36
jE04nsaKveSVrxu2kDSJReG7aUu1ZXWmNCB/R5ig6KsCkNQQXNGEs3/CgN3Ww1Oq
d8Vu1NaMPglTjOos9cy1okIAUJ2aJds5dff1k206+Yw4GqNntJ96zAQHSlcyi9rg
EFKNbmW/OPLCTj8Z8jGbYoZarYbQHL08LP1ER2+IIMsVBIPruGXdeo3PfEyxMD9Y
cFqjNWz3r9TM3xC1O0kBobkbuotu3Z0oVc+qDMKFCY4xuvwddiSO81joPM+lvIxB
dPP+vPHyJBbaN1zL28bAxsvvgDyV4uLRNXnrOqkeMbboXGFmhhAC/RlLGNxVvfmv
e54glKXo88hrG6JdvsUx0oXyuAAROCtpJIldAHsmoIT8X3LMUP3ebjzeiou1DUrm
qkdXQvHXMT12Abf2aZYCfez/rAjqQbdU2wveUz9jg6rWse/mN09gknvyq05oIogk
zjc2ZW86+z8qw0wjz60XvuJIuxGrPc+0qlnSGiLh2EMYKUKTtkWHaUe8tU15DsQR
TER06b6jru9hbsDnFFffh1is17Pfz97PFC4JdPDumhZSvxL+Lce+9LIogBFM9e7U
Kip9PicyvOotnx8a4WI3iT3aDnNC9lzDrgGkrGD03lMj1iWs1ZGBagZ1d/wWsqBV
DAh5OmFNdZQxvOrVq9vYdtOsUOZcxwLTjvrp0hT7mDBnv4Otq4AhFotFGCOyBh16
CPnXoMtdfuMeXnDHoe/l99Yz7p4c9zg8L0SF+voiyVTdMYQTmTgW7cgXCrq8KoYT
Z9GpyoY5LjV4wEUkk7hK7DMJs+/za3uUlFIM9TuXU9fDb/ejlDdijkY71u6EwSIo
5ewG6fYbKMwR9mIWRi0qpvmuGQfOfLle2C/5t7odkyOFYicT2M1UoWrPuvuBOofi
RgoIBrHXAKRCm5i08zE2OHhOyO3vbH9/TMC2Eowpz+kCNF08b0dJ3wJ6WLJnb9bw
A55Kp9sIcFVTCc/94inHUlFNzqsvmqnQzzqm3haV+F7eaupb6YKCvOMul76xLXko
VYd780lwp1Il/a5Tzd4KAPcbIMT4TDBE7F00f54Nur4B6NJWdDKTItVkwGToL303
xAaDugpuFbWQy1jQkWA4FEwSlz99smO6N8sqSXKyoMJKUtvEKaEupeAN5/l6X413
xLcajSnmkiSyYZbsZPub4xjR7VtzSd42Zx37tXNJ+4demYmYXC/tTLcx+8iwxfGV
3O8JIXzjHS9mOxozLZ5BJwKScilw0R6P1C2OJAOtm5PrwYqnPjcTnLWmmXwSY6QI
i5XPuOxPc1hQ7MsdxZUedmV715HuyoxXc+2nZ23PPdseU+4Ko72quWnukN0Bqe4Q
X7HXoH+jtUxjCf/PKptBjCWg0ai0NvVMLcBCjLhXjdb5RjlrT7p7X2atjLBTlPaU
i1tg/QwaW2tRuQ2hyp7i6wxbwMKBDoKc8PCe09HkaTS86AByLr2SUHywGHAKs1Hs
RzdqnbdIbgK+ybb8xi/vkC2k4xUvnP5fz0PA63+2uWMIRFIokUEXwjxUjKSz+d1F
G6/lMANleZdKC737W4mW8v+E3tSo81DpvvmR3JZ5o3g4Fc9Cy9RcxEN0aYMCKQM/
/QqcAXXKAWOu3Rg+dhU4BZE0pDnhESowy2hgMgOD5/8fvCrhL+4Jt+MxGrsnCiqx
hxkrcLOJZFn6mFwH4AuRtWsvkI5XeoXBIeZfmEFXLWfD2VI2DLF0Ch3uqELWqXgr
wGVi+gqKXWoi61NM7uGRLOsDEJbunZQaapnoY8R+xhaF+abAV24Tkfuc/g9naw/J
KkfeYNSSOOGcLaxUFS83hJRkzlVRYNtA8mC5ZTdNw+KMcYBSLzOCNYkD9BrICaCf
2eMEmiZkUKyx+7ILZrGeL2oVr7qvH4PCVxykughNBo+fti3n3IFTZ2UzZEHZ1W6M
LHuNEjawWtThVTVTyGhrrQbCEFCvmT8pd9r4g+ktmEGhWic9zPPicFeYIuKEhk/i
gBiI0yjITJn+vORYyj3VpABk22LVQLvzRrxf7A69QCcpY7nUIZB2XG/C6cjS8Gjc
rgODfDI4ucUaAvIht0Fv1+Ii4r6pbBVkl85xpdCZJuKD9NK1fCqIoJMHZddzACU8
WxvO6RbGbgp0/+qNFDoQFwrTfFOkyxGZrSiuxlfeu8dQFVMTcUaLwBjsoEMZCnQR
yhUmjqE3UA0CatBz4YA0xhEohKQzy7VGnQ6Kb/Mgcg1Z3nnHKfc3OmY8j/FuczCk
w5a8E5lN9vKOQCsw9s0FP81UN2PWzThIiVjy+0UzH2TfW//9di8D6ivqvpKvrUDD
OdMaKNJyPmsC/6oXh9jvLhLjpfpVFr/augj7PXKLTPs95Sa2WmPsDcJnqnapFW/w
JZgItXJxWCN9Z6hWsoLxhBv85yC2m9St3Qpr2W7qo2EDqxBkriB0YlbhDSjbAOKb
MPc215T3bX6aXFrTSXb8HwMVtvNgRIxHAGiEWltzdVeJo0EpL2i/OARHGYeyIWIT
asDaByHO5udK+1aw+x6X+Ism668W/dcDZ20TIZCTsPD3kxWkfgQbGcZbEyqoiaIE
Ww59bbqG6YdP1r1cEWcoe2vbo7eC8gl7DkKpTGLWGirFngh36/aWdKV3Mihreqo6
dtGISPOQk+IS62mIdrM7yened64SlazYy20Bwrhlxk6TduYH/DlyibRuHG5vUwSW
jWI+xK2DPhMPFk9FeeFEf1jT/yO7upF3cG63SrW1CrNFTWVlzB817uKeOWsze0uz
vvspRHLWlsr4CAgs2kzeuJJAlKn+x4qdIn9pxG7hDJ/D8qh26kDRbHtwFILPss9Z
EArLKiJ9aPp0Zju0//twHBEiM/I9hnXCJQYvBwWEupdSnHsqEw8j+lwEzD7ubgLQ
JVkzBpLYpy4F4ZAMIqXxlU1gHkO9rFSIjo9vDmrto402qhaYcEreTdkTjUthz63i
YoxnTh9sZWRMtw5Th/wMbxDXZD3FxsJx+e1sI/woHCnNzLSAjuE0O6XRuxM6kcSq
KryZ+qdb23irknh+ziULxs1NPTieeuKdJetATFynPDtU0//KyShz9+lO/u8xW9oj
tX8bLJdv62bH3nt6Hp5w9loY0KT9XCndD6f9Ji/6cGU8mFtq5wFSSEauKUA+4aiU
3uM9bE2hnviMX+2gjLMzeR9rC5EZNXuljEHmpZAwZzAKf1hzWCEvABrlth364nfd
Nlh31in/tSu0d4Zhz52FZDlkIloPOf1CXgpaIHaU8u2adv3S29szuOzIniSW+FlD
jxDFY83Ss+mXxrl40KgdpZ2VlNL+GeRBNaQAjZKx2X+9K8Cdi4pT69IBcwGaXtPo
Ul8yDQkylPsHLxudTSt26U2bnusgT4wlXXoXx1jL4fZb5wIGNQt2cKg5YIhfFl+n
fREve/Eptw+eXHPx0nQIWmtHt6rmTrGh1kZ/43i7oUhBFAbuMMttZ8288cNiaee4
H0q3JjKVRatYpv/vVp6qMkcxlgUO4ES0UZIZoIVpVcbbDCGxGnPaiV/I2Vls/Kw2
JSIY6BGVnYX3dDjxRnavUzCG5hm2zXlHJ0RgIv+J3xFKXh9L1kKX0QpEU7Dg2oTD
s6dpvyzMlw+p8b+pL6gvOe+KY8tIv1ejQG7JZMi/6dA6aPCgTHb70k3ie0wFRuSu
ntB6pzmdsEKu3NYaKEKcms1JMLCWIY8X6r71hPaF9PRpktqHzyRIazCSSDG6Gv+0
4CQDgpb33HihIGXdn610ZMXrCpnBJ5KKdLV9FwFtWJkczGncIJZ5tIqh5d4KhoEo
F4yo9C//ZAiNY362AbiH0i7xXCvOGKRGpOiiKtYB5Wx0YJ6Osq7xYZtvPSbJQQ+w
7KHL5tooh7Zmoy0UBKebwj125iB6pt33FosXd84lmxYu+gPvqkV23GwkCJuK+1qz
HoboFyRCEqM3Hxt9FroxorPyzmSW3ZyrkDeUJj5PXfADT2y/Jjti4W6zg2uF1x8g
xmg/kj2KuzW+quD+1b5Np9rlA5LAekeSKY49BuU7udCBfFy1Q85e+IuFJ0TyK1bM
dwIz/4FWL4u7cmlzSAnqpHO+vytTRIXp3coEoxtkgIz/c/+YvEikmnM+Mhqm3O04
4RPx79dIWBzDou5n43M+HqsRodsQuyLIu5h7/4L9x/CaZy+MnJz288DcFWmQNTki
X6dannwHolvlT5seRixrxEFDc2IJPeQDYZ/oVDtSd7iWGSuIz2RgkldMyPI31pBN
nbps+4RkVj/CZZbb59N/1HZfh+8cJU3lQKka4FD0WOHcrMOiL6ofcypMu14QbVGS
OPJ7n5/NsFpZ2DR9IXfgvDylDG6eycy+duCbsugVAIHu/FxdTCBWQJlAEUkMbMsW
o3hY8of9Rchg0vrycDT5hrWP6ZlEw0ZbKXzy0ixPOt3+eMAoZABXmkrs+vEy0lXG
WScouRSU5FTiEkXsy6XCxs6wcAA5sQ3eYpCl/IQSuGbKM/GmMTKdVIq9y0EBqH8y
twfdQSyb99MvMopzEaxip02rwMQTXqrUjqUAWbjp3TrNEaYw0rbaItg1T2CapwUK
6jcnu0XlM+uiiRC1btKrJ0CrYHm5j8HUy+poetIx8s4eN0v87urfwyjxVmEFktRO
031Uy4gixr0BL4PQjfxW3Lsi0qI6oJJQuNOZEUSssqdTF0uIPNrk0Ekepf68+dQV
phMQ+Pno/fC0lbrF1g7A65o60WNqxmwa2Fg20Y/FVdCtg99LCp3YIX5ZOxDbJHUb
RkEPnbQvewSamrxR/48XoabWt/i49oi5L+6YG8T3z64N3lwQRrdt9UPYVjzl3tUq
gPX9BfZxUB4HWp3tvtQf4rRnfLCJMxp/wym4yVLt9+kb/eCxtQauRh70NxtGCKMe
FcwZ2XeQkq3YptajivMQ75UQXc00YEkHPinG2K4ihJCjXawrKiXAXfkKsu/HHP0N
KBOaAKeUiFMwBxikcDAioz3LxzdIZqXSr0OsjBFDn+HUMYooXFMLGLPusjYsqCJa
N7diqCjA7FEscs13cNiPSJxPJawE/1RXXBahZVdJNCRzlAhMA2tYqctNDXVX3bk/
LyYxdzgXyvHRrgBg92R7WDxED00zs/zZhi8UDxR1r8Zwh+uVa377jWsKWS6EF5p5
uFonMCYk55hL0p4DPoUSwNJ6IfKP9A6TH8G2RJczatEstc491EiRXA2q2tjjKKKe
Kva5mQNg+6MrvI6kK2OUBz4Acf59or7VRYGYV3tn1G2RVV72mPryjJbWAU5fHVP5
Jb3I+ScMPxUqM20Xa0K0bNDLcswkBFUf9zagoWQaIBcm1z+uRlmc1OUET/MT6grA
QBYoND47mvC5+VPayCVF9QH7Q9vEzfLjy2WbBIKbsOt2iKtwAim82WUG1CWMLzzQ
qJLmiffN8e7TOFHc5Seok4QHAuvzi7cOywha6Y99qvyw8maT/FXEv6akDw5EiYs0
gSipwwx0XY8g1y/3dyhyKJduSodldrUJ5CxXsw277PtgFS8LB5kd4z48Jwh/9CVX
sh0nECqscDdoTyQ4b7rBndTQLLZDP2EGtTnYLHK3uufxop2Wl9S9RAhRA8S5S3xJ
nkBalFT+/sgvpsXxY/4eN5RzySW4tGNXqOuFuzar8nVnMVMCxUZGYzH439qdDd6G
SBUXWRe6l6oMrlrpas1LGdT/WLd7/tvx6EtDtFFXfJMz4D87WYzj8IegCNgKN0W6
/EjfaW9kIYP0SnRFS4qFmxeLdbPSjn+881RWoY4YvvjGNToYWRYhOKCYdZNG8MXM
WJBaxnWfykrnI3VJYUBeXKjliP4IIwvi/HyFoGNZRhQQFOsgOShOsntVC1NfSbV6
HQJBGz+pT6omZ+VAdJjEeFTheMSKVxoMJpOiihrEKSdpKSoBurbfCa6dRfVbs8j3
DFN1yRr7G8u22+2IS1Q6Sehyb69yFQMg0H2OGohBuZj3sX2KKUMoPjnZcIgRlRY5
0Mq6teBIom2pOUwjIvpfRdlc8jsr//gWO80rB8Io/IdiME93qr1n0mvYYYcWXbsv
LsaW039qUD1p7RKnDdqPqn7i7bHcH3n3dNz3XaVp3Skyg0eWu5XremtFsYL55oGg
uTPbdJu5/Q8U1Y1Js0xCHK1+WZiC+6tfXTCylVITrQnZi5LNSfziwstBRSYaH96+
HN/fwiUpIWgi+XbBKJII7VLBfH0x29TLRPGsLwS3wpqapHXh2RUpDOwTynIuzDk3
Mwd7iZjlQ7ycwBFSseRp+mCyhyy0ijyghCMYfiNpxnFMA20V0rwTe1tgFJ7MX+Ma
tBuwY+LW2J3EbJD+Mqsi/zb8QnuGABRjMJZi6+ByJSz8APbVh2vV9JBHzRBgSo2S
dS7Ary8k9Bx5dvkraE2lFw+/Euhb1Q2P3C8gkrieBU5gvP4qNikYFwdRpPzJS+bl
SIQxqdojiMbt6P8vnLKJpbb2ErBhjAlfRqhx4S0hOvDswbrBNIEh5On+0gRUB4dO
VqQp6OfnqNVYM/x19Gd3zgN2zuSKrZxLYBKHgVLaipFGokfkETijyUtL9cfClicl
uHlDuIMi+wrFJ27QqQCF5qPOSzST+csDRBUAqX2+RN2j7EIXwW/bYCJpN1CCf5ua
be+oM7PrptvaxJHcS5dKH1ZOLsiifBci33dtZwfTS43VlK/Id9TvgPrL47KzU3vv
dXNNk2FilxP6FRLbwBpPhhi5jjLyyyzfKfJ6sasjaUmLrSGtuS0xfscy88xfCje6
+7mTBR52D9M48YMHa7TREgnHA1VZ2BYUCfu4viQhNS6KIrnXT90QhivFoUVSJ642
hw+HC2Zc+SPTNb5DVC83MA00IvnIBueEBd8iN1U1avGygNJ6MYeDjcEjYWPchpJB
A0+g59saJIVflmguUDwrhqwoWO1xD9Q7LmqC05xrTgD4z/hVy88peKBF1977Qxd2
eRotG/OeQRkKtCj+kSi5tvQS2Wrhm4aESAt9fu+RK8+uC+oFdfiC9l0imjb8bvcl
Pktxf6cIuL895655k8qJCnJoGPZRvUB1isTO2DMgt6LzS52paGxt53bnTDMGVD8D
xFB+8KN4hwlVGlSE5qsaYnj5B6rv/qD/EKtbyR8moDWu+c2p7rpAC331DuonOl4o
3Xs7q9811/lSNKGEwCslYJM892fq9yyV+E5/KP5Z5/QfEkCOtSJlFqoapLexwrWu
cmYwkhdGKe3+eb93YRTUYS3D1YbzcEPGx9q0e6WE1MmOC9JNCs0BYnURuvZ1y+zX
9q8dYxIzcCgY8Pvr8v70eQIlOLNzgv2JkB4rujTpfHHZw7M6FdBfm6YvYOAPo6pY
sOiJGXOyQHzF85ccSuHrKAxJtChChe4ItjTk317I+VGgldrFJdL11KomqTuY7iDS
9nIB4GT3woPpl9n9GcgLPWR4t32MRoB16eheq9cCwICnpgQMd2W2Sti2ZAZRi8to
Eo1Qj7cXTAla+HCh1a3FPph4VzixteRLSLbJU+KGha8h/PLdClC9EStJUNBNlbPZ
Z48wjRMeoG7mplkP2WOasTFtzPTsCqJlr0N1OQxv/GGXP5VosdNImOK+iJSFOXlT
ZGXoasq40PoBIoDbHl/1dTUAJofkBNHHprVqHNYvqNEPciTqaSrS6LD+lo/c6T8+
lPXUnXa5OAgZ2StNHi+OcpVuwzqTt51qQ+FrydwswVaJhvmORoKxQwuvVO47Z6Mj
V935Ah1yeuZg2Z4TSt4yo5FHpOnM9cS1dsDIfRybomW/N6N8eqQ1mWXtI3EmisM1
T2bnAvLMYjWaKuJ2bn4A7t5B//CTp259bFJ3fvsFTbRQTTornR9LwUuw9k2GeKv2
SnTbFLjMZ2cM7AtDBRIcyewnJW5xDmO7VMdsPSI5kguvvrpfwliAimQwlgMW+7d/
On7a3XYsIlsA5wmUz0g6T89ZA2z89MN1ae91606TtKFbuzVJHZ58F11Xv4jnKzjY
5bt4lysAn9F3HiCPrV+uAQ+O+h0cigbJaZamkrcpx6oVfS2gRQMj4zEWazTncHjk
T978/fQJGtCx4XFoE/edyInM0TF/JL9sxE7rk1ne2fkd3Lf/8cnw5XOhbIZyvUj0
H0MUwbut2K/qFdrfBDXus9yUMlqiJ2ZDIBVUbgaXm+jLcQBgsYBNWGWth6yzMDQZ
BCv5EKyVplm4aTfRKU4ST9JZkwRWuNLRD715lG9yXhYfjNfiYrOtdWLdosnISJsY
nqdryDLjgmp8ksUmqLtYsDYHiCObg0hzuk54hoKlqsWzG4nSCCXLX6r//3lSp3Pj
Tbt6O0YTj3ke/o6KR9Qy/DNcwpmRfc8dyS6ndpdN2A54WPpzNSeHeG/KASw3np2k
DWeRVRbPlq+sZTree/hgbn49lu54pfOe4DU8CC9T3vsOuVBb2Uv31Rd+he6KbFUa
hA8+WZ/8deHm5OFOuthxCKCuv6RD8CfGPzAVgaH9x4csKeg0oJR7dC2Fxxch3Xim
T6GDaKpJim/r2yGuCrS7hZ/9kyAKxC5HD35qEvg7FzvYmEWgpPrZcEut4YPC9uhv
MfPcyB3OBcFk9teP1anwXkxKRxO/n+CP39v6yhuvpBfrNgz5LcFPiDs0h0VK//3s
B1SsWA8HReqSnBgg3uxDhC/0yH5fw2ok/9BF0XQJCLYnwOJnh+rO8zaHxtTlTc8y
6bhGBQWb2cvDNObQJBAWm6P83d6vYr+t36v1ZoM4tBqv15bdJyJgOTxCJ2hXGWFJ
ZSWwEGuzIvTu5Z5p3c99crNn21+0Nsg+z4Q0bmQQRks2B66pW0r/JoeVGhUFZsM2
PdaaQnJjrQQT3RiQm94Za76OTQQ75aJLcwJufo2VFEQIOPQCtMdKoTnj4Nx3If31
4cY5vpwbXF9icItbAIs9UEc22wDHRRiOjOaW0BJYAgv0mTDpuL1VanE63RdtRvcI
S9/R7HRR5XJIBNkn8dshtYOabOAWOljWNhyBHU0E0tZKGGtVfOcyYtcNB/2YXv5t
yzUF53atfVYlx6EYZGTSnxNeiglmlhyl+NL/Cu9wsyCCEIOvc1BBWtdbis56wHZt
YW5bMJeRqi320iPNGMJ5W+mAXDBZALQwYxL7uMXYkaa2yaRIqUAR2TT0QpS1Klt9
v8zyw+gH3CDPW8ZZRFJJgSQPuvQQW3O/IoxwDZr3ypEJPAvZ7WJGSuKtmP6akQBq
UM91MXPBiuvNe/uJxpRN5P+F2aCc+JH0VzOAxBDKNXVfQwdzF48Qg2DhlznPkZyF
DvaRptqcgxUseLMb3aM4ASs4jeOUW9Rm52LXIdysSmSrh0mNWGEeIiR5LWd7i7wh
w0Hae4Pgb5H8WhbRm3Q9fstKcdFzXFpEtUGMAYmN1YDQmhKmd2PhMe+YUTOKdxLK
SICA3C4q4VQlRY71MWnEovI8okD6cquEaaspl4i0KUXSCC53e8EWWI1E1xTM/dSc
rF4kCLr/A4MPJPfSLkCConWMXDN8wWVzYQwBIl+gYzrzgqA8/QEOf/YjJxLmepmF
Y1pIfuM38WICZ0DqTMfpRZRQqAQ5FtaDeiIuqjsKodPe0y/rXMQ1ypXSsO+c8dgu
aFFpuiwblY4TRszdTdKUkHxasI46hDeP9NfICSbHOlQAxvh6ETEoCdjUbOn15jAT
rJ52a0HN0kcOnBe7p4ShMh2MhuwShxmS5CmM7DOCLV1Gzd/UREKdXWVHbxBhtpZJ
/IeUTk9jpvpQLPxk9PZaH5TdnHQFZT2KoCPAIjrzzePM6QoTu6CH+5nbNDcfIhlj
UmKtzz09ZSrwXDim8jNyrlN4U1ArFW5MSBCcsIJitDySAlVS+j81MNSe0oaqYTRy
T0YEsQDsa6/Jx+5IdelUXEYyAhgzoh7ZXfV3Y0UWJa0DljMfh2rO5dY91b8akkgS
faNi/ng8/Jxb1oJJr6Q3GroMivh74amTWB/Ut+7obTn38jrRcT08koZLyzpqAN57
cnmiVyZhPZdxpJjyNT1mmyrAamj18awS66bhF0GVAC+lxdWS9a8GS7d90mGHpsq9
Q+3oFnIiajdvmeJZFzoHIBZaEGIPezYcZ0GZvhou3ouxvSPJL4FpXWQYIkiUdc1Q
Q3GOKXiUSZQ3QyoWHphRIe2ffxwxjq/UjpRQd8+geaC17Ac2JEtu9wGLnNvILEf7
uCeRApdiq/yXTByLWRoIAP/YZNU5f7PkK8+imAKfGIdEeK7lRbXZHm6HZmfWQAvS
Bbd74JIPZqRflFkVIU3mT0QTeZS76Zi9hGAvf0QgSBVny5p3miS2iKDvBbawEfAI
8qNJOLmsHYUM32OGQTejaBHIRIgLJrdXIk8lUJb3y97hK84JcrZdHsqi1fgPcKql
JeUc3WNyEISFRw8I9j5nhBz3yOBlP1kvDPsNAIyE4Shqzdru3sLwYMe3vsrLM5gg
ODD2cOgW8mnBVJu3PeaAvF/sslkGGrYYCC+aAzkTzQNkpllfVUk2pXMHXHoKDUUv
nyw4mnR6J3fnWZHv9CIY67BHGGf6tqmpfplnAvdfS+qy7aqBaT6UsFhkgqaEyNzv
1GEPYIW+KPeN1twvtDjtBh++rEcp6OExKMVvFhq8zEFj0oKQX6tlY4ujeTVrM3jq
YtGkjWjJRb73CTOuDWwuYXtwI0xq8HKupSF2mWIPUvJuwQBC3vRVJ/Sj+lgUySAr
tP039vs3Dd71Xjc9la+Twb31VbB+70DaJtrajZN5QmpxID3uIPlyvn1XokRzxna2
JRNIl5+iZfH97UVL/yDVu2q5d2ICYjuKyR+czKdsa7XrdkJP0b6LJXOME5sF8MWw
pRjYmvskzWDahjMkfRcESyV5ylkWOODfvoBicHe8nfZu0cPWrkVfdAg5h/oFlNGd
GXYe6er2CjocqDEPqdMT44iRGfQPAhmg1XXUreZ1FnYkqRpNSs0AaF79ujGY5k0o
zeqOATjyBuR3XZHJnXKn0WNNpWR0kpgkLTfuGz8GrFCz5t6hSvsq6Y1kwqSqcXiu
ZIuo2QbooSxn8xu/esIEhhfma6VnBpqOPYzrkcMOriI8nhIsLWHcVfmivU7W/bDJ
OQTv/KYo9rjBhVW3vI8vG2u7vdFUtldY35PrnSRdC9di4DZomDZkEB/7GsoAz7ed
7erYvlN/lszjkKH3Ys1BcUb2vqOn/l6tZ6AQwPgc+viEazU3AKswslnwrxxG/oVV
Pz/m+2UOMjJYjEJ7eBdZgf6djZZ4jSbO/jnrYZI+ZghndiWFsJBM3th/X4L7fxLk
91iCPzNJ9wQWUxk7CtOUKYDHc3eIXVe54v839/Z/XRYy4tId0P5ZUAixj42Yfm4o
OCjT/3xUy+7DyXdhermx8ir115Vv7TI8JmlKZH6Gm2HaufbTve78WAAp2MrBBo4I
AfXD3xLGjgADAesGRc0D0GLq4D5aZPoHP7aMyyBalNAaKm0bRg7nIKsyJiJ3pbeq
5ki97zKtW73cDjZhOaFzgpRfLftJFTReSa+EAD5u5SaUgCP8AcFVz11cpCBDVoRK
5EH97Q4+vun87OsnwHrRbNkiTri3jklf6DlY3d8Rt2XjpSllGOznHSSp4a9thzIK
aXeuFEFFsEYVkMq2kSD6McA+a24cU63Xcwgyrh3BCg7tOoeGPVhyZdmrLg9fH8DA
Eszw6zAhAaet7G+U7ZWK0wb/c7ym+3lFZYyjzNZQq5aS0+qqd2sXBxVOstUVGV7u
eYSYvAgWm4zJXUYeSeQ+SvAuLLZCmsbFcuw5umPxIuYIjYI1SJFVGm4G9kBSX8Ys
GMNge8wkHDIRe+mOBYYSb0BUyyf8YFPRDQ72WixNDGRGW3+9LetiwA20fSQL0nIe
kkOYzMUZXXnH3HCkS835tbh3JWIZdpAJVoJs50Q//PX3z/JiSTSI80KojpzRAhm4
z9XyTDrzTzFKO+UtVRHKqpJENvfG0Lrf630ED9ZoJ9NQxTMdOEQcnTR3gtUytme7
YjVVHZ4VTLejAtemhs1XqVGdKb87gueXDAK/lrM9tNxzx/gBSGZORrkmpprN/eOL
u1+gYRKCX+O1i98+Fzdb26GC30+Efc+TeAnhLYPJBdGhnce0lxc4mluBGvr0ud6b
bQrypsBWroL6YNmFivj35ApF6lG5uTRnGZLGx7I9u1Hg0z/HhM0ez4LMIh8GSDjd
SZ9ei08OERGPT4xHd/SeOXQQAawSQ8ELOdd3IGKPuVYOZbhT3WwEBRYWxbv8cMR/
jZf4IKiMSRNhvQBC7Vh1mTzIAvrOJ8nUBxQ7Rb3s+2O+Lkmy0pCItw7nzuWBVk+6
4tt2eJldCR7VBI8zgONxoSMJZqKw9Hi4uYABhZbkTwg0+d99JFRkAYNidAcKXSne
PIf38TeoWYznsDVyx93b05vAPOJhre6gEbuvpriOvf7yTwUedlBur6LMGJ6Kabm5
rC83Jf504uOUeHumuQqQZo4DWzoiSxIFG8XnSh945V/NghtcG6E9/5bLWZwTGM6Y
wQicc4EUwQs72ChayAqsQRQ15qpAFvT0Nk58gyuAbT0Hrx3sW4hH5pBUOjN+pTC4
h9G6wUp9sZ5J2cChfI2a/zvFTcLWPj7vhiFWT1dztTUB5yUzF/FKAQxF/5bt5ywB
oq4k8mKaEFQm1qiLGm80bI6NxfLFwC0NArdHK21cbgXQGqeebaTI5t3g1Dp0PtlX
4Js+c0E96dQV3HtJhQqLK0/X0LCQFEbuiv/+keB5mFc6G+WMNrITckz1gkB39Si5
o9K1ID2zmxBz1nMnX/aOClq0tQxpVBO90Jg43xxb6NgAf4C6o9w4xzBevlo28cAL
UKlpZp2pU30t1AF5c2KssNs4F8u/GSx+LlKwLD/hw74TjBmwj9+u/vA9/YfbV9nH
IzdTHUWjogBx9es38ZWKEPqsnnSmtLDsvqNE9i0AoyYypRT/j2GfiHv5upGmImiS
xA4B1LwzCCrlNq6GXuZVhCzc9rJWoIetONHh6Q0joYpCs3rVD+gCly6MRtxNm121
16Svg7ucQZvw6cvtaL9hIs+FR/Q9fueOJlKgU31GBigMCUpFz46Syet9Wqo6SFB1
pUXutQrLZQRou5/bnJGrbywJIiPfIrrs5urWNW1qnGx1Zg0z+vatxispKd8FEWPN
iAKoi2BzLipdHTT+wQ+4hypKyzD97YKbdgFdvjuXU0vFdWxnl12ELjIIRxtt0CJD
DxCTmv13KovReqvKs0zk6isRscnhOIHq/tRPozLRLfP8PvTvwNPro4hp7YA1jpXN
HyWTb0h5mrnnhp0IZd25c0yrvesfJgN71NKbtnBf6xou/Fjy6OC6DZ4aF4SZ/ajr
6tdCG9QpPtj5+NpBfpFWKPvLz+wUfj09yCa3IEjbGyFE8ZEq+l3kpPuMzbGIXupb
GgdeOgkVUrspWjL8nifM4BIHPN3b0CMOuIpAn87O0XJXoWWL61iw4RAY9GiMXyFj
JSlviA1AlNbmAbf1y6QWiSbZwQJCzbDWIPb4eKtACxZ4YtSR1txhtVAANqBPhtAP
LHQx6iYFynnNtc7JVzYkjCDDICYM+6AhtAaHWLRZNTgnIwTUL8f+oplq2esTXbAC
AWgNAuPAVcNq59G6FOvSrOuGAzhRggXlDFkBCv/9cZlhe5DAclC6iG5aVAxSuDje
c45AtHsyPQYZ75t7d7maY6zYGDDh3CYK3/UfpzZM/XVURNp8WetNuuSEPzdtif27
SFtgJzXhXkPLdHXCe04JTUJlUWy2xGse0+x3MhdvkEgdgW6sC5G1sJIOLNm4uMny
SRA5SQi4fXfcTFrNyVdDdnULwY/1hJA9MPfR5saBHnL3bi0dswo6b/UuDsMa+k8/
+EWwudg0518FTaJL6JI8k874YlbtADDwwpqOzEAv+6PjgBnqyRpaLk5Tx8ElcQ/f
sjgJtMthutsqQ9Z/y9TPEXSVXWSpzP/8jl70Kf7Jkj1ow+NFbuTZoHSC4qr0hwKX
gALadwlzf3UnGS5xmYEoCA5wh1Sb1l/qCxT00219K/8zAfEhItHwb9FzG0AyYHkg
x0AAbDgQdl7Ujo00QMMvKXkfv2D2Q/wgnzCr9h5YBp5BRL7um90zxEwOcIUOI4lf
LqA8TKVKwmJ+O05hdn7VZHY1TIkzNaOuubaM2K0hrBl/Z5HFAFa/FB1srUaH81M2
xWZBDi7SlZDhqZz7P6KdomVsyvOjMs9awlV/2C213VfgIK/PvhAJlYqABteoQ5YA
OUwcm5K2529mDj9f4qWM8JoeqMn7lcaqe64/PemrkIH7rGGKxZ77/YM10+iyzNOw
BcqqPaKTiQsKXvrXfqErPlTlTWN7OrNS8tp3jexuZlUbV6soOd+ArydCqWFftV6B
Ge3aF+KAOw/ZUYZApdkdb72aCulLFD5tc/k5V52ufWaQkv0I3fqs8s238eRc2MtW
7D9J3P/FK690f12pLDBv/F6NegK9fjMdQoC+oMIH6XiFVoMqvNSAA7626qgQXsyy
g8PDXVuK6jE5e5sh0ZzKIY7iIbN1d5pQnOandQfe7CV7I7KYrWPrE8AkAbhh/VrS
atjAn5N/wYjaFMAqrxdM4Qi71btltCup7N+czO7DnDObUjf5aZojgZ1OpmUt9ZXT
JGD8hMrpKfxLJ33yC2bexdnl3C69nLaBAS8GU2rEdhVR2Jf/GrhLA4xsSMIbawF9
VXg6hlcmPObZAVU/kw2WnkonHOuXUarIV/ZNmb2gyuKiMCKfGFR72gDWM2ikeYxZ
78/5PIr5J7dIgGfKGzNM6JGDLpb3iuKS+lGoLIWB6RB2jeJwPaW5A3Bag9dZ6KQ3
bIaURrAC973g0hupfzn8pfdH1lsV5vlb21sNh0m92Q434P++clRawUq0wwB1f8x7
s3yWB9Q9kZ3AdvTJX3lWylisDF3v7h3+RsMKcJhuE3hT5jKip8n3ribZ6nfeknJQ
DmIzIG0P3CvCyhxz90X1weh4RSgx8itkWJm6VWMun0NeCH3KGIg3wqDntkBCp5ts
QNkZkGq7Vxj8l8CfIMnijxMhKJisCS/RLHmGdU/LGGp0D5gNSW8dwx5kSl+5rHnD
FxfzhwA6xhVxB5Mx3DM6ZVNmtNevsgwYN/o8SBF79vIjnLKaobUgJ1vFvFXgbjOi
sVfwlr3qy3K/u4t7+iJXWsqmGHQwNZgTJNYbf6MZCLyizU8HEx8qUvAWYr80nw7E
5jqge17VnaOu1kRjNnMf6lho5SoDberyS71b0OJRVJk35NGfCZBm4+c4tGXEKJgp
x1KQX+EQP/zFAwAeDONrBNtaC+DLQ8NLgjKmCsuy0H3/cvuNx3brzDRCppKP+T/p
/3f6ICK04lnzgzVR/NJvh6Edeo1J5iquvmwhjMG11ue+uKlaQb0iefuKTeTyMEZR
ItjKggAFk6tY1ICxtWeRaovpXaC3UN+9oTpPrVvPItr0bxUFlghD5v8VFxwSISV2
Fm3HbrQtuUfb9mV54gnafRh+PCRrsEoctnUCyr6qAL6O3o5u98zza/zQHZMVZ0lx
qts1SGUHEtc0S7Vteroc8jlpfcNA7jYtMuHOuTT/SGJS2qosveVZZyqHKBkqKq7C
PKEDsixmDmFdxyBXEaWFszVsGqjQ66cCjXNXngHNJB7rowQEiksIb53gkHLQJf5a
lC1epdlPgCLLXH5IgLZZg68OzR3/u9tNFRk+gj6VEXRQQAh7AXMY7cbinuHL9SUb
5G2qLaR3v17kY2ZrSqHZEyHhZZU47V9Y6QeUght+7lg195+g23Q1c4bVIV2MtDzU
qjYXDF2Ddz8KplZ8tXmye8AZT2U3MwMCu7q71bzn3vR6DBmztmcGNgGgSGeARFSc
ntzisuRho/qhqSd7RTSHmzWVHc8l4gh9s63dpRVLvzmz/y9Ou3HyQW6Ar9znkp4p
WDPej/0DwVhlV7EmYr//b47Dbue+ILCg/HXr5F7Do6DRvkMuS7CHAk+VPOERuwmr
IDHqIka9MAxCxzm36DIZJ4abxmnYU/Y26562txMLhPV3EUWqFplHvGe5EONgwMWp
oMhohlbt1UtKFD5O90IALTBz4Obyc0xfunffo12uRVVzCGr8AH18cdUQcBrnZl0d
NaW9Yhe7JAvVxOZ8WwCWVFvkxEB/XvBwq//A1ToCdqRqZpW8okZcm0Aec7wE3h/+
kxcB4hHmj9iztFrlfr3qACn5SixtvVi3ZDY19/phubfKYRYw7vrziyCdoIOqO+Xv
ynM5fEKZ/ODaG6MF53EfnTcba0UfiBr10Ic70Z7HhTBBhispg1NYG7ho2Xm//x3t
9PW8fm+RBMAfTQ2ka4Hq0MZTXIfo6SCakJKLVSzO43RmkQotWwGw1B7Ey4zqDyMs
PX+rWVNA6vDCmO6F12mOj1SroHZflMmB7jic1A/EytcdSfR+FTdAgFy7Iie4WV/J
imEZsdqD3HPktaFvBQcXXgwxdoPI/GRh33PFjfmqEgJpKfk3R+2lsUr1pZuBuiaX
8HZ1/8j4k65JkjeSF8ujOGULMoqJ7kxGa55YdDDxIfnn2nJnfvTI3P9XTuWZL9Nr
nbG+dv8NJIE06Xo6Ek485Lj7NkQmlpB9lx4XETKd8Cyr1dzWLSzike3T7Pl7TddM
wSc8jYMmzChaVY7O+QDrj+Yzf0XxnF6A7dvrMu7MYV+ant9HAPUGjUhJyzjl1tBh
QOAbsLdk4U6mUYFUtHuTy9jD5oL4OqlnHz1sW19RBlfWvbBvmWCFXZCXjx4iI4Qg
6gDPZslI3DFXpuzGEsbkJtZr7Mn0kdGWLDVcQshZJJSuys09UDAusu25ei8g+rmp
uj8NmmX7n0ZTwxIPIRHfRUmKXrMy7MGblN5nMr1kEtiorkYDkTS32wgtfq4Jm/rK
l2HeHvtJEDVPQbKCvQsmM56yJctNuEFCaLXnvItdY/dN9DG0nfr8FyiT8rY7jWhp
TEuazUUKaXjfpX4aUC55FX44aAjkK+gcexFaxgSjjp+venUrZma46WZeX59Qb4sF
sZKTxp9Tbko+o2Oif04RYlmKSdwa1heYUcj4+O3fosXO1FFvg8y7hpgdZGu2cd2z
j66YeO/g8zfBBDZE0+8WncnCkUPGBJ3Zd15OALUf8Fy1eO/WWD9h8GALGUcbc83z
6KkAcx8T/X3EX0anmuGbST433WhqmbjPeSPFzgvfG9vNCd9QwEDumcGXNT4dmmnW
UsQvqScgkWCVqUPvlq0fM8B2yjr+THFUQq71s2BnY1QOTvJkfKWmA1f2IBQUh5Fk
VuDkGYgpv+au1ZY/ACXc4JR2r8OVRnVKZLd0QSDQG5D4xP5eMfRr0NDYA/5TRekE
hjmr5Wy6Ss0nNtwtt8dzImsmL9ZphNqhiGxFd3pcYL4bOfweTHNQB+56hWaNQ0pq
rLkqxuPFoJxKBATu/3WC++o1ByjlgdQ0HAAS/LGAOgbZigOLwmxwQkwe1eVPMQFr
HFoYF1hc8ZVo4SkJ5Z0kCmUoTtglBSKJNp2FrJ2CISEy+3tdCkziKxUYYSkbBNNf
FsO27R5/lNCef/QFycZPApqi9x8vwVd86jP4SPOontLfHrlYXnrccljT2SK1YBZf
aJkGcCaSQ5RlQmwkbLTxI0C9JlMekyPHE2Gu/4oBFckbjeSjt30WhpDkzQIQCIGS
UA+WU3YZXMl38Pi7/QPVoFWYgInhN9id35L/42fQlcNMwns7ZDhKhqFitbWtdCmX
7VZSGpJ9DxAUVkR92qUrcgxY6BzI+yYd+BqFxJhd68PWnHGua78gwfRx/uVT4xy7
/uc7cYJ/KG3UWAXtmDBXPER8RJlfPHeg8SxipTM7bhAiYIRtjNFOhfTyRnuyFGLR
k4Woln/7bqbdxTbfdgeashbVfNNbc7AN167iXnLBIxYt0OTmwE0jDVIcnO8l9rYE
6b+GIVK5auBcNpndZOEextTph1HUNsRtsbJM6ePfrLXXv3jBOIfWs8wjAL7BLxC2
ffZBEafoBPVP1J54xjJMXhVtSDOJYgNlXl6MVH0T+CDYmktEawkaMpDHGxlJPi7o
KanIroPduvSCFv3K8QhGtLMb3DqhnPuMKvdNk9r2biOrPLG0LOdBMRqJYCSlQ1Sm
72Xacr5ACX2RG2oIfbFgXCIEmzVHTaPQKB57rye4BNM96Ej4Ov9U1DoxH+GFZf8/
tZH2q8WhnJQuOIE3vIUQnBBmYjmVMwBVMq/WHVL1+ESXpCKIpAkGD54ZyM3crLw6
3ouTKDshzCMgmKi1u+eCP4OLjwTUtuJnU+OGqlWc0PqXoFKc9y26hU58zGPvfpMl
XdcY9hdCN2+Q0xr61RelKMyX+2PHMMAL2Lc1ry8DBhR7CZeY7a7a32ub4EuCytQO
t/kcjH2rUGujxXvkXB942DO0tx6NLzdaLHpsdEYsl49WHNgYGtjNkiNBQ9Iac3od
3wWkVXRPm8zfefMygbXLlVbKCHEwJ+mYF+5QcYSwdP2h9TiW9dpFvmwEYa8lpS2D
8gGFac3z7tkNQRa+GReQap3J6BLGmODWZDAMoLHD+WT5mSZozOPtifOoYEr0z9Dv
db7vKFwhTOI9hUNNHojsmk/xsrQGhopqca89GrecaadmT70AooGbvC16BC9V7FfA
76iTLylojSkKk3QyqtcRoNfYtieqCiAHG/jOGgaHGtac/y21CYdzvKUA3VPvGAFJ
zjl1SPZlbQvbI1QgHRXY172bzbDWkT6YmGT/s7ADm0Ai1ixsc4zRpEDbH+jdArDV
iDkcxr+423Lh0tIT/Ps0Elh39HMXl6ijx2tK2PyjquhbD9UYj6K5R+eI58FWc3KW
j28KroqdOaNrmry5wfgeZk+7Plyxu7yoDAY8JpY3mjVGKtdgcbWE+CD4smkHiBOq
4c30tGNBgrE8KM1w7DoULCRm2BrwaRO1jZrUeKTBMQ2P7gLynTBKQyU6fWiJH8NN
1Pv3vYn0eVoN1mji1mkM5PFI9mq6ESYJTGInUQstanH/XvB8rcw74j9uU+usMwkv
yfWk2QlhIc9nXjdy7kPp3U52+OfMqPUIkFiJx7NFzbyNPuR+eV4IToYZ3qQlm7tW
hQaKKYp2xwHQGTFdarlJtlADi0aRJiBGI343OJAaiVHGSqF0iPpIGbDHicdm+XFq
kuKH+teKGTTxM07XVy20xZZ2Eu2bWVzjFJR0kaVjLKtVeyz9rBBLtoji5ETXlJM4
WO9JEiOzAKKf2/qPGirQCxD/qS7b7SHGct0pYcgxzjseo5cVfhW3wOHVoZSFT4Vz
1E9pdTAnjVxqaBqWgUiVma2ptIHV4usbPvOCGnjOnxFVeViJE3faKUsjy5Qxu19W
UwHyiv0GtXWAvnLoW+3u8AdZuxa+a4/o327QD/wmsAiITSNUQg10JRMUWm8fb5up
TS0eeyA45XGDO0Lwvgy6yjPO77e5AsYCwLOiy3BhlUcfuPkO24/6QljGh4EwYt6f
JqTxzIXGowrRdLVZB9I05qukm3p98SriIhMdSaZbOsRIXzfYbgcMljHBt9wbZCib
Te1JYysXLLyA1DRXYGyIKY++TAPZWNBPC4nmCAR5nR2YaUrkA6WOop+mkO1eB2C2
7VS09Fm3vfvGeTMCJUyf/RtdRyjw9rMj9CUHcBrpt7Yi90xS3IEZeU+RDqrqBqtb
MNi1H8KX2z6s2l+Js0yLFnRb2ZrY9gpvv/DYPJuv86gyenpP3YkqNTHhDpT6Je2C
N8100v9o1JdAJ0jcM5JGZvfPq3+59ypgGEXWeyO28ILpGIbhCsWrDueLCV+kRhA+
PKHk28d1s75s+UGF9nXXpT1uEhO8cSz6marXylBIDrZOojJZDs02/Q6ip/D+N+ZZ
C49q+jGcYSnuyVA/PV3jkzE596SDEd7pKe2elv3iP/SWCDsL5L20tfSvtTjzd6TF
S5cbsh33t1F1o8cfiJcyX2b7mD2YsytjQDcOXxkhWHR15c7k9OV+flGSBY834Cgz
T/jgtI30W8TFT7cGFMzwEumcJrReK0gtoDY01luh0n1oTDpD91SbneSM1sWFTRKh
yqRGbUN3FfM6Y7E+3yuD4rHUHxK2xuh281rDP5HEltIzjs/SfAQcp82VPpX7JzOf
iIEjOrQGX85I1ncLTN50DXCOKr+bKhSmSAl7WhU8KJEADnX6gw7a95Pu/Zr7gS4N
f/D3VqEhyUPXNIuXWdfhDTkmGdSoGcgclekf76B6+2bPY21t+rVX/le/QP2OKWdR
ghZMmIKdPIttyc68tF6pIQvqdH/Z8Ntgk2O47JJ1dh/14ya4c4zm4vOd2YCO5baY
BRpFPWo4mlU0OwVrFBIzmT8a2CIuC8sxhk+xbgJEkUOBahx/xDxnajY7rFAvllVu
J67ETWBcjuGzbfxXqVbiD3BlbCekrQ4yQus7RUmMfYzcDtuni4QzBoa6rZ8ylE+S
30gU9iklpW4aDSUkpdmN0E5MfIykBBygMlCgAp+XBPz8Eg6FN3a9xnPU9xBnB0A/
AVLPc7HfS0bBlDgvJcc18gyoBbjPaFS6LkRoPcnSigDwG+rgUsEyjTD7L4cfd8ej
kmn+3+JHXy2vnoBwqewrJ8yW1/DkzEAH1xUFz/4ry3kVL/mExTJGIDBJeBU61qd7
BOHbg9pO1wV+U7z6YdFdzWPldFYrmNvrLlbS5jRl9gTzxiqIJ50ynJdPE9AfzBR7
h9IOaBmDfHFre9ZKoKY0wYaVJ8yLAcoNxtcX02zGMHzpo6Yt2hwgfrLHVTd34MEC
d2zRLrQFJNL4P+EE92Xm/CjYK7x4Xng4OJ7qTujwF42W0Y54j9TgDpfQ5obnFkJO
dOgZMF2L9p2B7cyr7m9jBppDJDHs7AsSjtZpG/GESp315WUO10E3LcOn5silUTxo
lyE3tjrLSv/Jx+3Kfrbp8G+tVQR4gYbBC431G4pn0Ju1aDNyQ/4Mtd4vWHpvyWzn
FSA3u8Irji91XPVUBy/ZcyFzzDlstUjHUjefdHGk7uC6h9+SBSTK/+FNq9WE1n/S
jDkJBCKkd8BF0vLF55Ug0jIaFKKSgCF424p/8sIzvKhe7nRO/5meTVgF7xZ3Nqrr
vm57aqtoPBU3ptf1A0P0h0kYBaxTy/EU8TcCnAYUZSrA9Q5MgrKUy1/7htAjVzu1
DMCjoMJ0n/reQE6cyuPLvwzqHBv79mk/skQQRuFmJYcTc2kxAsF5sl8J93IdqBw5
jLLDrT7wFTrN+xoWZpXRmyrZr6GubYYgk6PggyQaDVvbqMtG28WawQv0JRWM/Z4A
A+lZS4iK8K0NRhYT3X9JVfHkeL9zxyrnIwzh+0jmDH5aKh2rNvkGNLSezw7eXPDN
encNDhLRb5k8PlbZmtpNu0hofeOppiXcA00rVc4eZ7TkDq/m34Uvguwphb9CUnsC
JKLk4lYkXWRKr++60cWQIyZygauRn95QO1TCmNFOmw6ETuuRs2URafBJzZdHVmAr
60drm8ZAb8IUQAjXAUPym96bM4UDpM8uw6cLM5nIcY6SotZgRACM8GtOuoiun2bK
c5RukikM9NipYp8J22DwJV2/Tyylsoi80goA/HMe13QNVzb6K7MsudiP2tTD9oAS
2PhJef44BlYqSUM5+ohXqa3UElQBqU3VVBxki2cOsUXpPJoL5R3arNHAlxyWr18P
zutVsGwcv2E+kM77rCgmmEk3CsAvUeATBZ62UfEBxQ2GrA+n7C6b7hAhu7q0sAf2
t49IeugKlYFy/oVPCPFqCU3x2sZyopm7sgyL/181CvphmgohU+ydpOUDSYZhdgcU
8QOrcygz7+cfOXYnhL6/5WS0+nX1hphgyDva2L84H6oB7+6OixptXiAarXbsxFzR
1nNdJHEM3JyiWmumPVvl10I6v0AVf/oESwp+LOw7RUULUmsAMnCgjM9qM0L80asR
zH8ktRbSdWT1V2+AbMsbFHFpkuzCYQl2umtFRESuA8nrrgBpv/37dexXUmgB5JSI
ojRpF4eZUXhB5CjpOShD9bo/UqmlVV1EMlv0gJVP/JNxvrBSMS+mTj0o3erwOEz1
zAhsIaKPoDjr3XvTMtqEdCq251JcimTWeTKyEwPVCuhAbCr4IXryGYf/Hcl80u0t
BBdNzkmyGsP+QZptrybhebQNqIERgEyBdnciAu5i6Ft8fFscFXgv23+3eeoV2eH7
7bUywesysOmqbF7qPgFlHs67v1tWy6o91RBZhsuV86yeTsCR/mq16f4RuceZz5gM
tQrx9hwBzfEZhSFZzVaUHEUiaNM8ZwxCe8052H3uWrNN1ostlSboH/H5ZcDH/5KX
s0kBaROvvlNCU2DXVxG54oantCKFh4GjaW8Y4NDOQVhdacHLoBeL3q4pRcyicpEj
mJ3su9Mqa+/nRkxi00sBGl8sBvNiqc3AJB/P1rPtSgrq7Mdchdjzu+TmuwYSiOTb
PyxIznlZnUCNfm/LJGy6vHFNIapBOxYPVmKJeVOiXT+Cgztn3KEFNSN04v0rlyKz
wNJODXbbEq695NjriCaHHRRQKLgCIytccQ8qV3DaQCtOFudq2wNrezYFKYxZnCTb
Ny92gP04Z4CkvjXERPBIL7HRJgrMPEkrNO50m3aiDWVOtenec8t0kzQP91ECcJjp
fjrpYAYnFF5kGFwFf27bEPzAm1cLAqtmEXANvgjHHVeUmXUuxDayMQLKY7KIJJr6
AaGSXjCk33RB6tlEtlxCbHAZE3B0cOr30mBASF6hX8sScACRlYbFMQxZ4FMBiUd3
r9SkTh7r9806I2PuN5+K2zAmvhjmtVoy0GuHD0hx+mEhAoJ0BMma4nKxQdMZpqf9
KmdT/TmahSaF3n5yeo0E1BU1O4I+88FPlCgZEoqzkieeIBDeICEhHpLTGf83DzH7
8EgHChgHm/ycdzRK4PAr28xxZDb5+pg90SkMrmplAoWKLSmiFioJqhHCtJm/F2Gj
6e9MSLSw855G/qPhU0kBBl6QRxgju2WC/z0WRxhTdx/ctzYTYK8DC8XZ3kubl0a1
SfNXjKZp3CCmMIweFtYMgPaVdIPA7wYGRl6h3cVpja3rqW8CnH1/tNF01AQTKzMu
uvFNEg+wKxW/RLyIlX+RXTI3rqF3g6aHPwdOJEDSLbZNLep+h6aMKvLIjiRNvNB2
s9xI9j3xbTA5//02lq9c8g52zvAvSZDZ5/kOs/lpEHMRSQisFH7hx6x2cRINTM8f
C5KqShcpXWsCXdUpbb8PlFGth8ka6bYvkDgRPdVHMQXEr2tGzxbzM/Etenmmjkuy
iesPvCSbr99U5X1mRU+EyMpgtWYHdexXkceyyLKkj6Jzv2ay1LEJX7xYv8pHum9g
dzHASM/VosJmo7mfCMq2/E3s+io3nvQ3Lhc0BU0y/KSDqB9L6GT5Xt+b1I5Rf8I6
AjtWGFWbDoX8TfwvYIbuRly25K4i2k9BdO3x7FKs8Cf7LGrS76cUdEwu1XxYuvbH
KHPDzdsGzGxLsFAKTPZg/pEgoUDY2QTxynK0nvqSJ7TyGo6L/kz2ep6eQCD48+u1
2tP3AWGfTNggBIg5CPeZmh1IWndw3a9QaQxfKV5E03NcMbM/qAEpDWLjy4jUuaVs
Ym145sokWLcrYODFt/ukP2C4/ngpB6Tnpa5Bj9Hmw96S9tmOR7uOYKC2Cv7FLbjC
nHSSwK6krZdFiM52SS4OcpMJ2DEqMqZuax0jSPKJCEG1MV/epAb3dFVMHvQrCp+9
wjKHzgewqjsGsjgbpjeQQH/wwkgyPPxcywHVglXJs2U/Bv+amJ/P2f0aEw/O6ySg
IfhIZx1Tseh1/zt4OUcNMwTHGzz1Z/j3zoJfXCBOgYXZTwB8tI57e/4SoSY+LyF2
r5GnvSalp4GR6Kj85EGac54tL85jW1vwBw5TdgWM5FKpl7FaD1glwECk4tRkh7zR
jY8O4a1DWR/ng15gM0omQlTxlVgqJOIduzO4ltZeOiMf1JS5j9sCRa/p2qTmrFBp
PfspspratYblfLxQ4OVLlBLDPfOf6au40co4PT9n3Yj1m1QT4YEJiKC9LqcNtk7A
EDUEvcEC5aAPiz02MOKiQw4ew5/4f0tZuRTqCFLphl0vbh600+1qZrqPtgojxfJU
4UGYemsJdIK4Kb6eQcxvgUVS1uwl5pIM3ZX5RUZ9hnl8MGVZVef9v6Efq2cDRqYZ
BeCajt1iemJyoIIMKv0Zj+OqRq2Rp30Q2Et8AVqA2iPs5k4yxYStYNcBKHZeCT9F
iUqwg/tCM6cmqnMDbXkntVYTi9mr76GTaBqO8+j0yU1GcqLigFKIsx1I006DGL54
NCN9sw3xMYlNxa0Bw69IPiljVJ8ynFUHWvmKzTlhkoZZk6MrXQ3b+wUprTY8mD35
0edNcHrIFX4neihy7eMw3tvp9r7cldwagvsaIIL1f54fKWTtzWrXQfEqyPMYLdpL
CCLSeFK5s884uruS5Gq30Ke5mJOtrRDplZBP7lEeVyHxZ9j7oSXooIeOz5l5BTMd
z2IxFbnQk2QaMh1uKdxQ88NDXx/hGJEwOA59n3GHz/aqEy8Wl4p7d/bYEAraKS4/
uFcdNd6bWn8pJk0HgF5ZIxCTQ5VuZXLlylYjm03Rl1sUEJ9udLf9LCt0Qp77vpT4
0gSgJZInKVzYBJlhD8VYpwZRZUtKJ65sG6bVM4V3DfBgW3J5cGoGzaR3BpiNA5Mm
Kh3oaOSRR3N3lmFbk2mezcWzuqtLTDmJH82eMUc2CaFYkF7Uay5ays86KAJWlw++
BqSeNBBrrhO065ciTdB4wbunv//gQJCMXvwsZlqQkuZvWhCjAy2q2bP9t9eAKSxQ
gW3JYI4QdoecMiMxj0LA0AvH+ZvSl2WiNIpblML92KEBYMtFHQbLmoUllGD/fS4r
XhoxjUD6dHXIPcejTqaQytgVnHK/LPGGYiZm0RcZiOD9zgcW/VeT+VcHSWzHNpDa
DJsmKFk6GSnVJzHetbpGz5ox71h1TZ0c5WtS+zoTf3oaEkNunhY9iJnlD/YPBhaC
dBMcZRcBV2PoLy+6qIszgv2Ew08NvxF7SOgW8vh749kcqZPI3NE2M3cGFkX38+qa
fZa0eJ8tMU9+7rdEshjauMX8St7/+QaYwXpZvbLvPLneGT8AbiL1FvspxHCp67uE
PMAe5jf8URGKRBRd5DxrM4zu/YVcE8uLwqwCJb8ZIiAoXQr1g1PdTJX744VY0W2Q
BjpatnQx6KoKAABjzbtXGkzo8Ym7cTkhmlY6e2hfszpx6dDZs2WK8SJdIle/+Jrl
hqLyy3Aufq9jjv+NZw0O+//S1AYv0m/1luRQocrB9gCHYYXvFI+KzHb5CrRigo7+
jinCzGdbIZQ0cbdcQgku5ScU6H4uSRyPGiSeISMtvbY0motp9vU6l1rV6WCzRMV8
wBvECnCnNVY+xZc1yKoN+sADGCc7SJfbH8psBxsGVt4xd2ADcNrOV5s7EDSybIfC
dQJEGwAkSl4di1TJ87J5QO6pMgAKsBSkzJvC2WBi9Rp7yhsNKBf1ilsyBYBj7IMN
bstpzSMJRO3wg73nyUu3OLCjQ1UoumM7mNOIMhKtZ6bEueY7WhUgm/NHptZJaoAz
kovKmLb+dYY6Y9EBxFyzW/DHZbNLwE8BUszu3m6wnbtUfn+xwEqt0wlF7Ql/J7pb
ZfTg/WDLd17Y023tShG5RrC/9x1jT2rgOZXLGp6+ZrZJaGK910zHjMzbFxS/rhX/
whbIeySWg2Dr20bbqobNmSDRwwKVOId0JhrxN2PES0/EbmAqr8A/647SiyWrrm+g
IO2TMjr3mdTwIm5cvIO5dJm6atiib42Aebpq/aE6CdJt5zBB3mK6h/08MFv+PkC5
39eEsJrnGkD6wQjdnXoxTqMopRFGgJH6Bp+ejQz72AGWZ8pKg7xIx971HbT/PUfE
4bOXh6Rn/7YvVi09wAb3V+/TFlCi8xvHhoEKP8aWLbkuaCgrvAblACyFWJcbIonz
Lhq5SHdOPtjtbKKV5EcHToMRpKWodvO5tfnvlfZ9Tux3KfvRCEPMKpA5XfPFDmtq
6IQi+GqxMvevkN/JDPJxxy4HNCpwOtkWcoqBKRHy+hkloFez0jOgYe2A/0TZVE95
aVYtNSGNPi2H/Z3JecS080Sx90vNcXOws+ZghgUuBK5rM//zcaOAkBzVfxWZeV57
p3hueQ3er65mO2SOckbtYbFWlpBtttj+xJ8x44C67cAf4vUaZiC6oEGDufyH0+sP
FVM1NVXdHwcsu5BwvhwVJKAilGas5krsM9afWx4Sq+hZN1ouPQ1gcB2hDbIfOxbU
hF1841+fMNqh6Z8sxK3J43aAWCoMZK66fDGgShFude5HhvL12iRelpafui4er1Gb
cj7Lz09BHB3KKlyJlPdnaDoAgSMa+s07s81R4Jx3e9wvAFDH5b0CbYFVqXCbdkKz
MACsSjl8kWyb0m91b73Qf8JmeoaQkMfplPAwIDZ6ZkKsoyUp9X2ODcbgW6LZjAqx
+bU13nyU9yP6ssxrsqBZpdt2ctst9OWqjVUPAt0ljfBhkawNWlvs7cl+YQ13XDbX
Vp5Y9A1Wl2tddzETNt8dtFWPwABsTBLrAJHortNBlPZT7aR8KZF4Rir+vy5qonHt
n4506ZcuxkW/RxniAxPNjPIy8ooVjecnPCAl8Mskx0g9uVCuv4gKNl0Zf2hv41Nc
2AyfO7AurcHbKURhBCVE0tyGkYOqlgKaE/2J1WnEyxJKL4kZEdcq/57/IHYAGGHJ
baegdfwyfkb5eD5iW0EbKcSO7LO+yc/dbIPZNgz9oRNcB2/M0y6x6WTFx0XhjFf7
TShhXTL34IwDrW7ADyK0jK3dS0DhclV9pMhlDnLqyLgS1CA+i6x4/1acyriplNHY
77KDs3A5GPNYr8I8Z/I9fwsoRgTupmCwDy3zGEE50bgMacgjObi7dyvThEhUfKA+
zBW6kgGWN1Uoo3Tyi6EisuxfZkvxzPV14KsexrpQhkgqyvbaJiynUaBsWBG39CWR
YYp57TFSOHNmn73tCUmADp3piCXg+YHc+zzeJkwNM76fTmbiigE/LeoIvH0N+Buj
lHb58wdwWSLHzr+LeKAPmO0C1d3y/+sNcEFqFqL4H1h3sxpY9zwx7vg0dKcgaIdw
ugNnikXdYODwjBjMJ9NbsGAJUUSiWSmcYFsi8axNSsScnDr4G//yxKVvLk44zXpO
nu8cNEKVPsVuoU0mXB6h235ELculsQEZBLiPNwsOGu5ExrEv+10Y++5jdeRArdRe
8ti9JHrNs5cINcmH9LjHnUkItYbUN5XmuRMO3Cnqg9MJI3kpY+Mu9vQtV5Dp/xPx
ish3+diK8y/w6eOR5poEIEBgxINWZJJ93OLHMpqu1JxearzMQTAyAiAY7kM3uEUy
pkq8g29BnG7KsULjCCdYiOKmlpR0OiHfHpqVciEUYnL5Xk0KOzWh2H8003nixvxO
kLjK78fU8ICw/FuaZ3XhHaq4GQfn53/AF6OEH9NP4PAgBmlUMm7AaY6VSY/QZmQm
Q5IlaK8T2CLolDTwgpolQU+kQAcVfQqOi4N+15pUM1LqK2laSLCuux+EPT/oCqSP
IwhINmv1dagvUl83qUsWsVpMUzTXV7iaz0fGRQmyWp0ld6MPyhrZZncGfZOx5Y4O
SLFRjJj4cMG1E32tCJxFOmWRdaEHF2lgm4SehbbBI4Eai/YVK4FolUR4PfixIGSJ
zFYzWygJDSAtBU3RMC1k25fj0rF8g25o5TRXhxktbqbwBtqO9DWU9aYyBMGZrzg6
WPwQ7zhLp/fQwPZyxZwnqwXElyWRE6lMyGa9VGuRCuTU8OpW0jy56LCX0ZTUAYi5
XYn+tzM2G9o9OEV2bydyo3WDs/TQ7CUL89BcbWnKqfSJe8HvFU6/AWm44xRsiV1k
MhxKu9QFqXXUhwLHhgPZLYjG9XihatSljKa3J7ftAe78UjRsfK96LAW3d1nYXhvl
iJf7GlzInwkmtd6o/Wq6mdEbB4v9010lUmDvRfV0hncivWT6l15wrpYSOU7Z0MjA
HDviXuBmjY6eCWt7e/BeoJppUimQMgwEIXG5aUfbX0Fpj7Py1c8+rAlHgIofTcaj
l2s7f+Xs0EsMa56Q5WhZg19LBtuI1GTvNOzkTHwQuTDIBxUEZxxwIqcQngk2duAT
+HKaDxX6Genxd8HZEoBoLKX0R0eh4e/hnlypWmtS2OZPAsRDGgAjbsdpAY4oCZmQ
b1gyyztqGclL/sDIV+vqJWKQorO2xi39kZ5HmYAwHiLz7YoKFaColqGWLQnMn3b3
1z4hWYI6uqeN3c8vPMdglgWvKALw6oPTenIMh6NoBkKm3MfRFZXhJrZKdy+io81X
0fJVdnWb1wraZ1gwqgzD7wFIjUQRmMQ0xjDV2leowKBLZYbspTK4HtmWbBkjoYZN
yWtCqYqa7FsbbJgHeWHIzD9mmWHo3IXcUpn20HXf4RHp86eap09/iyqfJRzX57WV
YOP12M2wKmU78tSAfwDIc2tchVAgnqDN8oSwNu5SBudwphmUEUtjBEMnRHwtvwqh
OVoaNQ7DweK+JFYq/d/58PoHwlN8MTHJriGInE3S5zjygxOZQ09WduBfyQbxgiHJ
24JVNZblhJj3m1axJB7Z6Xa9kBaNlv/ugwx4/3m0WsrLmX3hWrUkhsK8voeZVPvC
AmAHTN+lQrwJkl4w9uq4dtQVdNdZj/8R7Zwyb8sB3B8V6Iwx6b9T9ZtVLLK0AXLC
LMvuO5RM4o8OU7uG8iRvcZJPeMlk+GJz+VNRI5Wlvk732WlYUz5qp1JXwBHvKTj+
f08k2W1KGfQXHrfctykMzZt0yYPj7jAvEJ5zmtv6633LgAGSXWiwuGknB2QD9tlp
pAuZ23YngswXeZS2Jll3+v6OJGhIVZB5Y6eoXooZCPTWjTmPGgothmwUg1fig7dd
BRdnM/TC4JIjPpW9fYbru2eKxdKpxQToaBuvf0oxxV2nC+U/tiM/9DbLXrWBIx9l
U38BFT7BaQxd+JO4dR9i0xk4Ftc1yof0GsrTOSgViZmJdHmPIpqyfRlt4RbIrQze
SuCMo0hBbAEwjJ8vWWqamA74Rp6T5W++ZWuX+rDDvzayt4XYe2D+fWc7urhIqB8v
1kp79wkvLbBlGoDPNVfEsiQqE4fg/zbX/ytEeSP83+FhbL/XZ3bus2XxpgzuNMGL
be5xm78l893sY4IFolvZYa3MKgqwzcXTaAI9U9CV5QiPAjWA99auAJDcAGIJmHaZ
WnkZa/BWpRwFh0QzbQiZkarvrfOMSX4TxMO3uuigbu9MhDZQgnXpjIUYio86hC7y
O4L05AUOdB5TriZvrWS/E+yzBb4bWjrgdJJ1xKWNbWGSxmubZ8xWmEwm3/fbxplp
TZOjRrWEXaQrZMHZPbFGIxzsQoyzDu+mNWLVcv5U295GiT6GcnT/URD3vtBQVqur
E9JKjO6Ww2NB2imQYUhRlkJ/MwifnmJpPDyhD7ZQwGpT7bEwvSffnHu/ezTSey+6
bB7HX1PsCWVvG/LYY+FHVGKIEI09E7FnWdoQy0lRUbKsvFcsprWYSN0VJEx8r9gy
Avi3KEWkcDA6MNqJB3D3T94KLhwmjKuenkVLHRRXNz9AEV4uI0jOGPzItQzGxw5v
8jDa+NIwhYz1ZZePGuq9ZgFgiuDLbCCgRDyKOt9gVTcYhPmSP9NOc4KDeVWjgny2
+eUXebVFtVZHo7iYMlwmiSAwpmU38jj40JngUZQ3GiFiz/v4lWRVrHVxZNaK1sCo
95Lhw8ozkPANRaOv7HUbo1qWVAlL6F21dov+X7Yg9ySfvZVgPV6ABhmT5vqY4EzT
MfvWaXze0Mk5YGoblqfTvgp35saUvDeaRm3463GfsEKZBmafMIiyZ0OXobwKfMER
hny/o+7+nam6iZ/nWk3LOTSZOEH1NgZ0hJeR9M3YbaApElh8XElZi1twlP60hOse
GJ2RYT3lujm53J9xiIQONO7/sFT1cBgyrbikOxZpDu+exPfz9VTp5xMFMk7VDsL3
5Ojp9/Yw/7u/SxysFtShS4VmBZ1lbIdBps0Po4qixn8h6RcMMOCm5mREkQgoj9Y/
2BO90Vf0uXNgPW6v47QiJAdTQKasMztfrmXOL/fqeIcmqqnM1LraQbDx5YplE/QJ
j/bkTZsL8EOQi+b8tmzaHPRnBKH8N2EAupv+yo0ocA3WSoeEMqjFD+Rq/UdQligm
v8MGPXvyV47y31Hn+1pHURA/iyReiVosbqqs5SjyMCLwD7U7eub1hGks52WMZdRk
b6fVUw6Ld0/Y0zH3fpYJcvkFrpdKNv70y65FiA4HWt16Q/j1XSynB+EJuMLGId8P
xE9i36XfCT9H0EFUx4ntiJ0d79ldjRTPRA27qoTBSo2Q+iCb+Tct3bt/1kPWNPax
o8YLA2PcFgTO0NGqqXfBNYfwNiBgXnbpYQkhfvqAGyUomAwZB+PEfOpR0cYkUxYJ
HXVFAB8jwBnvUIGN9jUxURKsu6r0E0EeM52HRXkvbDD5QCs4aWimrkH9d3Be4Pq9
a2qLUNClFzHCq4l2OpjBApzySIBwyExTtf9S3stYGP84qK4l4DCvHuc5TXWGiV0L
oAOlEIyhfzzQ8xZbn2agJsnL/MMDpjhcFcQooQPQ9m3QhtbNKZP1DCB0A/nfAU6O
TXiotKS6DhqCELaCPrtr/CknntL6PpKqxGPLnMVcyeilmfHIuS6WyvjgSdesJE8N
eK47JaO1Nw0zuEIXrW2Ry0RSXdr95IAzC7tvAeef6pFtmt04ZakJn0esyJmx2Xw1
AgcgdaSl+1nnMWfUMHtcMJ1XvGn7YedRWwvD9/qzRqVDVuQUfOcqRo7dZQwXF5mq
u7DmQyw0+phAQvWfy8gvVhdb9zgOV0mgg628FmF3KstTY/kIC3k0y8KrkJFsABIa
Em9T/VkYx53ez6cNPjAv0AoUF2PFwgIhxkJr3s6TcGdakrVMaEg+MSNYgm13k2Ey
bT5YlDZme/Wp47rGxf0f79qZj22MFG9kEnVLkE1j2EHgrflRNYGmjI7VuxMQwOcf
x4Tyenwfs2RdMzhYpQgb7FY/ScRgeDZgYaFq4l+dA4AgiG34MAwvfIWJRg5hUh4s
5teGVvbVz2mO6HiAg86rHaAha3v8j3xRE4qRbl/GGdRJUIYHE/cvh8kApNzLd4kV
AAJPhRiZ3LVsBVLxNdoGlrD9KwZTtpzoiZvK3GB+dMuAw5VcCocwQF0j70R+uSAA
RJ1K2IAWeIpfhGSTHq4zG9PkkAWFHNv35sFxovekXzu12mEY7cJ9cKdoC7pR4gMW
RYn541OfYoxfup2QREn/DR2p/Kz20fKRSoTS8ga2Hzse5RX5VsKlKZuASW8tuViT
MeQrBJYBSAZNsCsw9Lu8NIuMuo7Xa9qVFZ6U2E5JvMOtMlNUJH7oINEeLSH1medD
1GJORftwif/FN6EEoI/UEtnEyfyP6WOBY4AGViAL3WS+kGYOVufoZ8B04YauO9mK
aGKeVRQRD6XxAlHepg9YRTcqxWxrsRTyTy3+5/LEghLEE+E2FB2wJ8Ch1vuil8V8
q0DAM1j5DJfxGcqUsAoxLg63CUVZCcY7Ka+dDAyGH3vUfrhLacehPcXNPK34LFxY
Lwyc1VT82Grk38dsbq+8u0a15lXWFYJvw2PzBJZb4bPjHzj08CKT7xejEonHUDq2
Bu7osQAjRobNFR61I+n/4gwGBup5XMO379RCuI5iUY5GTtjeGbV1L5b5P3vSufdX
/Nl2i4nt5HWNw1cdYJ+53w7j2WCM0IRxabKXO/KcMIYW63ak8K+9yhKeXAEtMGVN
za1toodMtUmZPBrSH7IXXjlDdGNjNRcRxjOy3zJohApGMhrOg+W5MAeaKa2kxDU9
XXStys/3oEBKkGg0hg3bqyK0fDjTG0BBG8q0sSXtYBlWyzGORqwxfa1gJoju+ynv
ax2Rj/2z+QCf2TivUbWU35pwkBOefBHRsbqs4cGlIDTTPvi1C0eCH1eX66qkeGnE
cBTjjho7WYhFyoBDChNZ15LMZXntFCCWa+Ph6HFeENKe2h/uKANu4P5q71qictRX
ds2MjuZrJj2fxHlpTycO5O/UxvjTGGauOJQp1FevyO2M8aLJlhF8hYe3bUjIEKfi
rr+qYtqxl+SRN5AkSXfoIH+6OMs/E0XgiUOm0DHPRmSQGjETBIfpRE7zxzllDE3T
i713httQxY+jHFi7boYpwGkBtVUjW1iZYRQR3UGh16GJ0kV9J1nL2wBgeQ6lvhNk
zfpP8fPMAQPX3msGKiVgx8PDWaYrKytOfUVhhi+Nm4nhe5//nSySys2KCvn2GBiU
yecrdyskXcWAdCWhr+XJFfBmf+7so6DACyteTGyFgyzEIoC3IxtOt2M9HKoDkMRh
jMqNKgbQr1FyGX3pF23KOcTZEdZVgVc6WtY1uY+ynfOB5jlclC2tmda/geuoyqwv
hi6aJL685Vh4Y5d1iZFdQPmMdRZMBFBBeD9TMfWhqydcvaZE0vwf8LWFBfm1SRQ9
hRsggNAplM9NDVO82jx87VunG71OZ0jMgeqAApDb9mpTaY6ha4tz1x0+rN+4jY00
9s6sz5DNrzK3pW9sb/OZX2P1ka3vdpBMJrFpYJqRJ3daJtq5g4Psp6Oi8nhMiJPX
ltTlhhwDqF2zip8/XH7IS7eW2Fsu1JOOBdRiHUIRTlIXpuy8OZ3QP5komdraPIsK
UJtz0NNV+WgeZLD5E4SkCf7VLEyWldx5gULQxfI86NRUK2mXk5+DNIjS+fqNN6lP
ulDhA2NE0zmR1+hYbMYTBZE+IkxeR5/cIUKKGNLG3XKIhgz+xiimBYs7RTDr4a98
nzOeTuWEI9rtVPj/PpTLGmY4yF6Yzasen1LtpPF12cDXGAlbDbSgcNWNYXJaMdeQ
PoDK+xdP6pT+uE/dHGcUpWX0dCeAxIQES2Byd0BYxmlb2syqHCwAO69N5meHEd9j
llyyyN0UmCnxyiGtuhYZOp32VZYE3trpeOp/mGgedUxbtHyDzaLFXGUII6MbzMfE
4I/jpq+xp2teWZn4ZPArtFDJ5Cujds4PSkwqCRE1eOFrWn97o6/H8LLRLv6XXCFn
mOXOPjBgW1wT7AQ3X5hoCCNKJSrK5JADv/j7Fc3tLPJoyQEDQKutWijR9/cVvCJG
KY8oJ5hmKkQ5OGtdGM9AjP0yf8WmmN0ehizffSu8Pj4sMp9buNNaieVPnk06mYOp
POS4hvRqp6S91YpQJNthFTc7VaWzmiBSkRgoVXwytrfR+ebQLwJymJ0bSZ8YwQja
EFA60ZK71xRdhh6fpyzt41nY3wWB6xl72PN1b6/Yux3oxR51t5lgpc2le4dhYZuT
CH079SbbD3b6iimDAZdUf0NfwzmqvqmvUcDrbPtnqLHceN+ZvSDyUXph5H1hiPbh
PV0jN6Nf4ZpmPWEuCgPfrb7bP0Im/8gilolQe/6H/E+xTfzFY8c0Qljqtw6qw/R7
71NLfr6JMCGkTltoQPbYtwT8h+Lb1kHHR0gmbBzJ9RhtdiDis9KZWKid+7/xhyMZ
DnuM+l53h6Owz5iwzgOrhibPBsRKG1nQdnoExPnSnrgfVPnwwdb5DJHUnpz85AfV
8pT91iRzOs7rJcX1rYJVj8WYdodrJ/JzVE9CkCoic6apV30bSIsQq3JnT6kzWmUG
eepBE3YXir0TXLD21DvZVT4bvEKEJX1VbcHhblEr3UC2KoxkS9I5V/ztGoFVJ9xw
v8hBN8qVcKorMVuoPAvloj+vaav0gZ52hibfIhaPmNPeL9PzLQV3hldWoheoXxZH
uCKyoe5te6DT4Cgcwa/6WQiLJQfPMZ+UkugQuwskWhAUII1YD5OnXyZ00SJjZbOn
deeH63z7792o7Duzae+MPFlv4P6vLEOG7KFyFYYcvBzpz2ca8R8yVuniFBylPcOk
Llial2tE4GXzvBq+jx6flcKwjQvgFradvCVHLuECr0egpsQnLWzSf/YcL1PxWnJM
2+Y7hi+0Yea2+I89BXXCu+F8CLWsP8MLjMj4zdqied3JGiyiYrzbevRnOcHQgwOW
G/KWeGBZmNCsl3HA3y3proCQyOR+ZjOP2kW//Re94Uez4B76BkNszO+0rPqnG0J0
N8swLqCEDS5Pj3aFM/nAwRY5ZWoCmmEIEKDNuKD4kbflY2BbjRjHK6xFF40J/WY+
3X0engu7BjuWCZnFEsIczbmDoEreZ2LGziyhAVzsyeUipSC00pkCZoEtuM+trNpL
6BKlDPuYkuoVNtwVcA6aAOu51HvtXt92v3ktxczhwLXuksn9G4+VP59o7NEUaJcc
wU8+r2MyY2NiMlRds1P8xDT/59JJQ2dPALVGjEIULDlEXoD7HqrAfMld0hHIu2ZT
t6GuN8HplybqdQgXF+1B3hB8BPHb2gj+5rvwG6fteyCJKNnoFqRocNeLAB2SQH0w
goNbTfZcC4l3s3BAeoK5Z4bnVAmwrfwlAM9tck3NCOJL+rbWcIMxyAyUj8pLm2ky
oC3TkT/4BskhUsQ4JDk8piqJFj2FC8YMy8296XW1ZRudOf+AscotICA4UwknSTo1
5oxSeT+Xo33sMxp843yzBcISXV5bP7Xf7Rw3figK/s4MzKQfLw349qTftS74Eqz7
ELWra8NAoJ5xqQbqd1C1Fys2CnVQgCRaA3na8+suwmwDabnEaVCiU86fg9749LAb
A0iRZh5anGCwJL6u1SVR0SCxPMt64OAtMCdtwQ12RAw2rBWk5AtwS57c3canbNQq
x2Qsxtq/MrYN6uoMoNUtsBlkE732Kk9ZMIldYxP7Eb6vPEfR1w4zW87wMuWFXNZO
X1PAPmEmbFcCDO1I9id+EAXEModOoljORnz8S61uuM+p3suSJKJ2bF0ss2C7btiN
9Oq+1V4M++Q0QhQTodlXQNwl79sIcaz6VpUKrc+4BimoRlzxKvkMLjcGusfLaqKH
sPFW4Rm143vH279T0Fyt2CI/KmfeIEGI1dMl9CbWveY1bxnrQDTeW7IEg6eBS5bM
zPsKQ3yzGEgI9VPECTDPYIt4+3S0vksPjD0cU8PvgxzY0t+LhTzIJZtatYrhZFGM
31bJXZjUTYIaEH5wW1sdONbQXX+LlIiRhw2nu/hajzgHdTZvfxQswkE75VKZxrs6
d5BembpF4nlx3028ocpQz+Dnssc/hecY+mrMYfJBXMN0YjWzFn1gjuYkBtZOTfyd
YjE6cmkwdM4zqGq3iMJS0/oaPVkPtgOphnO4pgF9suXRkGdP2VhBTL1PW+znDaxC
4ZcjuUhNIMsC5gb/H5ndibxdZfDTpARb7wqSmBwV4EjTo20UV8tX+jA8mQDeW7+T
SfRfc+GlXjw390xX715VfJU1D3k+fnBmvVcU9ZYIjnFkt3/ivQmtv7OOsHZbfeSc
lVDND+11FWYfqzjZnKvQ3tPFd2FBY3LJGBQ2F2dqcQ0TrWSJrULAzzOwQLmAW2b9
8xZO28G3WoOCvDsUpuC1x/cK8gtBP4o+b0sVtP7E2/tlRDyyfner4aIrQ1dNb2Hf
TmuiSgopstc81frmXFH7arbwMoStG+1pp27FJn4RWpQ9CGpmBtHMwUnDaf7akZDF
adNpK6shEV0qd+yA6HgFHVvfGxYN+0hqi/3xugDXZgLITKQxQG/yfgWxw7nCwvto
3Vvp2qRUVfHdILWjjqfhwbIAcTGMw/5E3tAJwXdT6A2Kj9GGQWn84IpX39NLUxiv
BpA2aPKPGfvpwf1g8Hqnxmb3WOOQtS+/yTsudcZ0KB7zdRPD5VYlbsdk3EY+T6qk
RK3OwBHwrJG/5A7SfZKCImPk3yDC+dCxrT3za10tGZXmdlMp28WXg7S/MV3H1v0Q
9VfH+SSHy9SFwIjOHLpt8RkzDGMvABk8w+tB/N7F4VI943o1V/wiEru7eOSf0bSv
YnbkmIh3qf63j24GCKoryqcYOhj2Otpfjaqmqhh76+t1kMCDJv4maQanwKvc2Jlf
hHarl1GujekmSzvEEDaqSNFCX7hslNxTd1gMBuzkW0ahpcfvcZlJsUPIld6O96Ma
UKlJn8CqRveWK9hwBWRVL5lE4L9aaEHsxfAoMNPmxDLyiGrrwSIMniM9Hg0VE+Cc
1hrp9Fz5A8oup7oUEziqGdeKYRmqIZqF4KDkIajPjLS85TSe3Qs2flM9Yunw0gC0
lqPwGf+yzWbz3zbgBSbK6AdtQs19fc+mLSTTA36qXk5/gxYq++D0K+6l5tlUDXFh
pHRC9LC12dMQuwe2hyApCy8JgGLn+FxdMUiK9J9m13bktYn1sCbb2WDTca8s1b+k
gOvyScc1++nqpJ9JZziaa/Qa9cXpistYe70qLiyOWRa8EmbJ9DM2/+Xfd1k7LgLR
fZQ5ejYVPJhzN8ps6QaFkKGPve1n5mdPzJ+0oMlNY1tW/bRHUEOY5/Kr7/dcCTvT
/WE2UJB1uFYjkMBLslrGT0rWxSugVSRclz1pDGxQZ2uvhLZsAtgMcOv8eD3Xvb8A
6AZv2dR9ymluar5Gcey6/l0ZRCucSWVR/DWXtWZDQ8xuqF7OsXGJwF/MCJR+RBgJ
oSPCAugISx8u68lzZoRUB9aFDm6GKBUA6avOAL9kzxWNWVSr0CJ5u8j5mSCey5Nw
eEHK4UtxH8swZbVf57UXZIiPEfS1jOB3aPKo971CFLgpicYnGTWk5BBWIYC6eLMW
AaDUYxwkewSIjEQ7RdJ8SAfnkP//N3uTYHNq464eadxgpRwqAE1S1Bj5a3OrbJcy
NyM3HGaEWqMbeoi8WW11MvZr0gGNJXVJGRCLnv6Jslz0p1p6WIvesDWgSpdRRnEu
PKFpcTnCsukRq6YVh4jM4y81ieAYFL+ywOSsCGM+Pcycyk0nwt7sq+2A1wtHf/gz
AmffyvMrZgudv7jKYtMMIHplwA0fjWFN109r1irh6O35wBARaCFZAe76yNp0mT1Z
Oln5zynyXjjzhmv5QOukBpLoI02ekMgJqMPKp5uPaQjW9TYkDo1P4IJsxlL3rW8d
wM7p6jfbOz1MyQDB0qRdMEvSPmOFpS+YBCSnckWv1NNzl3/EcOHvDN989qJ/73pb
hN7T+GU95bXZAXYur6K2xLqluWd43hntHtrSLlkcFL2YjyoFIWlxEw4MiGnDUxLc
F6i6SlI3mfmJay6yqraeaWgX71hdnJBNUepfVG9AcqdGRVIme2Oqf3LX2qfXNuTi
Jl0UG2QxajRK13PibuZpdIaPZ1PmuJmhLD1TffdGy4izNdX/e0XHEZFbSjdZLToO
XlWszMm8qd2t/5a1dxCVSl5XRP4Wg5SVRMffyjU1Q4y244kdlRtf8I60cdyOtDIN
K1mgbSeFRLBlvHKVEo4cGB9r75Q3nF/4dyA1YH1FH1Zx4lQO8G51axcdkLAohUw9
Ad6C6sIwreiw5bCDAKOhTeU/RArXGL0/cq/3jk/rJ6MZDI6Cm5E3zaL2836IPlR1
MECq9+6ewUPytT5s5ncB2kZwUL5lmwx0HsTHINli7OwIjZfqA9L63Sk+QY3YGoS6
SbiUIy8fIFJz1pDTaICSP1vxq71ntnGX9iPi3pKqPsANwabhNo3gAkQHcZLxod5w
Gk6/7U2Vb4MVJ8+WP0TTTIftcdyM0uEElpwzDlh/WcHXSh4dEM74pdNafEyyYXRz
Jee4q3hpdsFKGxBFGUCLXoWZHjLVJNjtTrn8TjCc3S6tigC8o2/EoVbCNKOUfvRY
KBz488pBAMwNDqh7v8M/nJTlhekpMb/sTIKEa0QLhDXenpBYKg517apD9udecBqy
k7HRPgJeTxN+J3muvKSHhVXaEAA18IM1N7E0RrwQ51P+mFuKPCcxkZok4PpwA1yq
A3ZthNNmbPbOe0DZZDHod7XDBa9bZLJFDSXGwf9UlsDIjyWXLe1zknGrHSzI0GVo
YR3fDMHpuOBvakF1aLGCYbZSdHJkuc0hnOqaiu+OaBLWv27KbQJ4iGYM2xQZkc0d
ApBpHlqLiPIpLFMmN355af0Ha8LYpdDtVivtgQm7NZQajNPm+uH/zr8adW40p2IX
bgYw4NE8gy31MQA5kwU6ej6GUrlJc60zUESwyeHxtnNgMJNRpZFQFSLscPfWCs89
H6gRYWb8Qu0I29o93MIJoMiWE99yHi+pAfNWBcg3PrfI1DeUaKoVMEBqV30Yccuw
d/4fJ04azQgs2t4tfS2H3VshpRwpnu5lSHZDDCiSqROJFf9WND4c/HVPAf7n46kJ
CV8REEEsq/KDEsap+P9KO/msP/U8Cy9M0R3pTvHmaHyNldfQtqwLrtKSK2VOa+wW
C35Wq+UwynpvDi6WWMcw0z+eM8HuvY3U4neu452bG+51iA3PHt1wNOC4ZPx09Qu/
FkC6Og85Ce7MWE9NmYzmOI+0DLNxooeS7fOJyzce2TFkDS1p/xZkTSDoivo8G2iZ
iDm+xYG3ISljaonsW8wLAiZXqLp2RhBTAVSfVJC3a3skpsTR4d5d7cUPJL1TigVj
YdrUldQUoSMOf6VkM5Gf7i2+yRUXhHFK7uUpYckiLCuAckp/7v1ChJghgAepPqPn
r5f4kEvD5070srEUjoMHqLy1bn1nh7n341YoxS/jWoHnf42mEoN2p/xFP8CDwiAd
xnFSZkbi7Toyh5FLaznJzdc4J9IjbP8+4FPmFFftWh1DpNHiVT/ElVcPsj45D8Ku
rBC8l8x+nHw/5BBSD4ydByUj/1/U48EmswV5GZdb9ABV24gpJM94BFEJVKVJ7dnR
Zji4/Exv61K8n+dN2IuO3ZMG27Dad1w5pz0IVof7wYgmCmPIOq+rcS8TEi0/lA4J
8dMXtcl09OqhxXvgr1XTEw4aVSoOssJQuB2J3jbVwiTaUcR26Iw0UcdfD7hKY7eN
Rlw8S/TtLAzbdLUNRtYtGUtE+pW52r0shEbO+BLejueBHvareLbChgt30pYgp1WN
C/s64hHsogdZbMIkArRgGPueYw4TzPB8igpnazY7rsjwSWIlRyWAJ3L5vlWtydcG
LGBSFc+TSnpDfEnBesZBQns5ErfkN+G2Xh9lnZQJo+ov4ALg2lOoUeEjIu59Jstn
ohII+8azmAmu3gQljiJeY8hibDP8mNRDND3TyDSO0ETLj7nI5a09jgGfqCqDdw2O
QHaxfPmtE4oMMdhMciEUfVGhcayHRkt8Rct/XdtsuJw4gsnRnp8XjCY0/OBkqhAu
CwnaXRWVANPH4hprImvt8fpi7oHmF5DI+ixEKkjFFq94nWJizoBC96WIKTm6W78w
mTEETZHG+L10cJ/jB+gRhD7/hJR5p89au5tFR7UKhPQwdzXaMOTKJCyuVG56veI3
oWTcGkazl+rk8fQ+eOVLxt9Tv5pEmDDl3Er7FYX8xgeEu0NyYvnGinKHYj82U98+
wEqYvqgcuRgiGzUqPRUZc9VBs9R9pNhoG8HoBRpqWJc6MvcElj/8dN6Z7UTlY6od
e6poHOXTyJGwar5eLxp9dQ6+QajVK35wc+G25kscY2Qe6A9br75hsfwjMfpxH1Yd
JsjNMs+Pui9U467/RF24/r4N6t+RZJ2MCS9trq7JjldY4vDoXCdxUSzn5Z1AFWUf
9LAgN9xCSzM/MzyP39fNkVLGxhGWEPcsPvBIr9riOMxA0VqfTrGT088k8YukZ+C2
izRrxsqmnebzpiKfJvYx5P4G17+q2/k/cbzfGzYZZ2KaejhV3d9ZbtVLfn8Gy+e/
3BmesrTMZlnvKcKlz3cGxEI+vtIqvY+A4fwEb/hdLkESrszHg7+Yi8NivYujzlDD
X2nWS0eD71ktga9ATi0qppxaJK+uL6X1cuaDWYGDk8v0CG1vrVBQQiMQn17A0T0I
TMosyESMdrAtkny6LEDbWSmfSouL9ohkjXQFPhFRqqqCvcbHwl0oLtse4uoECG2G
LzO7ObG7vjnPOqB9a5asIFlen74A4oF6x3IEreEaLkT1gPPsU4K+rmejYr3p+GUR
qLrceBwdbrv0fkD8FfHAYBfrBJ8vBT1yTiAg44dn1ilt6OACaaNana2bAhRar+7o
h7QQ9uEKgC+soB6F6pWWkDs/iG8hMBC5o2hL+8ttKPL27IJjkptvCIk65EBn0Pas
vsBS+eHYBebyiFb+6h+miDLrib+t7LB9HG+a7MNtr+7K92x0OQFFmKsa8J4BfFSS
QqdwPLptNEjKuQrDjbz6Q1OLfbut+a5CIgB82wmOJdgzJqagLD1uqbUbtJe2Ph0R
3WLd/Rr1TXzudjUNQmG6aOzSLFqCvswEuMEcdRrY3kw9Jusl4FMRsyYRfDHp0jES
DXa03XvbVmzUWt0/VM8ZNWRbIY4lpgb/HPd14EyT8XQ0CjsiCTq1QilII/xSLgYW
Fov44MNV+NEPlVEhE+JZGKN5IdK/puX2CVOpFMsFWNmXZwxg4xl4dkGjc5r8kMyF
+glzNxHvptwgRFZ2MdrtZxzq3XOVwEttx6ATSD8NSBqbrtguQdr7R1ub0QC+7wJP
tLRvSv6PXUTS3t3yU5AlI08sHiHdi9HMiwBajp+9hIaiq0uNO7Rd8JBtmV0sDC/7
6bdRmNfz2mekRMhslaNbUORlRV12iDDJhF/cAb1wlx1egWupmdOhGWwNdC+LKanY
DldT6SjIyqAFu/r0q1Rhf4abJTphRrSVpoB18UFoehyDMP7USyRDDB2NjKDCW/T8
IQowJZ/7711Y3CiYtLQnkwR1a2Va56P5jkO4KxORq0eN9fSA6JO4vZX57FUdNe+x
MDkcUWqlkjtM75JMjeScG7NkY9Jv2iEeXtAzk2cNDXC6PaGrm1FuPZVc0Bo6DTGe
G6rEFbbpGN4Q1lcgueuC8yGLBMSCLJFL9zkT+geMRRzhXY6GFOnJO9yUnPhIs+eq
qlYAlXXSscrtKffD51C/F9N5DyT8IcdsXxteT/hi8THhX2ArpEUZqkNGG+q3xPlM
r3EJ9pqhUCtsNoSJvUyXXHwLiS1NIfBnSSjMZMAOoNm65Qhjajt+vMtDe4j7/8s2
i/1ZRICKfvG5ejsbji5U4S9636c0OAkMoUsPa7s3LDfC6c25iz5ZYfYKxN17Ndb+
+ChQIL7cU/Ssob5K+HO4fgfwLgkLi99wPwoWX+UP04T5vdwTsojYgu5lObV568MD
iXUToMCYtdlTukZ9XsunhDEKuyof+FZjoMgvk8JjJi0fjXpbXoKHBA+5h5K32Sli
cugDfNg+A5jNsRDyJUG+KTQSVQTKGTFldp8qi0EqcGPiE4De1eiOezgwM+pEzaAZ
DFo/FqJRx5hXChW22IM98p3pLhpVrI2Jkn9U3wdIom2zaFIljPvAsKu1hp+wDES1
4Tj+8h5ttS8Wu0HiKusMYbtqDllbvS/5Umn/cCWVxl7O8pKBcCU3zl9vkS8z7S3c
qA4tj9ybG/CkT/WKXDY0HYdDkMwZw6a7ASYUYkd2v3PykDB2AOxf6HqLNiv4BXvc
A2LM0CIlyQLNFUMMxAqTszc8IkMa66H81+ztC8ovIDROSFDOE2HD4K2nSKwdERAc
RA89/gfQXxV+3MUPa3HYp6KB2acMxpy2TiydcYUb1AEZ1HfGGJ78v+m2Tk6Y4KfE
AT6ZkUONMfudT9PRXeLXYvQ/XusuHIfkzsjPLErwwS6bihQHBMl/nkXiEFYIEUTi
BDClCOhMTcdd0Ze4radBHxt7NbUvDDzTd92XBcD1Zc7JkIGcLn6/Ccfkegv3evPl
wp+K6nrDc9Z9SRR1oo4mY3NWRvhKtLAWux7V1eYSSFuzPJz/X3ePIHkp/qbkT+vt
BB6NAMMAQbWrmHEHLDWK3lHVGr3mjiQMM3IhSzCSOp6o7waLlT3IpbRn6/1m8Iye
F+vYE4d5C6YInzXLnAdoT3BzIkRAwoLVz7ZyxdxKK8SAfnW9uzvm0m33/+HdWFoR
8g7T7jtUaNQac3C16EIa8JMa+44suqqU72eddd3BrV07ohjOAZjdv/4B6L3KO1ym
wL9BAmPXRcMnVwel4C+2en0+iCQXHhQQpUI4r4Psy3XqcBTIWFCuOTmxMkq+bf9Z
tiWuYZ6P++84tsuY0/KSGSFRCjUnm7hl2nZdkJek2QuQlU6pDUuAE3dZqbb8+QG9
Izpn8w3CxARwQK3V/e0s5GtQFmwLr2SglsSaIscLJ2YxyoUm22fTr9MviHeWZEEN
A+lkWZnc6zPcoXIMv33M3Fli1DTeL0Z2Omy+JKKz1svBFEDJWIY7SilWyfDBWlRD
XSNKqrGeH4KuJ6OmEaeqvqIK023mVd55pAVouZAD+p4AQJKu1md8tOTTBfB3grNI
EyVGlzphPD+ylhJ2Slh3TgoWOJQ7vhPifv7hzYL/0OJ+Qbq2qdZx2C/ia3Xaa7iU
9H5JC5qn4GYl6XwjagiogE+0E7dlQ+TSjw/HpJs5XHs5jdKX4kqVa6X/vpcen1kN
VU9Ygvu65rMPzh8aG/Ahv0yLNThCopAcKz7DoouSYePjMRpfFwk/1y9cCcPDimOu
3ecBvvrqww1oGwrjUmfEsk5yM8n6/W0uga0j14/jBheE7HIY+/yyUzcaeOntZvTt
5hTfNTD1a6hjFJ7PesYFO6fhoV46p2T3HV0b/4IiU7YpptJfWUeB2hpELChTlz5v
7gIz3320D3uUje0Ro4wCMUuaNf1qfokl2JxQFZA4ZjKR6TL6UiGI/d1QFGssXB5j
p+pBxeVYZLfzZhBa6I5a4Ah1K4oZ8mpE+1yOPqV7rtike3Hvbfn+ZFfHrsAI32Jp
cZ8/u0JvAYTsZF6qmhyNEcN1QgXPbRQV4vjYBg6qjkxx/tZ3hUPoNH9EH914gje+
2YDRepKipv4Zu+Htk4qyx+/E0KG5YWdCQ8LzcbGMgIVqWgj2N1ene4If6FnK1hty
GHTV2L1mq9G2mtmfyTq92zofEC2+WyOSOHa+/uCBaheun/JBVcDlP8VnJnOfjtU0
+vthlHKCLX5zWWAUPKtwUP35U35WLM/7s5v0deWBipYryCTrOTEdYDt0bW9naemj
VzuSIYP59mtEh1D2o1SbKJqQHKLPXEsoKXRMTQz9yrmz1GfOwxbNfiyDsBWiOeRL
Ws799GnY+ZBmSckIL9UlgldnJetMWBxTBmVQTZJnAE6zDmAG7WsjCsLGYsDwv9xD
QShTR8maP+Y+EyvodYp0NEPTKlStzOyT4RPHo4vh3bZb6etZwm9Y1o5LNw4WfiLa
XblxxeA1Xg2CPXR4t4IoJyXSmRlL7tKgyXcR0i+CYJN6R/WH5oNWDeFb21ZFQgh7
r2kWe1J01vvjpsyQ2nstT0qXZzQALK1tSRcxvTLqZUn9BnPjQcpag3wNjQMFecpL
uUjSzIMCA7wO9NNNE1pASW5V94kkDQTxY8r0Kh+yNnxmlB9y/r+cYJpqzJFF83e1
FCa4Mj97tqUHrS4jVvMuSCR3mpAB25avVcBc1OGBPMJm8TxvmlOqdfyzR4GFXeEy
pi3yRdLngyUo2/288Wzo6JHLuN1cHOorW9T4Lg/FJ5Q+ubaAPLecoMIMqvq4LTpw
8QTWB9HB4mLSPsFs0GdHVrUerq0TadkX/8u3JKSWGuGQPYZHxyhQo7EL+BrMTl+G
UORvBw62B5c5Zggem4130g4Ws3bVn0F07hlTDrerfAnvp5rRZQHWRoGHGq1QamTv
vjKrStLBR1J+gIL+WCDTU1p9ErQbqYuOIlVCrvxFnlviw78cwkfmPneVBSLWEGzL
f97B1CHC84l4+oNzED3WchdBIU1lCskQc4N1RP8vEUa5zdOwXxI2eI6GlfV4Vb6K
5iTOEJpjPYNvWp5Ua/tsD9hqr0CO8wzEbJy9M3tLBjKUzSinvzqRptuIw/yR13dv
7YUEVodzXFHI6Ca4fudchMRL4WcnxvE1ee2mAWykLm1vZE+Hj/YLF/rIyrTPKIFj
vFrLa7qAFQTGUKnWkSPFT3RFY/gNZHnLu+1KrJVv3ijjAd6meWIuYVg6OB9G+lWc
8bqLdBQCmt96lvpr42Cg6j16S1PmHmhx2Ls/T04reaTcOGYLOxVXcrEo2VlkKhpT
0xN0tq0uBoD0Dp/7QKQXzL4jN/FQDOKwoTrwr9y4Aeumf7XMzwm7jCndhms1d0ZO
Duu6eHwsjjQ7VUt3BF97hQlwQTF+iViw/Z64kfLC6vZO6Xv4aNhKwdN2LeQ8MTRt
N/FzDdtG3cJmbTZIbBooodJcIPdn6+ivjx0nlIFwYUvmyebYZTKVKIXCEj+bmYkT
9tc31qHFDqGE8DtkZdQ40tgOCEyIn+VrHnqVzbLPJw4Rej5CR+CGs9MSjEh8R+W+
TqYArYbRUAFXkjx3uSg7LGt4IfUgExn7f5AGiTT7/PYSq8wFG7uo45sWfSqZnZh3
hky8YwAYOEwJMA97cjHR7Ogjd9K5iLFQ1b7cP4+E+q+xWhlcfg6yQuXKK/JjhtSG
IS7P4KCkEHyslaE05u4A0m5wbIku7CUyH2+chi1jSarVDCqI+iL/JMtlY4OX57+u
ut5PQze3VGnKS9SRlnrZgLEgo97WCVYdWfLLM5FpZ3O8zwzZ9gd8bREBUePIdG+J
FOUoCfpn8uzNds+s5WmdX1PFm6cMCjqSEGRRkM7vBvO1xiN1doPW+fTrMK87JeWc
GQO/3KjtoJ35gWOSBfuzmTzqcmWY2wO17Wi91y0WSUrf03mC1aeL9ogrnplwW47C
xe2URc8uC6qHzdQxoKac4mDVdizhREZJgu4n2yU0Jq/wRRRyUDxxOvyDRS+KMDJ5
ryUFgLTYr1FF3xE8kYVMHBQT4c8szFpqCn+6MFTDQ9/eTbgqrfUMx5P/NbbQfT+I
05q8YlS+ljcWRhYiH27TEok6DbxnHYIlTi8IeL6GlGf3r1jpPv5xdk/Ltduzffvo
z51o/3PavGboauOfKgOSCVIRDJKKBn2QBOtxnuEmpjIO/e01HpScrWn7pT8rSgOG
mwBZo6tD2HkiKUohCJSrykzEr4L52TPiU3TiKuwCYoxkgRINLl8y94pJDv7FIass
OtKDwOtPtRavETKlT9HRN0R2bYMPnO2Q5Gfdf0831wDJiTjvderYwYFZGCPs1Xbt
Dxf9nvfaezGshXxZdZGwTFgUz7I11D3kqxVR8GRBg+KkfQCtGq1eA8qOWmPFjX21
kChan0iJSsU2asR4SbDpJyyFu9yPQzRyDPLh3rGIYQpYygUU3PYKk9Gr14Ls2yt7
ne1OlEqGju7lq/pX8hTtUMupu0pzD7jjUy7l6HbAGNvUixMEOslTM5ye8/NrC3pn
x5smzq52kOlhtJaq8w4D3fxplxxk+jGJU0nSvnsRWZ59kYpTBUKb0mNgZJUQeTYX
23Ndr4hae/XC568hhueejdFA+9EaoaQdKGFVZ0K1fY8KfIpdl3V80JFXzjsI+COf
XvsnArX3iM7boOMqi0HeGxKoE7ynm0GMQ9ZjWrhCY0ZCrc/x4Z6BcWn/y8CuhGAu
n6H6bbvcKpRO48I5+/xVMUmHRBmhblwd48RZK4rNdYonfeIatWJjIDMad8e/nWlM
pFwb3abl0+cUkDQGWVVka9BdHEQVzufNqteAuHN/ZZhmGlj31qTlEQxqfwL1i+vw
gjPN6cDdSMAfXMnwirJ7VMdjtFgaJ9A9qS99nPH3+Fah+2GEQSmqZbH4r7uSHTQZ
DvKYH/hXg/SQqNdRXAgNNCBCOoSEnDQO/gXrNbui8lP7rRL5zaFnbY+DPOLeJGe/
uNBJPz2GpBkDfcfQ2233RbsAXi91NtDLLNoB8SETkReCJV7ztFtdrZzqCFfeprJO
XpByusLrJ8dSJ1yZk66G8WZP1kjUPWvuzJFqWgEVCYXrvLs9odXu/2acU+E/PYU2
OxBEljRLGBBquZ1k8BYwAp/b97IJ+07bMLjXT34LOr2E8nzNSLT38Q4Sakow6nWh
dIjStVZOprD0W8RkmoXI6Z6hKyliYmmJ7RAK91vJtMUid+Ze+pADJzyH8vJ9hVA9
+F6a7YuBMyvtXGKgf30FdjVFrYoU1Nu+qaC3y42ZjppGJLIjTsGqpyVYB4+I5Qmg
Au9wW4In1T01UtCZSjLNtYO58AYs4x25im4wIjytZ2+YPE4hEt1KU0TeWYYN6/Hp
7qIInEKU5/d0VTUUDYFq9l/iIzvoVEzkriBLYwiCWoktRrj+WnUgIbRf9PMu2JFS
xfIg2oGTLYt3yLqmMN6WVqJcCE/kw7iAol+NHEXVPH6wFpIw8f22MzRJkkJavUcQ
QNGss/uUfFoNTYSDtWAPjJBJCq502sgoTBC9xoZHn+WFF5kbxCQO54RXUnREzlrL
+YG4b9o3aL2wzGHapHJ1tsMFdBRv6AcqFiFI5ndutiRUcl8XyrAFPtCLh8XSupiR
S1xh4PRFNibq5hNV9CDhWUbCW8m8RWQxBt9i7/oJq61vxdCB2sHAvCHzOC1KCDIo
0uogtLe5QTAxbKSnDeFYsEseUm24WuzizYaMhfl5ZigMl0hykxR9v6b4CXDTa038
9eKjGf8a+qYDBkGfkij1LTipwQhPxt5ZUDmP2xO+3M4Ct9xNIP/1ehhXGuGDBLfp
oYKNxfTkiBTQN7kW9nEFftow9UmYEUFNqnj7H9QCT9IB/HqM1kPlePjlp02gqHC6
CF1GwPt4aKT6Z8+bCqi2NAW52bCAaNwIZHfKoPpljcaXMcMhERPq2CTu5YaMsHzK
CWsGkeNJ6K+EaOSy1OXMtRJ69Zl7izrIs1IrWpDi2JRYMK7w3UmMMQS25HwzvjwA
heNKRmma1Nt3EXxi+cgWQGnCtyeMg70CV6Ejx/OSXDw+uRsRDzn8QsCUgCwfZQGO
ZEVe5dgwbk57e8k/NSfRnSR5KU3tyX7bXgOBhgRbk28d2Z9GA8EJfSzXDFt3fcvL
h/0hrOpeeWa/6jyAPfp4y+NWASZSGE5nkDSf93rQwNhtQDVzvH5NDMMcGgr+hktF
Zuw+lG0iG2xl8s64vSxNTQ3GG6AyduWRLlb+z7N5HfY3fYIOjiaNxBP1/WGQzI70
4iqtYdzZwv/X7Z7B3fpJCnFGNs1gRIZTxXF3LqKWGVK5KP3BnmJ4C2JvMqvm745P
uzVtKbfAT75jNhNuqP0k743aOKNiyUpwuH2kT0HddA/xo8gNTffTGDnSmjqrTyMm
wozkbwz4O3DmvI/3OzzKFNJqFHndtNNowQq5h9AVv5FrQfy96uuDLLAU91flPAkL
7QfbOvlLvCkDVFvgdzXRHMXbBI63oO8uuqfrEgMUZwAiZUnLj9z1XZDcrCBJA0Je
oatcvYEyL7M/7Eyp88a0bFr+vZtjYZ9tEf66AbfZh5lpWt2yh4ja7fssDgdSEkuB
kJFF3wqvTsTHmKQGWPzTrfr2WlsDV5ZTTM9bMJ/WZ+PBFrpS2Mu7VTjwI828TVws
tIP+3UnCvcufUgxzyszofUJ80dQolJcV0O3CXNOmtre9XHi9u1Z85iBWxHVeIaVl
gYfug7U0ManFqVugwNDqa3Xm05zYN5ZKRdQvI3Zr8sAr6xDYBmM8kGGM3kdJVaB/
XPC/zLhljOhYvnhr5OMhbA3yuI9hnybTtubEQHVtyHGFQ7Qm+4kelKsSlwe1x7fU
YjVZ1gPhRa71oI6cz//Xe1MBKonaszyi7SyARylF9P5zwxtnxIFEAY12NjbdcXr4
9ShoK7VTSvliy9XIl+tV2sruNjer9RoDBvoIS5q4eSI38xFhvf0bucAV7zfBu8Mq
B8JHk3WrEX/kxbFEw/56lQ/Ju8UXqvO8STafnJ9jgZDgtkb5weS18GQ3iaQC3DFL
PYDgodjscaAnDUHPlvI2wyKaGgSObOSwzu0FCzvxGXFJV3oaf3m2Q3g52TcCUpO+
A7BazasmEOj9RlRi10TkJlPKAFFc7BDlhwVzpsbaS31onCB+ipRSTw9uGHQFqrMd
8QV2s6oTMIZV4HOBkezstPdw78YeKWG9M649JJq4KueVQVNC+7XhWt0NaS3U1xFJ
RC58kvF+rJl1ui1iuRRAptRnzW/nWb1IOhir6owfLLRnYSHFNHtAxOqmurH9bGph
MNIYVUPMkJ6lbr9R5GYQ00TTA38mRPlrW8zL6LHd0YXufVzB+4IZrrbAREZEUG2r
qmjrq8e8WXj6SzbAm94bsaDx4DNJOuLjW5QN3DvpNchGsq0bj6Nzimj2V0rH3/jB
ZMBaj5MzRAOhVx6mxvbFfVJXZxPt1Oz20ojCgsFtGJpmMLCic7Qq9+ogyEaEidM6
/eO555RX0eiXICFtz2sUFMTGkpKo6jI//uUflIN4BmK0JAyQFBnGUG3SjJ7/ZG63
UmAsEzwi63k5MftYv2MtGyNNoAZTHZaBXtHiy/ulmjiaBPxfH/PWjDxnmffNFK9l
YjRPxWs3pzrk6KLH6iW9i5bigupTIxuXjenod5CiurYtvGb1DPLrI2cPEp5RigQh
re5vDeY0iOfaMcz3sX9eZ6XpHR3uYP6RwDVrPW8Vt74j5YbEd+PNcLh0TDuGkZfi
7a/E9Vkfeliavoj7ewtk05VRFr3WgWSudshAIF4W9UwwahNsD9DfgRSkWe+bwsow
AiIYjo9tzs4uhPlI2O58VvNI4Ygyj998V7QMuZlvodxEdeBXaUAeFGHnuY6mu/Zy
8bO8nxshhTO3K92jAtMfjP2w0WVMmfROPA1cvmtZgg/yv/NVZV7kSaMI8I7rqjJd
5Gu1I4mmDNigBkP3hsS4VuogHldgtt32GFfOOUHRlvhEsvJoSiZPJEHsSPGnJpb7
P7VCOvkqUf5NdIPhLi6l2NQ/PBbzYs7Z5Z4Sk/hl7WEy+jnSN64qnPc1kXa9e9NE
EkCMMKHGG/amsCsUtczrWUatvbRO0Y0o6UTqz9/F/XK6ZR+3+suPL7WhZGjPh76A
OEG/Kd7BKZKtlVome0R92EhwoToJpzDHkHYBNmDVFT8wARCNlnYeXcwoqGj+zwLf
qsd/aHyT2+f+2t2F0+3uhJ7y4+e227uf8OpEFlU384tpQ2//ZY39FF7dubiR2est
3YyQLtwKRuaOnQls0/p/4FdbhnKpfnaivbpiqmufRcvKY33hWZsiCxNZeSmJ/FMH
bRoHWIIevl5ozpUlvuQQodq9nTwPxHLkRgjXvZx7faYyFplLCGTmybF07dkOxiGG
eHa/avvMd+24g9yJYz5smpvrfHdsD/T4YCRGdxNtCrCszRBlK9IjJJQFwUDnm7gR
HuSHDCPdrEPzs9hu35Ox984DZoQYGcJkDzqOzAvVGfgfYITJ8JetzeudCUAoHidV
Ep6DTQosHgZEnlwBAROesmhg/iwoILxPYfYfhQfkS29ACkWvxsnFnv8TsILZM8Xp
RsyS15NAVnDehjT2YLXtW4ktE69S406dz7YjhAnKpI91Tog2meHXz8Cy6DVwBT2e
wuopI0O0o6V/Erqzc2u+6CK4T21Ext1H8TqtLtGElD1uGNjAyib0DC618NcIb+op
WTW9FVPgpHu1kKNTBSrykG8GyNOfVVpmzuZCNw/yXnrifk8ZIfrZaL/bJW3JG6ZI
dvJeb/jYPaufJhEqhVgRjdZXIAdeYK+9s1YVC5zKCp6DcwKbAc3AFMGJ78jz1MDW
t4y1xnQwXsaOGNX3CNot35lc5wbk3TAnAG+HHT0A0nJmNNulGn9DuQE5c8iQ8HtB
1EX+ECCq7zmJHIk0AEoXiQ97Mol0+fT3d6bVKTxdpbd9qubvLyyIW9WHpvypwFfS
W4lfZ2dGzLy4YF5GGbQBmzcGxgJ2c+3uq5JhO/Dsh5FgB5jAIruy6EWpWNyDw3sb
KP/Tv96+PfrAuWD5DoI7S+xTQotYVf6XJE6Z/5WMfij+wJhFTpSIj72SGpFFQnKI
kBrOHiaP3kON4SKDp7PbRVB448asrHiGGRU8ZTWJpYuRngyVbu6+t+0duKZ7OyxD
8W6DIXc9ZdmVtAzgX281oP7JWbyJJ7lI+q/3rhdKNFNhCw7BiB9nM7psBTrABQ4h
dSVo1+e1HSWv+ei7zz+RN2BRgnUVJXnK8WYSD6a9ZUW36Wc/gY9r6B2QEV/aO8dO
9QKRmj9FFR6ttPmo1xwjY4J37JIor3wtRWtoiZYKA1fS3pGGHxfUBPQGHNrNtgn8
O0Gb7Q8a1xy/3nfMe3UU2G5XEvBQ6890uibHlxXNN2PVNRx/ibcrb9YJIgG9DCOZ
67abay12rP5UBwSKVqVVTarx5o6qGlBYZIJ2yZC98OViwfdQ5baB7W8xjbuuy9Ub
K+Xe9kxax5kj4XGLOcdapvjsKuEKT7dIyntBHhpybTvfQhxaWOr9wO0MBKuCEtAb
dPGr4sGmBcowyB4q8gKsQNpgUtVNtHf3izMyHRhmMsBAdWVp3SOI+/wu7mbHmPKU
srp8lIHbNeCS7G4+0l4BYd3zDlFoqTAQP+ZVFPJKa3K/lVWOOPAWv5bgfICXuvVm
XbjMEQft52KvJR7yZjSkwk/v7OdTb5+pKnbaaIK+LphedTvLy7fXQMCOmiBJRxLL
4xj85EjIAlTxi603JhbsfchVDhpjbKG1ojYDVE3ckzE=
`protect END_PROTECTED
