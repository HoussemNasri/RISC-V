`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dfahYW5uWBGOJbfTJTTC91S7fNyP+2ojsiTwKZokXG1zThdM+kaZFk/JFruxaP8o
SafacwAzblTbEWyY9wQqHFFsqnqaSbvEFACrLUQg+EpJpATO4J3rwC1yK9UkTmZm
j184acTAcuPk3lLRgyQbAsDiUgPgdJulQJuAHGjOG0/1ls1MYD9M7Q0lCS6+vG3B
JIxMTMr42k1tLVSkbxj1CSWjwMbgcVFV89EZvwIh5B+Q/1jSeTr84hTh8+sYaCHZ
V3HF3fNrQz87YKMvACzGaCqLgA8COav8GYPQTX4L915XotQkNS5PiBLvJ/ExNHTU
M4ZesV4zb5obFAU8Wn68M/GReWWlHodGJ1WoLlSjUYM3HrGXjlZAoun3gFgZI7LD
`protect END_PROTECTED
