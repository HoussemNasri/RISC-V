`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/w17BThBY4rhhrM46xyUynnfNORr7JAFaiZ0jZ8WfvNaOuR7OznNg8GbvcOAROp
mcQIRNws3QPwfyf/9bjPEc4/EcAjpae5h1Q3YTUQSniTk6vpe7dVeL/FHXE1SBsR
yfv6HLG4qCNQBbvJDb1TAD0X++5Fx9kBSuBrKvues7/FLF9XyLtEIURaXvnN1485
Vme2zcGJZqJmW3A8z90iHdFxUmfVJRmEmE72XgynDsM5j8936Yky3pMVYKLTExDs
9CAfIxiYevQL+uwCrvpql/bAv5N9pM+3r0lb0ZnDeAHbrH04ZaandCKRZjWC2jHL
GASnxvGGlKh4jZ3WgMllbFvflQVZFNYDJELapP6IA4yI2euZ7I/g/bfaRIvu0QFQ
djdspUOurKrMcxAugyBlh3XfmxCNd69ecK/TDw9zkSlTM7cMdGEZuvH0Xe/qqb3L
PgDozzqiDH2CXV7UhK/pZi2O/zrai7gL+Eabud9gT/F+BR3NAIXh11D8KlmXm6mF
v/ceVCtwb/g1qxtPQB1NE8ZhpomqZn4fTXoYi4Q/AtYDSrzJlwpPjOedvbvC/Klz
n1rN32W0hLnUOsiyCAdPAUCm+77lcZTZbCbmL1KFZKn+LN9RqEEvWJ4IZXHhdXZl
bf34D4V4tNwGVQLZLl6TkO24URyoNZ1yRBtsZacMZ0mZ6kXiYMy9adDIAo78zZPN
bvfR6RdcTHdQgciyoAV7buJ/FCfA05/s3iuaPbY+/ycocmfdGDqwRQWZyDnNz1ve
ZPZjTq1edOZYEdzGkR2w4BKR95Mv8H+aJeWiz8xXMW+aQpRHDyEAaNU349TRga+M
yni0wS8RK512TnNqcOy5aUxENVx7BwqYgqDGNmagwxlABg6ITJyL6SgEBuaeX28F
Y0z3GlDDovlVarRnVO6AEmOibHuX8YzEHjtssGvXYzoM7EPI+1LqDWiboGC4k9Tr
F62R4SFEWj3OgudcbiNDusSrLBPLqYkQVldOxRWh1ruc8Sv2bNh9/Cy0TiCqcMDD
fq/LMEFnutzaHBxRfpEYNYt0pedpF6XRf1IblvROskRVxrPSaHrGkIX27xa1TdFu
bTD19aE/zBrjLtb5wDxYxk7u6Kf4v0+yo2yUePMqcnpJJ/CtpzAG3+nfGtWALqma
3uF70zLaiHqtEB+fE6TOyOfFyfl++U5+5ebr++21cJMquMb0XvO/3gzCk615WU5L
vrlrKMdqtLiH2i42Pj2K17ucZhCXmZebn4WzBrcbX6eqnNfUFx3qrpY9QNo7FuzT
oEIq7Z5R3QXW8F9nOabxhqplBkASrlNHDAVZAQQFJk422jgcN6cAhGSS422kb+7x
czdYaIBfpz3cPA5OzQIBpO5cNmfgj7olIWqbxoHUS+Nkow6NRiisPkIdJXix2Wz1
ncBr+sE69xU1CMbelCGhEcmktaczO6/AIMSLTjY2QR/K6rLw6sc/eFaIsOQFMJuI
9juf4NrzoXypBVQ9iUEDZIehlkH7YfF848nqFzSUS4ny5jAO/VvylDuuSFKJciNo
SAqFaTox8i8tbymBKTrEmX49djjRnqziBwDdX08wZT1p2H+y+G6zLxFaJ5aQmywK
jPPZ1sm6vQenHDFyw2xwqfK85CN+dgh4NabhWpPsUj/UBoRS5DyWgXzDHwUPKOLz
5gzv+Gy1kpjRdDP3hjX7GInjzyd8MsGzWR70VZmSrDb8lV59/8jNFV1NIpwpwcdg
R1ThoPvuhAyPivyP/BRQ1ZzY8t9EacLCOkZKnPt1/9kNQfx+GcSqgauA5SYaTCDX
fj9+5/dURW1w1F++2OsGZkFi7LoNdcbmfFBkwPhqpXXrRAUMzqkvB3sB4ekiiQE2
2priTmD7/D8HHgktjd8vlG0OLrpt1BQOxdE1IjW11gcKGnItGe7px1TpdFTBM0Se
SnLt+maRL3IBJ0yQe/eGtrqY5cDCYITczMl9ZhP02tP00L2uXLbPR/HsQWiipMhg
Il7dO0jvSoXkEzT/AJUibSDxhe2XSKakSNbXU1I7xlZQC56ln2/8UDSGolBqn08P
9b5S9AXYvDiIjoPB127Ns5EV3klXynUCertgTNUfILj2IZyi/UDyi/t8A0atkIQL
XLMqttLWR6/RJ2rDhqNebFEbcHRkGBrV64rtC95a8o5fdHuG+f3jl7MDWmUhZOum
EZu5CobUUeDuTqWNbmEN5oLuQ8cpkWQ+0lF/19WNQR99Hmzj1HQhfMcbEDKPKnBY
0r833oR4oPBFDYtXsmDgHQ+TZHndc2OlimiqU2hEjRe7RlDKM5Al1JU67SOTJj4K
4Epxtev9v8I4WjcEjU9cy38kHPlm76uKF6mL+wU2KY5EXFBXcsnAH54fq9zXcgqC
Y4HMFG3F8SsGu6xvjCuFsui+X3VUcQanFWc67CuZhtDsSH8B+qo4NIcSTDmlRtJX
L8N8Z9BEB5IA3G4hKZCUIcatSc+3B276po/OML8cu6mDhYeBAgWP4taHxOPpHQXj
2Y9nj2aGOQD9KP2XX1fI9xHwRmYKs0K+vyRRht3PhKlnr99C7kwl3NXtIlCVKd08
S9fApP9hyPH/6uP9Kwyr0OoeC3G4YosYbenm+j5J+t+RnrwjQrtBpYN8iUcM1FXb
w2y1kJ28fczRUi9AcJXWXiKq/dXpjnm2BA2sX/UKzLtWPO7TrMxwIvm6AulXdsPi
HcjbqZ+9DTRRi9S+q5gxnMEB0w1S/N8EiiIueLVtD8p8oBZS++RTV7AqQhVIFdWT
78FZIePySEaWtAySmcf/SUdc0p38L3v6C1MsSYnzaPljbVqXijHDrDz+FxrGY6Uz
fBna/Rnvp09z8iNvENhFd/25Rf3Kq+o7UyF9h/nCOK5+5wgVrfp5oTt5yW4tjrq5
hQQxBXG9VmsUQiGRD7McQOeGOEiePdQP9CIovi7rTqUZz710YEeK4UpDaitt9k5m
Y3wh/uVjap26lCAD+lFwH/OJrtdvJN85nxj3pyF+iXmRvP3qOeUDdtFdcd+7Zrcd
5YA+vGACxUQY07HLH5ZVZxFZ7K7++H8oYnY1vRonL/0vw8EOEcGDQa8TI9ph2AT8
OPLaxA3IbxhsjymLO6+mvij1T1QDWXT60rgLEzHaZleEXgaucqmUOgR6Rd3qqnmy
AQ1l7RAAS5TKqowJWRjjCjZ/8XYmC1ZzbWaYt/bIMx/DW9IyIiU/XGr0I97z2Mja
ZJ8x18C6KQCRPOMTXo/R9BHsfxJ3lX2XeQsADxV/BKaLgS1zvwpyvpskPTaaC7sW
Nd1FkBpT2WQOmIx1+dbRDlYnoFmYRovr5OMO3dKHslYLNAWjhUuDIuPKlrdvb++x
c+hmNhHFrIih3S+/dGBisv3GQ4C5zSVU/BMmuqJPK+lM93JZdOqcFbT1Lldl+WOl
DvWTYcoWdMCqvnblANgneaGDKnHjUjkdQa6hdwu0d4LEsh1CTeo75DBa4El3Ae61
0MUSBEnfbD69KW5foPCUypqbxNB4TiHeC6BPZmQdqQ1qM9pPbLydrqyLW2kkPp26
Wo/z29Xw8j4/dSDWz3RC25kvQCdfvUQnzlOmJiJ89xCoqw56lV9EaOOkbOzmH+hT
bnCzpXJFd5bOsC57SuFbAlOy9dSdzZ7EvzamMpnzPIVMiTd0+P7c+arMwH6v41uY
dcrmcScGuQWHMzbnlXikAFf4BhBtHKbY66AKhJ7Y1Zl+BXGkFnsrouWuMAEwRIvE
ZUxpEleal9xclJP5W2azTo71ITGhY1n+6W7MHi49bTvVBFdpBWxG9x4ZHY9XvQo2
yXH+vVmfvd7EtU1sQH42hJPW5seKVYhb5PINLQPhZpTiYZPtz1qcJVgqupFPX5F8
hWdo4vQ7RnHfWwQvZzrIDs/snhXMfW4P8etdeY3mVpSw4QsCncbQPoKLtjf4WKZL
WVPqisY3qFBhAKLxkMB7utCP9fKSmHEcA0HULzhlwTJUOIqWnMWM3Q32n0VwBFnz
hdR99MWTui5fmdn0AO3DoII5nwcatfk9UO42BZDrI2GzstJWYXSQTYMD2frb4kXm
HUFy9qNZjIvyonCU9jOHkc4Y470pO8j6qbDtuvpSWN4raQPSCVmMUoFUEryojEBS
ACIvPd1n9w0z//1u6uG/+1S5fvSkwNEWCkKwuaYl27S2BblCHXnOCofTs+DWm6fB
bETqek5SRCvhXbeC4NBzxFlYJPEg/wF3smly7K7P0br0yOIu/Du0nEKM4ejfaa+8
AJBGTXpCJ/P11XMrFldFEX1wCCoI37NhTIJn0E/RZWMkfqx5Y3IMsD1TuBQ9NI7q
bXMB86k5hZWh9OMKma1/cDl+5TqwgoScCGitw2v9JTHHH5zrmoTktdIkq/lvv+VG
es/cCAD/7TliYH2emqnND+95ATG7/uVt1DxpIXnmPIIwaUu6amXyk7+HCyUpP48s
56dZWguEXZCbLIU9iu7sXBBDXWhIQhkzFvxF6WlQyVRvEtswZzrtc+Mut2oj3JCA
6gCBVMvHF5uAwdzfdnzpHmVIkH8Y7KoDtqCr0MpLzYdb1Fzbu2tin2rHUY6Je42V
RnBDZszSnr+60b38s7etyoHIGio59v/bTO+d4phch6EiXLnwzkkOLDD2J8fetv3+
fGXFRqWmiQr88bcMI9AkHaUr8xwhQruZ8GYvTYhHMj1fqm+r4ApMWTo0jskhBxcJ
nx/zyJLFniMcC0KQKbNfNL+RcHTmyGMINiG/Pm75m3JcmvVEGtXbKbPTRv/3IKMw
kcMdgedKAyjnEOu8ntnS7QzmGmYxsPdl9QNKl4R+0TZg4nlgXfH2+NqPX2Xw9WfB
Ik/zSSB1gxgzhykCEAEQ1Kcyc/PMxviuDMEHhWfRhZ9Cefoa/Zgq1EdlWm8Rkl+0
77XR4f1QUvTpITCXXIel5s0oZ1bwKxmqfTvEVtsZ2dAJNDbLD2Mnc1kqXJSJgroL
yF5FceF8uus5+gumzE42bJfhV2og4bGAD1cI/8hqi9atx9Mro+09K7538ULscxlJ
QxwK0Y/VS6AyjkCHG2nxWk/S5S5Zq94JjAEIG2zgToAvSRR808Qe8/PRFnE3kNhx
q4FgegEAbb210WspBd5jHwxvZ4fdacGopAM0oup9yWZpqHZHZKqK1+ut77+csxtv
iRtIHJd8nWrwxojpH2S2yCCC+t36rK01+GM9bSkJoFOJ8VKj9bVVwzhhhpTjWvvo
jdvqFr7flm93AY638h4NK09P3J228JD7Q8dVwJbyOYBHMbAzNdEqEHL20QxdoOly
CPhXZR6TrnfPlQCcbvovWCHhaKfy6rhAOilark8rjVCq2IfByMf9BeopEoxDRXtR
SewAso2gds5G9e4XLOK5mZkTa31gJ70eOKM8kNyPgyNTb+ex71c5DV2kAZCJIHoh
1JJJ+1zB3ZGXJUuoyOfUGTVxLILCExO6DyAjfHCaVowAxiclyjymXHIMtVYOhHlI
ywVQvGPua5Jysb6zpEQbRHsuOSekVo89fP9qDa7RM+BAh622VCnm5sMRFlxqpmlw
3z94yifhqijkmsleaWgd35dmnP9ramHC9isz9seaaTVWMIT5cRHek09Expcv3fyP
U8bU179oS9pb81RJv55oEZAQmm978Ota81Uu9mI38+EcJOAT4qxz16knm/9z+1LT
VccnmKTEIboryreZ74l6sycrENgS+3q2clRSxXLO/hOALAgfmLBs7WM6g00q2ncu
AOrAp70KlqDY9KFQKmu8BqrbD0fWZ+tPe5aUJwd1mJCA4d+jtIRA2VOO5lAJrc0u
NyOkNaqWNhzQQV/J6vL/PRRTnkRuspz9ovOOO+c5vezMF40njVPKwvhHb9p5OGRJ
MXXQgtBK5FfL1T3pFljPWEYyAoJOkIXlrCA0fUMqi2jTvaXUO0YWyIBERTzty1nY
h3uIKHFXhZGVM88blGLSgWlZKx9mcVOybf6++Ofp4ELbRrabVHQ9EWZOP8XiuKy/
2uy7hrHKHUgSpwjhkM1PWMaomnBA2OWvXP+pRiYcLTg3KLGie7b4JXt14iuSmZCi
YUCHZdR3JHF3vSMh/V9djyHpjwsuPVSNRaj7IIdFRFDXWwKs2xIXvlJzi+bMnu85
dIlwT3X4Jzj39cgG5E+2/8u3GJ7vvst6azou4a3VKnfbZh3k9++tsxUCnXADqxRV
VVvDMSuWrOaDqsOnyEUG4PcBm6REDzsq3zOzg6VWHxfh2ICUgYelGCD0RA25FYXu
iStekeO8emuuLivt7mU7GTTNdARNmtr4U3fkKm1iE+dKHcAHG5CNu1j94IjjxHmJ
vy05me0RjUezJGv9Qyw1TPIAhvmHicm69pQAzrs7A3dWHZ1t3kDKpJAF7bKt6vNT
uVWd3d29iauOt3xx0uStAM8+MB3kAoUl8BzJhgFQ33EUN0ime3vgydouuS/KEwNx
BkkyAMTWzOF0eLSjcLW6/wmv4anBndb8HfX+V290+ZsN9rglFkPevbs9QNKj8E3c
PCuaIunXpJOBt/bNGX5BN07+nxsc15RGEeK+Vd6D+XV2vYQbDktBL4h7Qa416qFZ
dTKgvhzC4W+xMjQabi2LyJF3pY+wdMknCqTu43WJJUoyhhQulE7CrdVrGuguVzMr
7Ulf512P9SfWjLifPKWJ9K2tCs3It6G3SyssjtkQIs4LmyEWrOQYFqt6DFP2CPT3
LRmciCRy7mTDpk00oPeZZD5Y5e3NJAFIyE3UN6Npp3i8x7hncxfeUL7jm2jKDLnA
prS7T+X1V8kng0ZfiRKwmcDOUquQgLmj062mwhjWaKfAfxHF7rs+y5Bw+8eR522N
0QAYhEard353X3xW6x75pNprVaTKQ7fIiDbrrsXpyQzDQwBQaV61cjKO+p50t0pW
ZAn/KOJDvgm0b3tL8T1byltSR5tMbqniZRzFOPOOun0fytUmIetTWAT6lpzRA1hC
ZPe83tBh8CEA97lP7M9Mi7QWx1unE5As0rUdpLzkdtQIWl8G9zHu8i4LwfUFPGPb
PJ3IPSvtk6V7pGwvFB/x4gjr4ZGIHVMSYeKcYicztHnZbF2Jn7nuyvW7dnUyYTOY
BvoVHy4vnBPVpGx2gPBEwjZzQUvdS99fjE+CkjZCA8c39MSyRcj3414C8+nwM1Sf
/VmuFZrNRDf+gZFnZHYSiRt17VCBRnzkXlTlv4eqoDcTPx/peCjw9qubIj18IiwU
bLPwtPG0oK0tKt0pF7DICVWllziF3lJKUapDmldsDNsu0ZPstVMy8rYqmftd+Cgc
oqXzmWsOqoovWCwCxbDJWH6WN/dBlHz1y5oUS91kPvCgbG/hX1TAD0PvZexVMfFd
NVZLsgBSHvvLa0R+8Jp056Yplf+y7zE8Nq8nanUtC+UseQQyLWqgYGfgOvjJDmY7
vzyBWglRBTLXrVdgN0nJCSn7GVAO++8PTKh2b6NSsDCQiIJzCwOOlByoAXE2l6TO
s1f8L0Ki2c6XDzKFMD3Rqeaz0wX1SiqQqh8KYojELcgSXB23xtxRntqQRWgLdK0q
Tu+xywMRQFkuf1yUwD2kzq1PJ7T5RDNf04qaK+AxpwxP4Qzx4EuaAqOKN41ljJxX
+fn7Cs5ck3liqAyR3P311z6xMU57l4CWhSWCiH3ePRH8fgn30LVny4RCEZU8csSz
cvaMBgA/WWR4dxAWhtQNGmLvgRFb/nHKF9NJCGBzaLs0EKOyxwJs7ioKJNcuVKAi
0X0M9RllqTih88zE8JYj8uFwBOcV6+0aaMRC3KF9PeGG4LdYdkqJFPMdSv3IFE9c
RAAdbMxy7RcBoIxxllUDnVKj/SoFFHs8Ihh4SZJ9o9GXwhOgpe57Pu+FKojIFuR5
8UP8vKtkUp0G52Zmv3Xu+RXMvIRMEtVnXeWB9EiiGjp1pUEz+F33NwlJJCs4RouR
shgPHd+VAD5j6xzndkijTaPwzPtM7mi8SxAieFJQ5UwTLLd+qpsch5PfOohArjd+
tNLOJluZxo89aBvaQKU3f55bHJwG8D1ZZ3hQILi1YAyECNqSnmyL+fyN4D3/y+c/
PjL4s99j56hL9RMz1FE1fpdaQ3u3+Lz21qvJAiUBQHi/aGkPgb2uc89aEYKKOlah
SQm7RUfK7/IXfpq/LfLCQ+KkPUqkXaPORvzZW6Y+L+yAUrEWcSRwjUIgmkFPural
sV9n/IkyHPUTk9JACUIsVdkH5P0Xc/mPCBr51IL7n9h7u7J+xhUj7giDuW5DUjjm
WgGWzUz2GLqWlJwHk5dT3XjUKxANkc+w0gDDqxVXqkFuKr968wz270Sp8oBH5mMs
HjxTrgskxwenUN2NjqSO43rKd3KbdANciGmQ2SsGiaXOJM6IUIs9JRjsAnos2FPj
mJEp6Rii2JUV/HCNcmDvjkOtQn0QRvcFflwa3P82O5b0nk1/9t+NBdxaKqUIoqPh
A5g5szYahjWlF2/x27Sj2pw6GZ4rrpV9u1GGV+p9mGUpnSC7XBT5Y4UgHqea0DgN
8Yov1u4ZQGpyIQ+EkBSxqpkFrm9xSNMRFSB0JuCzsOnIGLvKiKS/6u1Wv3TmKsL9
n/bZsfYnxEB66Vfx7ej1CH4H49bXpO3C1zedYeiRlbjudv0Rg2MRkT8C/iNhMkr7
ip+Fsr+LHQ7K78AqhG+x9qgdo7paHE69sfPj3bElirQuPF+futd5p6sTtUctn3Hh
4epSKStoxSO5rmA7BJGAfJuO59el29tl80sPEd7dstnQiD470FDwWkQIUWScSXbz
2lk1pO7n/AiUFnTiIfe5RBiy2+QbyscdRgPiZs6F1tq0XyyFhq4Rt9QNQ3BC8F0/
quDxrk2Z/MoHxKIah7BP1kkITL/5cKbPB/V1dccJJtbAX7ynJ2/xpeuzxgIZz2+F
WwZNuLBXkr0mdB4LSRx6L0UJ5duocdH7rh4uWS/5R4HttgRHHk6tCfjjld+DkQq6
aLeMFtfVpFTV4aIOBFXfLKtFouakWyQZAN5jMHvsK2wXsablzkXvBT5QPTY797ip
FxbR/TSr/nhcZr06/TtXeRtGovYAuFuObrvcPZnmVmcI9c/iLK6r2aeku1Y8rO6S
ES1QNTIujKPltEMbczYu3JNcvCdCX9OPrel0ujSyANLVb3JkO4QJO5xgsT/vbWQV
SM5O3NKnfjmlnroiEhoEvzPa8Q9ACjZ8cmsgKi93TI4xKZLYMn3TxIifFdFM6r9t
B4qvVC8GbtNzEXkSisURaMgtxHeZ3TRH1V0e61rrAP6W9FaMK6PgmONkQdMF8SkW
bO+HpvBcd4htefurhdIJegXhA4HtkiysTd9+uC/BA6IVjjyMDLYIITYgp2GL0e0x
xfXF7xzxw+3vUfxibSoH3NIBaVN6muzYDtgWUu3IAYx42jFrNXld6lrK+nljl81E
CRoyZCqngfdROAv//JL4DzH8mtqetpoCAWX7tkXCV7g7RvAUk6bdPnl0dvZ7A1cZ
6mfhTX22XS249QgliYeZ69bGzLjIOE4dCgB2IoodGupuFBhj8dL9W6GZT+ABgQ0y
rJFpGdbmsk7sOpmosrB9pOc5aRH1gCSKo1ZE5XA3RRpcXm5MMFSVYY+/Bypac8i6
n926oMP1h8cwv8GOcjNZvESyRhpmWP2P7S65GH36WfFWfHOtTwCfiHf/jaMaYxN9
VRqF18Q+CQhaP4nOKeA6IQ6DRXP8g4IbAoWcZLxdtJ1FEAa3VkFrIisKBtiXKqdp
LUeHvJBHxIecPv0lFarAhiNa1OnGrGxfyVk6hfwETMVNl+H8Wfo3ps158pp2Vip2
rQA5lIa3unFJ8OUoQ9cI51skmB2sc6+mDiIiYrUTSIMP164k/mDXQ7UeZ2LBIkpc
ECRTb6I1CCHMg0LWw6NveYa41YIx5WEZtzdzPt0rzrSWN9IsweslnKgkj+8M3Oyt
Re+dT7m1CX9ql86oaoio9Up3TpSYi1V4Wu2DuzIA/KX2x2szUezOxGfoXfpEzfuu
xQR3Q4jqI4YnUW+MyHSPlmAvsGdWQ1JYjAtnjb9y+WDb17GNpzEHHJ8fApQSG3vs
NqYD+elJy7VnHjQc1QIXIvTadT6aa7ucJoZ6uRQr0NL0ngV6WquFj0mOXxcNqNGv
IyGjCpbQ0W9RXOSV5NRsWey4JDw+BV665EsFYNwYJWNBKY3XrBpzJjgVrcyC5jse
JBhaspzHQ743aeKDvtgzu+JXyhcv3rHBejdRI4WuSverVYhMx9HLqtO6S4InOZF8
vTiTZLVbZTrxBiXecTFqGLXcGQ10iKyYGVuQbIcQ4Hek20ayt5OG9aKhtAdIOYjz
rUXjcdDysDUEnx6A6Xgli1iCItY94OUhFnM2n100vZrIYOF9icogd92BDHXG/2cn
EuAfWVw+Oi3tMksUzksPr0ycUMENc5a24RgEgzXPPP6SGqbsMMm2BEpfmDv97Ja/
HNqQlWW1MrSwwVEZAUFX3gycMuoIlMx3kNjjYobHgDBQUyoj4LWsyB96AIGXt/Hq
MpZBK5QLUij4yL5DR8+ak8dlAl5RoBzufj89Lev74pBhQMPtS2OUGHZMjEhJXh9q
4y1oIl4fb9Unu1jhTpgR+9CjSwcH8kEpnjll5rfS3eXfdFh75+XNeCXbGLdibxTS
5TOln+V0798YnDFBdPcNqpbqJdE8k8IpzRZ6+SAQnh7MKiJiGHXk3e0hA6bOEih2
xx8pYUS6fAsgTK+Vkgvt2aoAMBzyfzQwxBKk/ZSyQWhiW7i7LG6CuDoPfF6TLE/v
OXdaGeXdx4+5g58ULFVF9yNNxl5Ni5MTVrMYLlYC9HEA+AdQqAkWhhBIp6uXQaeD
fhDtsUZvNrClKgMzYBjk2nZjuQt0Tf8ukSkWcc+vH6ZpstxZVfnE8qoPl1MJm+Ps
qv7HVFJ9temdUexJvYW/lmGVZj+n5wr3LMAGbhXtS/580CNzZsLE8tWwVSLNRbPI
AC6Xm8cyp8GKQcBr32hl9GMN54rl7hZAfV9XcjQ4XTJPcfP7tJyniR2nUwjosSy+
zNURGLpeLwqcblPgGVKmAASkYpXGb9qFXw/F5r5SkckrmqOb7tO/3Ozs8iXruJo3
RlW04kcuNWTdSS99xnWRtzDlYXV1LlsSyZuHtLMlFssUXTcZS9QY4Shbo6f1+lOT
EhQycl0d8PoPIaEpo64c2xm5BhXe37AVqwPqgVs/tjFn9g+F21/gECN9DT9nqp3k
wvrwXsb8Q1Ymz7E6uxhSbWK50AZzvTxi1J0NfTkKHtgUW7d3suhtubVs6K96l0Ib
rjDv6Luvla7pBnO2KkvkdlLTk4LVnITUfZ37VQPe+Wi4Qvw4vfSF75XmCzhxmAtZ
BVxI0+DZwo7vGZnBwJpG3+49LQBImRxQRzc8ZDGSieyOEaPKLyziUmFwPcIpSyC3
HtXmcH5kI+lckLqRa4Hibo47eDk2X8RXxU3gECUn+7bU1zajMat00MpMlDwdgh6p
1AU+5zYUtKK0PAXCqU1F0MgjftAFXYbU0IeZy9j9cfL9YKV4o8JR4CdsarjT4q/U
cYfFYcXq9LGr0MZw6gByDuOHUKlcZ2y6/wcZKz7HKAMTLhHcwcROtR2/rfaZe8QH
4hHh327hsNIFIz5lIo/unS3eVpEcKD6CxjpSuPA1oZbye/1dJPnkMYhNLh5hcJjb
KKg6RI48ICWaIQ4fPTCizuwfztcMxLDspwBhl3OLhCpshSrCcPgNV4m0pPTrqyVq
TG90v9UwnW8ixJ0HzjcSIBCOroNP37/0AhZaOd5tFjCLTAJvCuo+hUrelgYwuZpw
dRszc660Pb7TZ67w8QttwtiIezATJ9qjhkH3DJ92St+khfYyBN8Pv/r543hmcKlS
o0HZvtvURqyaVNYmzThulAzxAlp9Kzr+wkCZO3FohmkXU7vMr8ApjFyyViNjIsGt
ucda0TizCKd4cdnCnFTnyHOcllXxqhjDGQ7C5rFC2iYn5+Ir1iMEPWAVtDFXN70T
+w7tNzvRLqTACwN8o9340iC90WgX9SHGZWmeJX8pkciUTdEJlKEyKL95BqLFe8mo
N9kFbj1HD2p9K1BgpRu7FeHrrlYcSsynNsG9NKzwcAdHh9ef4YwB7U5qAU90fdjX
x8E/Q4VMFGH/a/lQ+cJeVgoLtFq4QGC74Mvk5QEyUnPAOrM1GQwa5HTNNkAK39BS
HxX1iGWqtqofDI1DG/wpdrbSfKlmkOWbLslok8gxXW5QnuF2aq3pMIxit5O8bW5/
zqAnJTOOTuT68UZvJlWK7du6V3zWTEnvYBY8PUUEHGGrBxZSGddI2UNsZOlVQQam
gfUateYaGmouZ5CT1XYrLFTKklCvXYZqYepS6IyTERBLQVaXBTsX2D2Z35jdmE9c
NwaXpkBsZCXaV/hX40BezXeidTrWbDTQGnLws+Nk/PMcRV2XdrYvROpgG8J/zDK7
98eSdrHDhV/Hc/5tC6OxAdfQAB5ofajJqYHgdRml1X792rckSOCweuD+GuhqvhGM
kuOBx3UHG4P7ozDz+o2RPdCW7fSSon2jCFCdGXVZzpH0YCQaXpS/qDUp49r7Q57t
Ht+Qhpvlbuxb6Olm8nBVBtS4xRRM6lKzxY0YsFNQIi0akQ7piy3O1ylsHusVh34L
qkc3NguWE4ekhYx7Jm6JXxGMVjUyh+HwczeAjEnXNc4DiVp0kuSTf3cZhf771dL+
ilY8zwZdple74MlEh5q0wdxbHZ+JSootmBbK0J06c/ilNPrIg5GO6KP43ogIjUDq
dbcIzARnOOdF79AixmboBn3/r98iW0fb9Sp9ggMJlKhCDOV+H3joojmsenAtOlXN
TIxhb6F/wO8ShraGmkgA7gEmns4BsJFcyK3sefg1RkKx/hmt3N0JErac5RQlIvT4
Vm+D7lnGmKWh8TzgPByY8msqjXHUc8yKOrkBNv5dtONbDMI0O+ZugwMXefZskC1q
MuJ0LHZjNSxVIjdWcMYOTwURtZPlzKOP/xjlYDZG7MDi15gHmpE2pqNqOVg4uo15
PWcK0Zh4HyKodK/CR1MdGRtzKllhNiuXlf61aO2ZWgFN6Wru5rCzZyU73SHB1K6i
l0ucFMgn1IYr9HGp21redk+AklnYMWmS+7s0z2xTiwlDecNXjfF/9HQaTWpVA1yb
TT3i8H3GgomuTmek5Zh+Kwvp0fdRRbsYiFpNi5tzeKORErnis2m3UR2kBeh1Wj/N
s5dwLemUKjVvcfCfaTzFvjk0s2h1agXvEkTGiGb6lruQ3WYCAyGydrAeAbPeGAan
pl8Lt+WuKkPm1vuGeV5uPjyvK/J8gq+f5bKBK1B0soX/cD9jI4OF2ICZHto7jEMH
VBxJD+wHeboedOA70ExY0DY6aVxJmUs7CBrM5Ik7ZHNCJ7/HXWEMLN8z+T3T6QSE
VX3FyFINJDv0JKwirYgyhvwQfajmTcS/pRiJLAq6wsJ9uFuggPZ9Wwru+HxkIVHk
Er4I3YDM4zF2Nkk09p1gf85YwISeeVTsJa6RiJiCTOEpSkIDjsyShI+VAObpFMbh
PHXZZNF5BUei2X8xmrNjqfSdpxaGO6coi87HK7SdvDoNR8KRnOwDpMZiorGY7Uxj
nBt0zonbAs6TN2ij4Qc8LpkmkPNKu8bShLYijtjWkgSBILR2QJy5JfeuYu78knpX
btbv+IVrJLjvA4EreHE9Aj+X17efRWdg+6QRdsUH9OuyfH97hWdVLp2iB40kpFsB
OleTjDVGSr4DT9zUxqxoXGETkPni/jzR3amd+tBKOxXyi0+A1JFg1jJbXVlzgVPt
+qUt9Ybduz34pfsFwxQrRzbGbyOIZXEettVXhO1jYxODr/5wthm10bfWKXBn4p/5
pMorLvoW5jX34HjdAeZU/NKSkDP0oI/2SxXGGeW0blRxgAi0wwxU71FgZ3bgpBt7
AANCJfGItm7WAwNI/gpCIsuH49W1cLPhUsDDA+uxRmlR358gYAOhIhpQZNfd0ZBf
oWnLeCs+L8/6lDmG9Kde9QOiAAlVEGM0bV1lBB+fbPbmUM8abHQwG4Oc4xUpjzhJ
OY/7H0Vxd6Ae2RoaoJbsNGhXm//ShEvb2G7ze5Mk6qF5gJI7fYZPROoC7PqhW7h3
XnDSQYu5NlZfH6r3XvlyHzi3UbxP4ezjQv0khy7VGC7zE5IP7lxVBIPiA0/neAXJ
JdRGAUtIYwZPza5bL7xhgaFXoO5TfZstrfGPvCS7G2Kdm9gd4PnX4XuZATCLvHMD
2LJfgiN7zQcLC6F8eXvZXV94FN7rgkKbtlklIDvMRW7sR4haauo/cQ6rtK9H6uq7
cvdSKe5+UpaR5jsU0hClj+26ALqGFCoo2c3EBk6xuG1FBQyu4FPB200sq5uhQ/NH
qxejV0BGr/GHcdpE19669eloYlkmB0uibbjSa0pqD6jmvDzI67Phbagr1W1mQ6tl
ye+QC6s18flyJKkj46fpyzR9SlO9inVZIo4bmJH6AsVbMgqm/J4p18OJVvNsjtDB
awsPN0U26LeqZAiatGmEM5W3NOvwOLnm169QYvcKPt8ow99NPRsmLxBCdjpn7tDt
OmyUry6W1GdGKuxXWK04u38qJ1bLtbm0HWy1hFZnX5S2eA1Z1tDkRSGDfzPTOGk0
OR2Ft1mNpM/JDPwXKJ68uzV0yhpogvcb0KMQcohYVRWSFb2DEkrtgaolkl8kBp3+
oowdTODzQjPXzz9lFvuOlMzw2ZhfDG1f8HULHbdq1zIsrNjLT7iQBzM0Hn0MjpZk
UXnokOByTu3+UQZYd7boP0GI0OUaT3GVyuKJY4vva5uXSeK8uK+be+Pv/9s9l6qE
a/R1ulOxndgJ1afM1j7hqtpTfc+iTYUpGKvMIiuU4davSlrnsFu09Cd7IAKWDICx
HYVI6uErrjL1OyhEjBsKNNv8uPbduV2YfYmQ7A1nmzmuv4IEk1E4YOaXoRSp8mVY
flDq6tbPjlaOFjJIsv9xkeRugS6bc+BQBN9QNDtnxLTdynnllinAvCuPjVCrtDtH
LCVH9spOHq5WT/VtEAPQZFs+ulhWZxp6GJrZoKI402D1mOEaijMdxHCJvMaLdd9X
8sWFuOq6eqFsB4lFmhamKagE7i7I4PTIQKqcs+SMdozyVuO+03nm2DVf9FFiYfDR
GpU/3ZVXFzAsajf0x8oYRIeOBCSVh0OXckgSMy+mxUjN1vrghWUtvjK2TzSFGMEg
Vf7kVv4ZpaRQ3Lcm+G6peV/gjJTbH59AvnmJlfrMvpTcwDvgCLyK59+JSjH3W5mb
HHZSPMYj+9HcspcPrkOBOieayr7aEVgyPo7BegIREG34Qy1QQYaLgUysCPkoLZCD
e2H0dCYlnScsbj9wCS1jvlLy+LfNqnB1jTAxbxybbs20kPIeAk6TQMVyN3wtHQuF
CjQe+OzVwObiqfRa+lZiFcabm3O8iffSsDZg280gbG3yvSKl9kMYpsYFtTUYqZ55
y3vJyuKNn6hggD6tPn03H6PB9qXuLwGs4863Gl5PRb/gXxw7fMuAtalRr9WeKLem
q0UGk4Jcm42pzqnwYUR/fwlmmiMVmeG3iKUyKJIRM+aH0MhFreEZ2NGgsJ5LFpyS
lTc/utY3TjJhOtMV7AyZBC/VaJoKKWlxJgk8uzpdfWnJ22EHYmwSCDHVnSoomDYe
mQmwUGjoDJ/gAUNataPq03V1zZMSQ5wqioXQpZ9JYwgCJJawWG5DjvVttnuzMCSP
AYhznmy7JaFVDxS/8u9wlsEnCZEKwSx9hL9GBtJ/Vh4fE0u0W07b6AV4MYAnODGw
fRn3igBjnaum5kuPxx2y179n9sFKXl6JsTkl2t1l1C/5s2CTVLzImY5IfZMtRh8t
h0YfPYaiNGMROrXbknEX6Dr7D9uG0a2ZPY3SpRs9TjXLhCYxS/+3HxRFPhDKnKVx
ikX5CnuOz2rsKrE2vPwm1tRpH+Qj5cLn+9GwCkYRwJTaXyuArO7ktTJf5/M+ztmO
wgBkR0UpajLa+sWoXKIqPdky54t2utcs6lrWdpWWxemBYDNPjFQM/jh/TBlUyzBK
FvTQeqYYwUy/CJpNc/+JRT9nd9k7wit4MD+bK0e1VHk6icFn2KsP+qardsWmL+a+
pJILFJNoPH9VY5qDf2Err6LWLZFv9MmcIzq130eyYBYf6FMhwrkEqk70maIAWbUl
pxBvKoLMWPFUZ1HNIkwgZ/7PBYi0XMT62QqrgOckuAh9f3bpQ8p+4FOWE1GUABkn
RD+JgDRRr0+R4NkWdBXAW2Xgwej5A4ShHpOnSkZswsYZkDy/T6BpaXPIFGvsXs3r
m4yE73mJAGXNiOKFojZKroY7LrTED0u0yGpHPoVAv3PjQ64NdYS0+dGJck+/6MbQ
g0bg9Qh3mVhdNBiWgnsR1QFab03W+8lXDJaaB0JepnV8gDyRTdOpHIxqoFR9TGMN
Q8xxyE9sNy1ZDUCkEZXq9uDOvDFAc11KrfYWOdIyleoAn9lV9s6Xvv3uI+CDmx2K
8vXv6mRH+b3yCXkted+4SjS5JsVLJoSRq+V+2Hece768o1BLTtzcG4Xy1PUfOSqP
84eaz5aQut3QbO0WyktnbWXoFib2VnK6hiYtCuez+qFb18/xYGrraS2kCanlwZ52
CagXgqsgHImXpwwE/Fv3eX9v99UvN6EewexZd0a+se3NRIUiiipBwV3jzvXF7U56
zBhSIkkAosM8wCtKWvtHtrGh81CJ/OfCTL5wlbGFDMQwG5QWcCqklBi3KvtJ8r6R
1W7HporGs3nGrq66ZDFTS3/bHX3R3UEO5CxFxGGHBh76QDoIyJ37LeahzHlfZMk5
oQsbFUN0z1uu+YCwcOz72bds5sYDN6Z4EPb0HQv9CK3QZtQgFonu3BHk9xTcgAfB
PLRAOeOe/5IXoC8LLzox0GQGEJdnnpvrrqPwyAbGvxOg8KsI6QojasSxtLbfdRDb
LsGtsUXx/UuBbijXjjOXEdhRVm+kde8hsyXT5yNqwuh5rfoTN7HedWEvxrZ+OAZT
2KmVVmr9zV5KD8Rv4stJBDL6G3wpYgktyOkYIKg04vNq/N1E+g5fqiF624/4CaxN
r78kXrRg/UN22v84idSJ8l7vjaixyO/SXZqz0V0sxl2VvYg52IyKg/B06k7TJaE2
SRj7hqjWOGyvxLty0GqPkH6xlxM8K/P5eXAYqB68RZNr26He54x6dv3t3ER868Sp
4X2kU1/hpFfdJN+1BJev5QIWUWqU6e7RavnjrkElxUKUbWL3M3DlxeCUBWZ5hp/1
WLhIJ++eXyHJQ9Z5zBkL76uzqMvFqJE5UKMZb+1Ii5c++Htc4fhKGmkELxpwY4M9
i8i9gY/7C2Q64CFQYc8O7AqtZr3y1lgCk/nGwqxchUO/fAwMRS0hnyeIEu9GeSPw
XbsHjcDRaukWAustTTRjV/oDcP9AkU/ndiiWrmYOdx7GJQoy8H+u/EyNRBWBlprT
mQtuFZNEOTc1VmRjT6RSTW3TiV+sjlQ3YOIqix4hcF72LriTSL8/+/dQDaEnj5Oy
/Pa1m4R7By+Un+ZdRGEaBSL9i2hsgDMIub2En7stVA860+bW35mmCeMBl4dKjP3v
3+dcwsd68mHXsfmZkRxFx9sN9nlUP8m7qvAn78YqpRQ6zMV5B9EdvaeQP9Z9SJN8
oL38kcaXSqvU2l4Nu/ZI//0R9/W/xk6QIBadhG6aAaopd/7CfdAeLVuD0brzkTH+
lJyOMB61pLyuyexh6r5jLEQYgkhjy63xDPNEKzUEyQStcFL24YV+ayRoZTPvz2/f
4YNcjKs2157zhBtiNYrbsHc+rXFfkOpBaKKJo5jyLkUoZGhLw8yXGh/KmYd6IjIH
II2/S/c39jZ2ogtfmDkhXE3qJAE9n9esrrwJbigH2t4wm8dngXdmFQ2i5fuRZARW
/BdoAs2FW2rHXRIbHsyezluNc7Y2fq8o5qd9zEiSlKrnhWseH/nPHQUW+6WLnNF8
AkQNbFpPHo/Kezh4DNZO5VsH5OkrnU1TLInjbn8syMzh9RdvRbOePzOmR6GuBSoR
rN5M9klHVq+nG0+YEpGQ56l7EmLy4H7ufIBZpHmJF9mwGpzJUlbGcjJgfPwNCX29
uE5y6RfjgwHyZxbRM3y3VfWc46mg4mxClk4kwswWhfva7mVc6SupVvqMtJdFjYzs
Arm9lTCFGGtjqipWXrJyIqToqFzc/f1/DFvg9aOgNutEKEfOLGZutC3vDW4tYUvF
2U0SAGgR1lUD4xs5QCuafAcgW0glXGoanIaLmV8B2K5OGcL5yTERK9XftJ3Nb1ix
DddtYtBHQ8fcqQVRvuC/Kc7WZebVY6z1swBmh9ydNRfiOghXSRdwIjzSPUZZjosg
pN3qOblM8/KHrj9LWqASFj5iWAdAaGCvkqsLeu9VoL+MynmPBbGTxmZfI9hvtzPi
wCVJ2i/LUqbR3Dj81qgTpjSwgQd5uzi43BPn2eq/XqYBVgUNk08LfgCyD8H9sIbH
ToulMjyQ1VQAcwjHWAerQt1yDcFEFj1hrHjvu2HHuAgj0JHAkKKB757kTCYIV/XE
qAX80rRLE24jWdIJIJYgQKoZSmGiuI9RK9TkSYXOA4ARtg7PmoeAX+amxnUdh1g0
v7kEVJzzhjlB9I3c/YhoLioqTiFsu0qByoDVs3BJYZfWsNzfcYECkru4I+THLHxb
08zlvVeZp4gUXISs4ftbPmQxhu47tn0noRGUoUIkuoY3ogd8ZFhx+hNdTU8klX/E
UpPR92VxcxsSnyWJCcbm6E5Z43HdIZfMc+oVrKHJFonhGr6jebh3Znq6dCcOyPfk
SsWMQMgQh2a+8gCnZ2bsMCJX39SebQbOk1gMsZrQZML64S4+FRkNgCCHUdA2Fsk/
I0gZekHu1tP1xniDlkeHBoKzukEq8B4rheyW75e8Vk8lc1aWBgTvV2l7h+aWpEvu
iKWk9O0YiPynjnOr48wCZA8JAn7ATfn6jkh5jWbegHsM/g+l7Jaj0XL0Rmh+rqxh
WAQFYRHy125JZ2j8Yk47Vq+g0JDq+ABn7EF+y8o0O3nEXShukwsP87jD2Xssho0J
jWQwt3RuPV8VlnNLugs49V2FW3nY9KL6an4iUaYd+opuAGA2MjPw0eU7RSpUZesv
iNGTjJp/olPB24dFXt5kkMe6QcY7Iu+fNQGGfp3SrINvquHG7Nu4b2JwfixfOt2K
tfLbRKNs0bFDXc8A+xPYA+yvDlvcemte5llH/POEML/k14PSa7DOxaTNPSNtx11x
pF/RVGZpIfc0/7nETf7C0mscuk49PD4FP5+VWbg8qk8gdCmGGukM/6a0wn4acdHU
w+JnNW+TwuhdHh0+U3HuDLWziZTzzdI79QOdNBuH8n6h4MZfEL08F6yv+UIDwh4k
qHaRdNNRQIcKVYBiQYDHetL9x2MX/HPznpmnrhf9LhHDIbWB5e2ibtK+wn+vOTrY
BS5W9f5BR4qzQiEm2/hE2Ql2bSVFM4Estc6SP3abke9tQPs4PKbFmGvnCnuAkmwl
NiwTlNC06UoNhYVkmT3eGCWDfWQxJrgKUdDgep7LE1RNuQWBZzHUeuZdhuKXU0Rc
DMRwIQTBuYp1gH2GhxXk3K7suZQYE2mRtS5Tbuc/HH+RcNoWT+tH4KIi6yKsgHp3
pYWEp/SBycdApeLWDrm2ZiuvRkovahzrdSf7NHrRQ6cgXlVnK1caEVq4ra6XXShR
xjLO4Jc60jAaL9fjThu83Er9KyKz+C+tZQZlW6XesCSPLQ+psgKvfXXe7gnZQLyL
be4yUXWNg0ElQI22Zrhvp7rsRYcWT/l8ffb8LFguNExbUrhv/2Y2T8vUlVky/pSY
pOnMaNmO6/Q1nki1Bj6uC2NaZmjOLmOUGmyuWp1g8/D2o5W+jY84w4+0bz5zRJpf
Zdy7EbVtzOl6h/LSgA43/+DYBEqua9LgdJkmznr2oklRueYHh5SLpeNFjiL2GdG+
hKVP051abqZp9uvkMrkBIhsPAZVbRMaBiX7DNEmQn0glqflMKnss+VtrgL/bYd4B
RMjkOIY2QwFn4E+mU4Pczg/+14T2xFTohg3Z1KIhatwER618jU/0ESjxkA1tuSpz
yI0efCD1SfcoAjkYxk6J7L+GelXVnn4u12Ax1RbnC8PZ9hs7p/naiN6jMevWqbZa
QrmDV2awyKjnDsxEkvVPNa/MG3OizkGU35cQ5x2OFx3owpnKG2ft7HIPLzCw8v7o
UT4ArGSA1I/h2qbEtjlM0PuDRFlK5CWwszYoUothXRe8WY6KX5681A5k5Wc31ARB
r/M2ijD2lmzuZnlga5Z7Xp8/duiX+hFQhlzbEL3BfhYxlxYdHgXXxkApC7jqx9U7
mZPVDPv0976PSNE+J2n7x4pFsqZ0N03KVCggqifQ7x8ES7vT6+dYTin97EJGQYmA
6SraYYv414R1x/4G1GP82JIbWhbedxwnlG4Q+TngUJ8kahbTHotV7CVDWYvNP+cf
ZFwcuPOTMgRMdWYdjANdAQUafj4gwGVn9M43f+SchdjaesA9/Sbwo6bT1mVWyp+N
XqN7awxvftJNpCgmLIqfZRr7uFdiw52Py7CsANY0WRGm9HKwDsv3yRCA1YOvszhM
gbM7MLu4yNMFjfUsLXzhcBTxZ+PbIlK+BZAmjC3sKt0P/PxMAY79BOlTiVq7SEbK
FJBkKs0q8WOFGkCSKxBakTrU4b62l/lrY1Wt9ZdFCPLsPhxYXUeI0ebXv3jfiXto
cuPe47GYQd7j22v7928iLXmezft5eMZmJKmgw38LqDrMC+g93S8Qa27izx4Ybo4/
dOmhmRQw0eEq+1xdvfCZipgE6bPYLnOYPpeGDrfHJ9Vef6WceA6MhHM3VTdcaPOf
rBPnO0uF6t2+nXZZlRpupwqFg5w0p6Fi6Cwxd+mfiDpJVyp18yqeoOVwtWH9m+FI
1ZSxuICB/t8EqAGunK2HhRgJHZoaKMKAUUwTa5hRZIw280T42XBF5dxa4Xec0A5B
XMsWbrBB+rgvdkfyFIUm7n/Q/0PJctdMRnuGEONEfqpQL89R5SlwhpuuytO5bG8F
MBVOwhIMRogk1T+1f2UqZ4k7YmAeZHM/6FLSo4EAvMyAQRbw8PfyCYPlA3tnTG5/
DR81ZN/cAm5YZOOvJ4vKeb5M60o4R+XmLN/rbwfXcfvZfJZsPJUaGNEA2zZjRxCP
IvfWGdq/4waVvv+LZjW28crl99JyVsicKEDzFQ5ddm72e7qNm6QW6iBXraWlLhbG
WYKmxEmKBqup1u+ksNhrGXZDDfGsWoOT1TRkicjZg/7g+F2CrSqTl805eMdbk87N
Z+QEYoVXwopPHDE23hsyTnsxMc0MjaK7Bt7mPUCeMekBe4t6ZU6ZkJbnR/VvtOT6
hQZhw188WcPh8cBJvmroafxAPE0+ZrpfjJoQaf8XyKo5j00yxaGpJAnWUN8zW0IZ
f138bDcD6s6pTJhNizeUwjZmuK45Gv5he6GM28EMQ5t05Dhbb4905dOfOvEbgKd6
hh4skoAeipQLOgQRDbejX5B8mVLnkBiUN/SB/8AnGg5ulcOXcOz2zFRMTXmzyWmt
rDw7n8eXSuTqFAlkOeV3jAJSil+dsVTtQlhA3zlJxp6Hhq4zWM/ScvTOB23eAQMw
8vgx0UOLGBdMP+l6Qpgcvfw8uDBRG4cfkzk9HpSrUGe8JpwzkHHWzXSO4cIu/CX7
70E4VHJ12hqLUeq3YonVgfmO4t+kqqCax+jxFAo682CQc8lS6TTlxVMnJ0bRo2SN
OV5grQF/KmFwdwq9qYE4PG1/nSpmyqumDCfas/Gypr57afsec8hOedosaREznSbN
MINJVg4D1BTFoeDq4zo7BiQf1otUDGsk5NmaUUSJPchIw4vgd7LLRZqimVMY+sHo
4XsgDxB22b4EOCNXs6x3mcYgZo+xw5XM1zOQE3IlPnwdoDWZREI2KGIcXLf6yOAX
jGm4biZ/2Qvp/xj2xBrfdkC2GOGoi7xzWNb2syaXWzaoCJBKTJ1mVRvilqpkpCHt
XSgKTChSuI+tZkMquyev7NNo2RyLEFWwKZdc5n9+yTJN02j7FKcoj1ztTEIq+f+L
J3WvNudx0ckcU8v4GueSXQs9QnxHE1mCYKgkag8d001YZABYqY8NlCgvOfBf7w5E
a1TalsSo0MTXZ0+d/TQT2qfkcp9U+YOhy4GHnljgng7C3wouGgsqvBqJE9AyR6Lt
zTtoSU4OpgziUymtRTa0E/zUzawmCEe4EGQnTI/1iRwb4UjxmK3JqJVYAmUW/RLL
IDo8FKwGfG0HTwgZSGDCgkeBt6PW53+lebW/54wmG9tZXw5PaWly8AKSuo1TPjNl
CHiqxorWM3Eyz2eNy+tFJrBeyxmB0w+R9qCgNfDDWPX5EDqKi/0UUCA1PFrjjfr+
fe4uy220+M6olERXih9cbecqfjrGHydG24+H85GJs+FTvlgPtI/Ie5o+mHqchNGf
xDMa4ICyr40MEDRYMvXvTDVZySx792cWkmQc9+URBeRITf5MsINp5ML6whJK946T
b+CXnkkPz2iFROy7X3ClWOhKYph5ITM2xVAleMU9AlNxhsSsFjpujn+HfnVFMrpe
KvcE1vFG4nEyQ6dhB0PyytfASmWxnbrVYbwHbxWrwsjcjoC+JZeoajI4BsVUhxQ2
40jxgaHkC4aZCB9w+Ntg6Uz5w4UX5O4O3AnbGTH5B1yrZlTP3IopvYRQNJ6nd5pp
xnufP29B6NSoXjisQqS6sMZkY7eDkUsP/1ADcBjC9IGdAOyqikwWEZixkaahHnEX
TzXXxjtSKqP0oNpkwN7Ibe6kah4b6VksN9ML6qiTaGnoCJ5nTH7xeN7apkNK+zbL
bl0ao/dqQlJssHNsEZVZEsPpoG9eknb1TA5g91awKVt86jV8dpVoSQZl8vYuie5/
kvwduG5Vpthi55ZNh51asvM/cmYScjqIT0bgOyjwmG548T1fL2v2jMb6G4TCpYlw
d4tqleWo61r6wJYaVlHh1nxC+uX6j947eAZopQ9izVYWGgkR03wbs1Byk3V7bw2p
NEw6M0Ee6MLSIOSrEm7IRj7wzl0jiR6473G4Ludfc+DgwfzhtgcI6ycjNDzXa5V8
zQoBarIcOMr+5atWzhkNaiK4eKRj3Sx+JWxHI4iSw8NvPUpXfq/hsOo+Kh2Hstun
0M2ELxLkN5SCJrvHyan9debzRvsHuoDQYrsD48NKpZzRwrWBvZpn7JxM7ZfNou9M
+Lv9rg7zEqvbQlqBmxEGUt70BxO8d53YTq6KnDy3PNylaAgXcnNDVY4DOVOTOgg6
rOx67qmegXu66FFOlga1gurFKaF03LX2vy7/4xC7ywCFeaqm8jp3KOWmGQpbL5QM
bl1SAtuisJCI/TotAGUjef/0GtRKPv3278GUkksB4JstoYMULgb03yg787BidvLm
YFa2VqqvvDsWmPw2D9G8P8L3yVc/IdSUXuaoGtCAQb2wSBrlmTqN2NrAO4JfG/ME
ALlsrigGsA4Kt2EYiafjWFlD0G8nl8++suUA9BiKNcVp1gvk7GhkOuwgFzF0CCis
Q1NVUnQ+UAqj6sq07aZaukloJ5dW/epQcKNNyChFnq0fOQRA8SB4lSIvkFHEm3bZ
LUDAdMVhb5mJ05hbOJ4wxB9/PGElSi4cyrb0iuL4mlr9CbIP1hJt9n/LRkYdIaIX
jhWcCzUyvCXfjc/g0c4jGz+w8mLN6rb2ST0lXJ+k0wCo++lm+4w/m4q0TmVtdbBF
IBBT+Y5YaY7MbH7DtBAyUat9igvV77cUKohOYyyE+UbQseS3ZmzjgP5gdC3tc3BT
0Ab/FcMkrEIWueLG4DbFr38jNbaSivCArOcvJiw/OfWLj70d6wr1Rf73aU98skaU
ZIdzRXg8nRumHkdwshB1/jJ7svmf6e52bnSASwIInhQjAzYg5YrJtHDr8Ro7mnSW
tWaqc5ae1lVVPkvVysxIIX/nn0XkARWBn3T6dpD4D675myltZwPHsK358DC6Zxo7
GfVMawOhqMq3knJs/SASfms4+zaKEDU7QGL0nrSlh2mNSaUn9pkPC291mc45843O
9CZzaykuJZMED/tc+XBONf1rP5z9D0A5jy47j8YaqwXvzHmSxkImdjaCaWCfmeSU
eJntJNvM3de+vkr8pr3RdZL95M79CjeNthJJlLATBUwfpnKvv4ePGIFrsEio8LHv
OUbB8Ar0WArE/18zxVCB4xZuKlBplqtw4EUvAt6plMTG7s8JxYkLGK50KdI3KEmt
Ep4ys7o4VZon0stkcrgqFQKBoXi6m0u9UEgPRAN2pAGbGmq0q5mToasz8tfMQtcw
BAMuiWLDNI55pmSJAJv1r+E6vvA/LnJtWvNj0ELEK/DwuWV62ghgfD8x1lPZyNe9
+wzIXdTiaxqH+r4dxaLA5OntG6PdFpGw2HD4RaAwaul8fSkDk+kZNTLP3At7nNKG
w+fP3EdbCsD0y9WE4Q+ZBcpstDdHnj/vRdCi1GeyowL1xFIW+c+MPQlyn3qgdVZ4
i75nP9Al96bh5mC/0or0EiwegnsafWe5/vzAlqRCLAEbfvTiKK50Y6qAZH1uJuQS
ERMfQNyR1PxF8OjgArlv/6Ko2vxJE/elsrJRxumOkD8o+wuX8ke2z66+1F67w7wP
Ex8HWdIayrXTZVAiPC63JztRLJteHiCnoJ/rRZf3MbbJQ1W4/q7YqApByBWsiw/L
YYZY9xu0fOI7NS+PHfSl74eRhxbOb9z/O4dMVmtv1ams1UHNbzosuszq5qubpr2m
YHEfErpB+7sll8KtNpyY08YqAzI2HObJjkC9t7RZrNsOK8KIa6UZLrZjL7Ei5f++
METin6Qk2oHFEagL/2DT45geIpTwTvzyWQXZq8drt8wmk3LzKRrIBag1nVi34Dzu
mc3U/0UaitpA/zk9xJSJXN/ATFGq05PeruM5wz0QU/sge7es/7lrsMVPqmeu4YFQ
Rwjmtzb7TeVcY5IuRYEsJPtAG+lYI6hNifqrBjUlDV1KxmoON0Zwa/QnRf0pfXc9
6ujkfHQRpRBdEkR/FAUkviFCRgkT2nq+KHFBrEZfsrtaAOz1YroNGye6ACvKJe5w
ccQMdudBM2lxCrgSokS+iO2SUG9klAbGQtn+doNxQVzGLs6m2ccmFmAJK8omic4z
/we6Fo91vOUYMsgjQUy1YzUMzs7jdvuqk3rRBjBrT6tDnWjFV0aVhuPoxg1z1qZp
F4hM0YtgX4MVbNzt+U46rQL3aOY/1rz4y+pTL2hppCq6e2is6bqONNUtTIXnLGsO
0m1v1TaeosSK3W3j7sgXpBogxDiCKaVTXSTual7irzXpaDNGrIFfmJvgJuq8GVcc
srYBH/qQKhT7tFyRi0bKAsmzq0dvNoShy/pMTflWYkEhuYyuDUWLSGWrgdV0dhJL
hf4534mW9st673L/UHmkH9DKp0rGmkRL0UIQl2P/KLVAmeB7RjHnzWIRs4Jk46CM
mJGXVJJRBWZ4M9HGxIN/aLbToIXq1hdnH+bsz6RkxslPeMgjVsS3/B8ctdFwLUY0
ma9ESoo9bDpI7jmjGzqYlzK7BNS2uaOfixso2Jcvy77elnA1dt26z381K/T7uTsh
qWYs7nbJIMjTSGD4ZBxQL7twED5zJyzp1aYrvsLvYdjK6ZofkyRAMT0ALZPd5hOl
dnbo6Mplit82kzI08n3h2r0HX58fYssSPJoXBtRN32E5+y9aVD7B7R1btm9Qif8j
eVsjT0QUixO/pVieb3bQzuOOwIoIKEtnPfMPDTSJkUkC1sqp8MzXlNo1r7DQs16L
aCeXW53hUTFsIfkP9Xd9OjYoIn+Ac0Ecukb46mp/h8M5r7MB2cRBQcIB/XE27rye
WlZ5sDtJTV3pmgWeOSylHkJdq0alza1WGbGrChnzehxYjaKyj+UJNKme7t5Cy151
7ksFSegLQVM4EJYWOeDBLulouiNhCGYuHfPIDlCRw47GO/MiFENAV4sZ/W35pazI
HdDNLvZwmEQa/kDoMjYwHpBFyNNEZtMbNOegAUQBodX8/DT9SM20Vw+M+HOdV9hf
Yc4xcqegeJgNBo+TBQcg19rWW592aZPIL/nHhofhOzbwRY5jsVAEM5FbFLAPA2Jf
B5F+RA0xKl0VpOnKFhqepBhxuEP3peZ9w0uA6UTkBmpwUfEb7EIJrgQBZNekQ1LP
e01h4ooieGYQTUb7PIkKQ5NCo5jHNF38ujFFEWITpq3JxHKUOumByEY+/BahyTc1
1mrl4jRIsE/Go3GcD+neCGtwTh2DPzw8Ph3s5cCJiGVp6ONOShl0Dw1ZWoBk7aOs
YhlaQ1DD3Nrh/y7am9INdrt6UwBq3yTupIZotBQlUdYxpoD6xBLoXg82bMwAfP0n
5KXSvvau3yucSLv0qCzQ0VjWqeyVcTElEgMBcJMLQeI+zF3Nzrsa0OHqggu3+C+A
J1i30rttoDjOz6Majhmkj0IpJHMYc7oDvZYC9Egm29KHtAF9P7Whc8gJ/ORm/9jJ
kmCsSS33ETFVCdYD0g5MJs4Q4DPrqe/V3Gijz30ylClTrVHCyMmw+Ic4v0Qcjs00
IuVO9san8M0uxyltdqXcTl4MnnXvTwpo9phk1+dMpq4Z1HQTnMb3DD3cDYO516eL
6wAJItBoeBQo96f4xqEZlPYX7BQR6ZR2eRv9DPRCJ7moWoVZolC2beiaNWM0XpFK
2EPSPiTKLkVgjW0QQUz1TA/0hZfgAaUuyuWi2IbEbnoSQ2cHXWGNiraahZMstnW+
gr5vSXp5iB+f2TAFbTDvmxEdsQpgPuQ43SNzQ92tzaknZ4bCqsY4245ibZxbdmor
lFeyuW+Vyj4IXmmuZx3T+zJIiJ9iEqTonk6YNkRVvhygC6hES/fMmV5Iv76UfEAR
0JTmVko2G9wR2qJjMU7m7wTglmUS/DWyNEjEPeI7JXfCLfkN08eAEP2jPQveJJFp
XBoEuAtUJFx90WXEkwBG91xpzfYx+DP+Uz177RzaRubMdRqi3Bw5ftq1IdffS6Uk
Ge/0jQsN7Ho/Uuoc3qDUWPWxh4SxiR/NVksbXaCvyCF1kDv8LtDVEDGPtffLP0/z
WwxksSSNMxWPZdFhAOOwQLrerFYbpjJD0IWwJ+VOoi7g3H4lgzWLc0fBabBcs/r1
oUdayMx+NG7AiMQnkRUjpoYzRVz5pJoUPqPr6NjP3JLg4cBOfNddHCtHrSRKU3VP
Wgl7DcnAXVXityjnmqJqz0YJHOByVsyCM6/oon7irGpivnt3TdfyDgrysTRiK/SN
yCO8jS5JCFf0VLWWxrXBChGC1AS84a9X/dtcq3Z89eD1EOSi8KERkeM1Mqvgl/qD
Tj+79RK+mBw3luWXJNQCASJW9QGUWUQL39ZHWZdMyzJXdnRVZK/Z9ziWy46KxAl2
jbXIEmzM5n0NIzITMI5LS4tfmxcny/UZKFysdYyPEEHPmLD0IoN04Tll7PnYS8UZ
rVg+8Q5LN04DrETQKUStk9QOTzOUiL2Z22pPQRyJT3wnDAtNTaUXhaQpKITx343t
ch+wqta4sgw82awoJKKbAWIKR55gBMk6goInhcPbiCQCk7hBW2mV8xOHlnm38QnE
53c6Lfb16ii7m4+de88yPuOlrvRh7fTDGJh/rhua7Ks8pHklBgWuP2is/Qv6OSdj
AH7xEIWTU8rpL0vQoalw1lKTjrneBxHte1N2O0DKS6h/xVsaBd6DcO+B7ITNy4vO
jGCb8qKfBUalkmEXOhWiIe18dmjOs5yOe8jmWpQYwDvyqzNIEvaL0vXMVprXxiTB
Njf0vZ/XCc93evlcjyBCi8jTKxpxhlv0GLWTE4Cw/ZUIySUFfa53RfpCTAboJ0Bb
CPZp5EZ+QuXY7P3+jM+7uTAXLH1KNVwYn++DP6a6GaDeII9NqTF/keziQbIkfLT3
EjTkGmIPmdBXk1rpuJ/2qOZ+ta95ccRMdtXWCydvfNDKKbKb39DGKaP0B1n5Tu5N
uMpsnYsTj572vB2oHTUly7LtIBpp99/n5PCI6xrQG9wHhj60kK1MNN/EhpKPGl2Q
PxAA/GAZJlRA9NCwPoS3UTlm0Q/ET3ZG6N0eH4ilVoWyk5rlFurztjmBOaNVsSxN
pYn4O0OvU8ah64oaxy8GFqvyRUJ4dHHrrptpeGQ5kL3aBfGyITIPkkrU9nrmauCE
HkT71h11VLR4zDbFmyv+ZUgjlOS1kQG4r+9oI2xTVwcoeDWVmxLruzBDb6r50UG8
EL8wDoLiiVpEiYZJ7hRgUToGHzXt4IfSuaIFTIWaSmBNE4/gKRdmX68fKhuPXuJN
kO4LJBiPiOFoNaGpqWcJP8OhCfMnirwnledzESvoUPTncMlsN7Bu/hYogo5xbbPn
4zrBwvjKiqdbgSzIlPPGCXdXCSUFlAhHWhQSuVbcnbAw5ZFFruBYrh1t4XfZKgtt
XGTp6L/lIvxq2M5OkcokYUq6r38ctBzexRo7ITI6a483xKoCYV7bOoyCA08ClfEc
QqrSeSMWsOumTowxFjARKeq/Px8MafD7YLxuzQvLKIUNFykvoBOUy4FWIVvJKwxx
VyZRu0oRPwmkKvwREWv2+V6lhZkIWSII+ATFtMRrs4daweTkoMIfXyGT9o/CGBoX
TM+0mgnArW0a8/bGiQaYOTQFOoasu2wkYnfybkM5OJvB2cgIlxw7I7t55iSwEtk8
pz1Qf08yN6QpzdDDTvUYREIYsyQuIUGMJ1iipIWtz/w1QNdvClURApDFewzbCU4N
XSUQyON4ajm4u13hS893/7lTCYzCOYuVxUiJGh0dEH4FflEioD1vtVQ84o4nB3qn
qmyL0WxRGA5vpvp0Ou5I5UjcZ3+0FHV/2i+vxGQU7KK7XAReWOXRT2HYxahf1Pmz
JiONBFgJZ1HAET8ehi90AZAWChll6TH9gmdNT9pGXwTYGm2iL5UHIuLYw7zExrFU
st3t6ibHLXcDy8E6Ne6jpW1gUsSFGG4cZG6lYPMCd+rZGSP4py8cUxtFR95uaIjv
obvLoLOLyERxSw/rBZP0C5IOvse3LBDv0g+qJY+8RVzVp9TSxTrmssWlzVZ1JjOZ
xftq52pcRh7u0pmRFa3qzGmiXt55LFikSvzpjPBqvIZsnFb16ohWD+yJPctS80qQ
TJaxuUwbxky3HOO69ZK5AHVbSpsKwBzSHa05gzR/soyyRAmhBntsysrgJJz9+eW0
PV5QYQArpl13e7dk6lFZdNfsfdn2ElhP2Mer3HpgUDzJYh4hm5uf4jtiGXnATT5w
l1O4GZDhkv0dx5e+m7yrHP3wzI3JK+KN3U3TcFdvonaYNO//HjsAleKhzcL48d3z
Vj8sKaats0I42KPU+pHfygfOxRoL7F7tUftX7RC9cXv2RdlzdcZvLu1nxU9/ZeTp
4a0bgts6U3l/B44vO1I8L0wwhjoD5A4ouMHLPAdtiS2SPQ5/69itrYIIIPTDXb6e
s2wwoSwZpgV+2QL9NARnpjZu80/demikxvgfLxKo9lUxq5FKGQDYpW29Nbt/Eudx
kjak/pGNw8MxPADEE58xxNLJb9TGGmwKaGFDp2ngMFwAy4Iq3C6DwbYG6vKJsafR
dbSd+3TUIM0hhE9H3jvYTNDYChmnh7VyH41y0EJuH5sy5VvO3Z2ymIvhBnl68jdb
wjlSy5DI5ACZC3BWLeYDNPD14hZmwrSGJqsLm5J0BY4+DbZd1ZZ44Py/40EXxhdn
D5atvzb4wiaWPllP2IcNEMJqE9xKunhpE3PF2nIjsgXuKe4e8AIlw4JfQCOjOHZo
xxs2CZrbn3BlLNupaTCJZOaabtAIC+ty1QS1JXfRTE3H1G9F/c0OrDCiIhLm0U/W
MuevVIEXEEXnQS9k3YQzJOARkwAvr+MsmIrYpIbxVZvw2tg0E6NyW+NE80u5ztDF
YT1kS2ZWTOHgjaYIZVCaJfZYzp1Yq6W+gRACJONwkK3seC+kvRlbKACo3PR7uNMu
Sgcz4qnLYEi6fBbPIgBc0Adwp88/YQtCO809BlfGp8akRQt8GC7NuOvfH4yBqVvg
hM9jzLtk8hBaBPhpFcZJsAyYN11uVU/r6p8MXTBMRfu7C/fyBRdqteEBNs5eePZ4
xe+GPZbAXoGNjqQ4QDr9a0Q0+cbKcew/exQIljLKmOm8ujadiVKksDCZ0Bdzs0RH
xaySC1UTgK+NMBQRoYLAvlMFsL2BrRlYexXl94Mwx74+g9mfjkbuSl3cacLnIzxC
eknPeRrRbB+ozHfeevhTU3JmPN2UNIu9+B5wCmMeajbd+iw0r2Us/mnJPaRgQ1pc
9sN/F8+MwCspVQKgV2nyXv9xo8AAeXcRkuyIk0uZIc2KdiTCzEdMKLoLqmAybTA+
cOQnY11qza4UmnyJ4P5T2B5Z5zj+bFKhW/SWmn2OpmKRmaVNxWtHi1L+nwQEsZLe
COc1AZBsHU7dmdyG5weoqJSbaJsWOSaleMQih/5MAyNSc+BZ/Nv863DTsuYtJdLF
voziBxq+i7Zz70g2yVt3zCVGvQbb7aeY1WyS1UWeVP4xj+mcyRTrsV4ep/09plK6
ssA7WdSCDP4EekTpih13V9apfnxjK94t+HkhreCL0RwiOPMSLNXcIadPNSDu4jvo
ku2pD2bpngJ4x1p5udzx4qrum+rhBm/h28ekGyB42Ah7/vn7laL7xEE5asQF+MTq
O8spxnNsES7MbyKcyMmfdN2e3hILjTFk9ZD2NSV1LjkeodBwdP3eqzHkZX92dWiP
u3lQj52SCGr2Wrav/RQdi581LpHy5Fy3fQxWNB56i5cKLxS8lsPmE/h5gJxNzEZr
5ac3TgpdzSP1pqGGrXz4WgHySpSv4Sr7yTO5QEPHpelxzraYfiXSsG/J2//81+sI
au6GAwhDvgl5xNscj0OFn7AAIaylkspV8hsMZVthmGuB5d/umnJ/4aonzDx8En6i
pKkCfPN7TI6ausLWQlhLYNStMeFVirDRSqRqcfhLv1LpE3Vh/pDULbgxFhjwzoYZ
0sqwVkU+tWb6VkLLZswbsZGJGIEcwGymOozgnlgnHifgJeOBJAK9S226mi8LU6vT
ts6rBAxgCeTPqhbJsXz4JKFbJiBqSVm3Nx3fdJCkPfc1iwyCYU+vwb0Kpv6hOFff
8w2+3hdN5InTq/R7JMuUtt9Df8ha5g786gnsBDY25NrGp3i/7YJoPWcV54HEK9k1
+uFs8fx8HkbuH8mvfoFk/8nkiM5tClT5GbKg5+WPM9efeP/zk+8fh0zRCTgO1u1T
qJQ7kTcMfYor3egv+83MdMtjT200cYRJtwLrnsSppIGrYofbfYe3Rq/NRMVoFKGR
O0Q2qbIagVNQkoF5Z8XiyL0gRKji3GbyYiBOkx1oXSYES7INYa13nrCNInrM+LJC
O05owVtlfjCdyvSUD7tNT2YZ+uslGfBqWAunJU9k41VLfuSe4SAElI6Elv/FDd92
n1wyRNhy3w/8K9zwXFeC2bWEO9eSndfb7SV1wAi85S6KRV0ozKjuRIsmg5tjDPmi
rjme9Jzvrb0D1LAE4Pq5Hwom5qF/sCcMT5EYRK09DxuQ5H1MzXWm95Imwk575H0S
w8obtxe+cvqKl1g4tVuIkCa9Zud1gQLunMsea5TgRwhNL4QWeQUBokLbzuKk4MLN
zwTIkNjd8WpQq2YO9lvNMvB+cxKn1ObWTkhbGKlL2v7kyR8Prcdmhs1xbDo+1Tf+
BPrkFeVABBsp2ahvUTPdXDVyMKQUZZ6Sj875aNl3+Co3aRcXW9zmfSYif50atdVz
gFTOjE7+WT9TMiPuNpApmDEhM2V0azhdf6mwTrOsaF8V5iKWFXfWao0LejEr2fL6
Rnet02r1AsKhB+kjOtvOQW6yyuey2z9Pe1WQgIurO795DuUou0XCEE6yD392mmxc
BL3fh7wbF1JuTOGSTE02BT7s3+L1+S/T0W1c46eQ0OgNUg8pOVOET0VAMDHxK+Tw
d8cljL2O4wFxAdrNwIEZAIv9pQ3GU1Il0KkJkIqa+Ix+6ew/NH49wH0ivJH5Hv+h
fFcYPSQZ3yd8j5/ZgsrN7QqJpQnyt2yAFaA5CJQ/kp81UU/k15TGTcARbiESEAjR
FWrqY9hRLu7GFUWbFtNKv50GfPC101Pf6BNwyyydAhPA2HVuny47N6NhPVDj8Rud
UXXTDKRMCNTSonjQ7Tm8IPIIJ+caqczmD1+eB6sjjEsz3t2IMME/wqXwtVeyGeVE
1OBeBuwRDrZ4MjLd1tCJQ39JzD5Mwnrp6xtjao4cMB7hh70ur83NVQAp8NKP9fq1
7yUYYna4BX2rZqMhHr9egkArxG4YzRaNOl7VJFjpWAy2Rknp41T4Z/kLg8NYnzzB
s9j1GC9/cH3pY2Ucvq29psImtRQ6x5dgm7L4MpSbe3HJuPf6QdWhH3CuyyxNKK8F
d/ZwnYDoFijtlAry9w2NLE9PqtuM18tTIC7Xs+fciP15CnIaAf8ucsssnAQ7FrJN
bUe6MUYhXCwSxtvw6Bd/LYApNNxYz58eBy+fwo5sUhO6KKpBjj/Tp3lvQ4ljhIWs
reLFY9eGHmDC/UQ/tlNYtMcMHKRy4w3hBhgJuKUY86p9XrgKs0m5YtHw1mgEOUvG
tJcudalRPMhcc6NGgpBpjShG3vBv1e7oR1+94b5DetiWaWNGX1X4ENNtRzevMCcv
c5Z+5zl0+ziYhIMHwGkCnuFuI71gC8Cqt1L8osE3hfvALMw8OMRUZxLcwkDD4l7P
+GVX4Dgy48Cu3VoKKzftDwUyCRX2VzCEtl/kbPtvhnrNGNEbyjZEdRhsDpxhF1Bc
V3QdQ9oH96bSPzYv1YDOTL0ofyoNa74Ub7hMHiPT/V12ZTbY5TlZhvN8MGy/6XmI
PD+fG4tIbPmzhfzfTUv/EWoDX2D9SpTLny68WPZt7wBSPSa5oS184gNjWE71S//8
pWi6Xhg54RREiEAg+5hUyMuhU4ho7O5mcvyIoNv6Sw68og2UWxVUSFWOMeaeiL9l
vpyrfFrVZUTgvN1v++Tu7ImSZGuwJhRRd7eZRJWaF9xqMZK15UTqZWT4s/QG5hTC
E7HNpBfCKswavvV7ENODZ81mF7Hr/Zkc9momLNg3DnJzQjNUrghG+v7OAl6kvp5e
lliEB2J74r5XYkSQFJ8FUZQHuCCt8800Hh+8SIXAPG0fsWYlVpCspHScwhKlzSaE
BI2N5t//Ekf9PK5QOq57d5vgJzbVaYQ/MM2z3VmowbAF6f/cL/kWTatrh2U/J4nD
Cp1c9aYKR01ORRXt9lJ18dF9UexaHO5m0KWbKmKrB3hn+LiJEEBg9TzNlo/LssR/
zVdyyvRO5+WNbSWBOoVk6Tu6vx5azHxJ1wyjbxpFYNlXN5D5T72gjZ/PRvFd1XgE
TOxVNRMPzTt2PpjEAGyo8OO8K8jRmAi2CsOojIlyqHJWgJbBjN3O/JH/IF3HRlIn
kk07hEY7fsgMvuhAk2XF9fl5/vzPZzKjK+mlrVhaXJZ5Jbp53s34eig0ZdcNvzpk
0D6dyJSlIrLtSDvmen+l5VueInZ6+vG/8KL+Ri2ngv51C18qqPV2Y/3quGvtmKJ+
2aDIf86qp2sNsIXu9W6L5h6mUh9wnG61SxdRUP5rIuverol3dPmyqF6lVqTMzuHw
IaDLZHDKcDxUbIR2HYUT3JqIfxEj9X3PXfml404eaRuaKRhXBbJBlD6B3SpKsAYL
gAl2kbbUgVxdWLcKEdrWsWgMlEyleJTzGhRmkIf+Pn3DQw94Au7WZSZt8v04HnLq
oyfb6KMB0g0GwM02ODTRPwNl5IMUmyg/Kzlg48negFeG4XIuUMzBTr/VO5wyS0wk
tQFKOHx8/fXJU3qzw7CspcTq9lDqqnHJsk4ll7EYhrdKsEITrDOwR7wzwS9+vR3/
e2qpPvcvZ+uhXsbV75gG8gb/EM1Gbxl5+H3c22jB9IzHVShJAMzpOaR5z2y9W3Mm
+ODXyq2+y7WGczKacqYSwLwqJUbp1PfxR/mlXfnaZ7wWDHSESQMJ+MQTRI2rYmZ0
vVxDjV8KG8VywKC9NcZit8yHev7mI3W3RJG5W6pu6VR5SecafKQassJBK/0HADtq
AdOyCOHTfBCINgwIeLgn0h/RmHoZePbJqv9db4L6PQR+Wsuqh3g7Td3NWbz1YKuj
DNeZVL/nFPzebTECDkOzxswjoQk6AJA4nDl/QQplr0LeeHcBNXXnRKvANZxmfRvI
rGDjo0cD8T5J9fShq0c2ADSYbXt50P58HWCnlvE79zg1y5pOqCGp6+ASoBYyodam
+uRvBvnlGQEJu4bX6csUE4suHdjh98QovCXRDI2whDffvVIWZLbxOrwcy0ysgXXx
R0UO7vc5hhXjITvSf860FgxBV66Cy2/yezbYY+bwds/VIXNhZUN+YxZnkoWimgUh
aGR2K3sV7JsDb+CBsdjNl3q+AEGbmQVknlCpX9/ubzIZGM3LptrzQubeKK1OHvei
EjAqtlo1kyjg55/6ugXdFWtthlwZMa7hzk9KIPte6me99GToJoPy3q3JgsbDEij6
HauPn/6SHy2Pg4bqbedBcw/vIwQ+/NCf7DQ4SmtaukdNcN9hBvwd6BFbPVhYWpU4
EbEMp6zeUEXGr6EeefuWQyGlTe/nz+iTnPXzUOkuKA2t+WXqs6niGb/O9R4Q5D19
V0N1/o7UhnsmrWBBzPPLhoBl7UJ58ICSol3rKWeo0GTLQJH47fH45mdN3RGRt1M+
IoPm8RX5tHGo+Tlee8n4y/a7OMGDBubmpRrFlzmUVlNgjbp2HwgLcbQ7g9IBQiOD
5QQH+YmALUC0t1EJBEo5gxQwl/PRfBtQPu1dI9trmqI0Fd35upX8RMkvbK8E7l3U
q3dZASSGOLfyYzrbXfmInEahAEk5+3zaY+7g7MeUZ10xPCQrN0yNGuAYSdIg/Ehc
oHWQidnAnLx7u1VjhqbH0I1vYP1xQWnqOatyuFpkq+5UIVB2yNhhl2j7MCZicUOI
fTX4KTJa5AXGmrHcaQ3V9UJmE6FUxDdGogyU9LWkcmi4imxbtewNkK4olf4cYlg8
aKfJvtZBG/lQkIGLTj6Xim7DcNlHPnf2kTJtmLr2Jm7TGYnfagHQ+337tgF5zm/8
EVkBiOxllqEF8juH8CQ1bqY/LVIAIjW9ml2ND2m1Tw48temTd4wQhKtSd+NPaJse
Kvczn4nLFpAvcVA/N4DAGZ+QmvqhDTQ8i/UVEcFmwgJlKaq6Xfcpkfwa0+QYxcCu
VIJo8AySFH1Wm1DG7CAsulUe2h9bPGsGdmwsO95pXQ5uaIXlGXYK9DDOAFbYPdPo
tAEYp1m+ZYLUF9xzd79D0ppdL/FnZNRHXgTW+h117tlrP9zcdYspigwDsQr9XxIt
cVShLicI1tVtyDGzAwCbMDV1DuYZXL2Y+BLxdGY3Sz2eu7O5q6yAatcAVx7TYA0f
CXSlVY2nzPvu6FfG27FYLvZbLWrpziOGwJVjtUknEeuUlyCbUTBMm9opAbdOSqEy
MtvSmGR2QJ3C1etHF4fhd0/9Q69LVXtB5qY3xL2x7qhB9R/IGc7jMt1qJXjg2RnF
a2W89gzaoxEi2ppdQ6299pqyA1zK8Rolxy9NK1fmL/s8mANvdpkIDJb+EszY4yRp
Lus59TBs8Vd1wrGS4UEL8f9brgByYnjQs8clTQDR/m06XTc/eDD1XAmxCb0NLx+3
Y1559MIkWUDQiSWPq7gt5PiaHWpiz+eqgw4X8ahy33GPN9yxctVsPB/g0mmPdK1V
muVsZqkpVpLYt07j99I+7Vf3LLy6r6CqnMwkw8GwpUvDxD8f1Xz2K3ZbZJYGKJx/
fd6h8UqI4Q4mz8t7JVr5AGDmh4HbJttRxVBbhUMrc+OpR2vyN0FDokznmlK30E1m
aZhxmS9w4Ne/0KzHYjPeq774dAsPzSl/BYxTMROWN5+a8YBDY9lekqmbt/jj/8vK
lszkw1W6+GqrgjCHD/CjaE5NdHKyJDVz8ixv+IU0riNP3eiehY6t2gt7qhYb8uaa
XZTfY3+GeY8BPe2A1CpxiHqlvvXZa6sGpf9J4TpTQy5mEcVvQ4pGoZ1sQU0X/tbx
lhaqoO+MXg+udbH12QK/tWrgqVTE+8zh+WIhEXTruOilPt2EyZnYHxigz5q2O21M
cWzh8dktNlXmTq/8p9rrKheblucfcnNkBU+z8mz8/hRQOChWnowmBT2Hxvrw4gRd
Pr4o2OEANRWVbQgsVpTCo981kI/wl8+Hp0xU8H+hQT2cZe9aYsQU+hLSpAJTsgcV
/TAxqc56OLncYxVBTNClbAfjako82e5k6KFpe3sJ4JTTkTvAzoy/V+Em8TCto2VO
O6E/ItjO0MHWbTSzYwx1F9D1Ec32sPswv5Khcr8GJwZaO7ZsRD6iQa7EYAzSS3CM
+QxmPRWW2TX0/S9KkzahDzwGMnOk4i7d6aNr8xI8+SXaVSOwraHEMSAIRpLkFl5p
8ljhjBeN5zhjLfZK+yhz2Wn7+QnpR2mU0NvEQSReWUxlZMVRP28CBZNLy2Taxr9z
aheHM8QuXOfFJIUAgEKGyBsXaxzTyuVhvhWYHRUdgFqyGwGRX3ELTxz+l9dErgHF
ujJmCTaB4zTdCtcGOfnoeKqzNzcSkpNFbWJbL9d8cq9ttWQQSxSU3X2SZ7Gw6mcW
32TJcbQL14OoIZZw1Zebt2IKAMr2LoNSNqfL8d6oI+wUrhSgZUnGXE4wJRqRIyFj
B65hYKbwoMh/o2wX8VG+51jS0A0e747s9w3QX0A6RhqOs9KzWr9oYFFAcUJ9ok6Z
8dwhu+llL80J9Nn0bPX+z7WyGCRIOsU2T/WU3Vvujf9PDz3/FR+DpELY+Lr00eC7
bsRnZnQnYGeVmImMqkjYVSawEOZvUlSyztlR01ooaBrLpx1GNP2RqRo5IDiLQLhb
EwEct7D3NhcnQtyn7JvJ7KcTJycysxdnvo1GaWTs6RSRDAl4JDYWhl6AE1AYGCFC
2VdDHuvKJ2nsleSd08jdPfOB6NYMXoox7iodbR0SiKQe8jXQIkKzDs26w6JhEnU9
gtAmQrjuTDFo8jQRXytN/1HNBGWmrVMRgYrtmISEOEPT31PuqqeOmn/JjCZOwxbM
kPYC3mx7Ydtq1RAw0ZPLtaB2YvmMwV6GnPAecoCjBFR/Du2ONINaL/i+C+VAyojJ
vxXgAtroyWDwdnNqyHefDYWbXFEBGhNl4n5lrdqZTOkPGpif0VeOqB+NS/opjkXF
pKlR4uB0zeyhYd0O/Df5okrW77RYnAfWirR8/ekKyWB33tWs6Hj/fheetwW01q3U
JXC2eED8NbdRJhGV+K0XMH8ORdIwQ3Nu6EvWBq1Y7/QcT+2jColMdcT6JrjwqVI+
KN3dBpB00VNo7kPvZcLqd7fU/f2X/gqmeBX+vsWztK3PLHWVQlY7pBz878r7JXhD
1af0ii1/g2GjgoWaboeXbMHuSndfwTR44ypVEVgjNYWi0ouzcEiFzKQqsSPHAgkj
IzZ2272fqqQt2uBZ9gXSUgefwUUtk9fswWTDqKBn6yxqDxi1ubPCLq5uXcoW3wZb
hhX7w+ZN3eqmBUKlE8kTMTPHqry9+DWgsi+mt7eMP3nSpXNUAoN63nYnvTlqy5LU
RBPLP4o4kglFwl1JMpe2nSlFIFmZjMzYbsrcI0X+xp0uKz9mW1hLjd2CXuYEZ6sq
vgPHnXR2zoNrJcAa052LnIX/sp9yhDzFX+UcPHjRIb1tCQEHOR6u/u3LqTZyKzGR
+4yhKE9xthEzGjXm0cLqAY5O68/vNN7aQyEJgvZBjl0m2ktXsUQtGdBJzJrUVSdL
gs/B29isOCAXEomDcTbcsDPw1keSismmHWi7y7DGzenZ/yjogM7U7PNoNoY7T/+4
52JCTLxl7JRGZUuuyTW1qn8d6e/hKIymiIaKpIUO1xti5qpjih9VBkI4tMqSSuXI
LF/7D3SGshNWBEZ/FQ9fjejxOVStsV9ZtXvKMgYhdyiL9NGSWbfM5z1CRnTu0xdc
oQW+jA7fcw8sh1YqnjxJH39JlyPvHC7JY7F5yXR0ro166Lan/5czDIwOJ9fqc9qV
wyC0utiM+oiPWDC5URwzSpFMxgRGLS5JnFuK3ejnQVzL3eEDpQyU0kjfMrYxvzz0
cW7Z14nRbv2CBt/bIUJ/AIdTSpE6TgiQf9ZH/cZtlEncAYm4vR9CYToCgijnIiWA
xcTD+cL+Pwagbv0/7Q2lsihOR6AZ7SKNWZpY4TwygJqz2La31kYfs3Onpnbkhpt8
SEC8Xf2sIjoc2S+f2DGCpL++c/KoRd6xvv2k5QF1EBb3rBSaKISXWwHqv8S9c1ul
I8h2zS/v74AEgzDWj712oeAMI3bK8MmgO5DJexq2s5YZvCVD0/AT8AB5MxSDJzoG
7TlQVUKFiySOIPG/kHIen+yIcTwG2g9hOurHf065uIwmu2RnFpuIPzPVOmOcS29o
BtNijh2HUsEEQ7wK+bni/dvMe2odwcaimHlOy8OA3snUve+YR0BR1fQs6A0WF6dN
vfdswRdKTfwPnffqeMY4UvXJMlu1Bj470Q//onGzrQiuyOV5YAW38keVKgYkRIJv
7R9QPSeOntI+pypZf/XRp98l8FtH9VXAehx4xnL2BZFJxtO1gYFi01DAc+c3xnnS
cIJtX/8n6fj0X4L2hQLv+5tpzZxw1/pnVG33Y9T8cEXmVxtyhZn3BGMtMECQdQ78
whlQ29S/oPjTqmqffE79Md6jZvd3vV1o/apzkQkrlcH5/HbgpYeUHGhwT6vjY+zW
iU9SKhpDbeaIk+5QCWqppnc00Ww7qEpOGv9cMbtYueGH6OnyYTREgylHl0yuG49I
XnVtyxkCew7pLPs72HeQp/M82BNNt4e7q9VqDXvS2GTaQSCWD6Q35eMXhhlx6gGK
WY5d+/ke11t80FpC0zJ/rUxua5yBgRAMuzmpMlFBjtwzvpU2Qo+UpompWm8eTKh+
oZXyuRwOmMBL4R6kUM3x7JzGvUYN5r2pkZyf2Bgp/FmXRBV/472msz02Usu4+W1l
I9dmOw2cjsPef0xdFP++UAYzzJuty2Wsq02hKo4wErwXtHwmYfj1nAz6Bz3Mi5rP
5pGIClFFXvaqT4rIMDwpmxHpzN+Am1DbnaMHauzwKb1RK/IivTo3Dtnf4xBLbBDU
tY3TdEhexZs94MDks1WaJU2UspIEN/lniJJQQIqeSk9sU+1+Up1wVbBnz91GRHZs
FOSLYI2S3CaXVRPZRCDPkcGdqOJgzJ7cTuy7YCtBijh3uLlfd6YPHCIukff7GwtT
YUnXbgTKh6fipwyTrKXCxffQ2/rSQ6sAijOcBfjyGCEKs2Lzb42U7vabzefQlgJC
Nc97kP/OlxOhYTW9RHhE1gvI8vRva9dTq6QHIZsbEK6D8OaKGUIoz20UhFrUwjTa
xM5ehgZzjJILelbIPCaQFZsvA5tczjxwh950F1QB+xcjMjCRdSK/f2B4VRVoVNEb
aQ0DrCYLobiXCgg1cZyW6+xNhRsvOdzG5xRGrDLiBguBmNvSok9QwUe9/aStYlBu
sL7tENgxA8JPuFXtc9scuQgW0bGMMUdbb2f4lFQkK1X7sklTyG7RqmpjYLvCUfma
T3LnPbbc69NrbgFeBe6gRzb2LO7biODRk3+cCBlloTbp7eVIK3/1Dd29Lm11SY9d
705RbvxMeRfdb30Ry9sbh6Mv/QR+2rflUmzmCKSs/4JYOzehB0cGNlsHLyPrzq8j
wtHLrGWaW+AzIGux3+BQGcFuCnh2JrnXhQ4E/fWkvJ3sUnsr0/1IsI9d550OXy6T
vgGjhat2bk/wjrqxiQTfSDT7G+3M3JP6BX5gxfZvLFhfmCAymTN8q4WUdHx+SQze
xYwzjr7Ern4hjTnR796iIQhQnm5VO16cs0OPGAd8W+XFdpDRTUXvcS4T/vfc28/z
CO+z4PfQNVS4ScnJUhRoEpH4VyJxK1y3cai4/q0GBLJTGG8dyWedULQuBoEypVWf
z3uQWRN+w6ZoJnQwkIVqMN8QoN73UWxbh1I1u8COQX4Lk+igvzU+qX8u+Fio7AO/
ksbpeX2z1SuLF3vL4M3XM/woTnaWS8qExFNeDdHrcY80LgYgDdiESyqOKGGmw8hD
AIb+drodEt+jzJ/ZpHPMpNfwr2KgzqADhtfoaLaGggJkdYQ17nrYT1VxlF/5yOKP
x0Rz1AMmEo63N4bx6HfH8/MtRd96wr4FRmnvr7aCSjdsubI4SQsPDvIEfUa8ECUW
nhYDCfAmtSMonKgD/0L/weJ7Wcn7vKJubBcF4WuSRJxD+pkEo6pCm3QkeWVQtk9z
//i6iqetSXNcJIwROk6NSVmdijVqa1XIvt+410Eoa50jk8DgwvQUlGqWD/f7OWjO
roOf6pu+izrRF0yB1rtQ+PKy9jn9fXeftvoWx4XJ9g9Hf8b7ki0nD6wYDsxwcSVx
wjfFqaGsDRo/BDsN6oa7sJ7Bd+LukMlhwNcfiDxmRKYeFxzhwlTdTCpZjo9r3ZZj
S4x7jvm8qrT3xE+ofCiMsl6q5sj8rbk/EKj8sEi0Ih7m4k9c4gS5L+BuMwAGsAAO
PwZv0mZ+7RjpvLl5mk17gMhpAbmtuyANTdExFKcl7FmWMa7nyfWSgmx8AIQk4zCc
hQIY8oj4VrDwYqBTAfNCuZMpJHipe1f9FCly6Cg93XBAUd01QhiWii8x9tkfUksM
jrolBD/7fKhTZpbzJIntBZ1zlJNVgFGJ1W5b6H+qNMxaao8FxjCzMe+vZq9Ui6yN
cfq+EXfltUvl9utE6gMcQnC6Nurcd9Yk+/zW6RHOXwBEwpBtiE3iQt8vyl42hnXK
Z2eg/78XlPGZdj09gneyCPL0uEoZuQ2denrVi0q1YakhExrMTFL1sAIc9lCOU7c3
r3TG6xvTTCtfSosenyuPSluExNWh9NH5YNa95zRzvCgxQpAa/Pv5mSgb33ds7Huc
0EMjlP6zVLYqzLY3zLK0my/EnBQqrbz6ZWsugWk7PglrQ6o6TzGOo2MmTIpDfxrl
MEJLI7mlsdDEc1KJCIfcjGTFAov24I5kruCEuPhfZMbI15/YAxCeGX9cxe++8UlO
ApqUAqlf1/x7Sg/vEGuKGCaolXpeRjyCqzxNDaZ0YIWP81FIGNaU0N7cFwKmbDl1
YyY/ypXMvNKMGRziFVgDczPDb+8PVDhZSaNXKna/fXFnYz55BrfTKw7v2ESe9Ehk
NfkNJKtUdkIrPq0gvHONlcD29zlnEgUnLHSk7QFUTYTPvpr5qfr66L6l49TsShsa
A+2ofpgMSbhwsMuYOsrJcmkqQclFXatMJcC+bLU290wSwarPK6WX10FrQo4ca9Y/
31zLTPlwOavl/9CkNiANxYsYGQRDZMYwLZkheIg41T8wA4AG9JDXBbFgvR/N9bGC
TjLLFSma6i1RI7DUQRVqSR6wLrRX3IT3FPuISns5MY8CPF9iLsQ7fCLLLCwDVXod
KhRGkUBwnu81jtS2OoEc5cgcccN4ekYkDWGtqkOh6OulbJPSe9wfek4YIVIxoyLY
YXxLrOgBBRLfOISYcTzhzXhukScVTjFFCrjq3LC4c0Fm5/I+Q1BuIDqgPU8fR+Yt
IwZwIdi8SXaV3mCnpeekKzGF2ptw/SboNofz5WUd0jKJdPvgRmxFuIRuYgr7g2JS
I6bAbyAcc+Yyoicj3r9Fy6Ozqar3MhLZ7t+YWQ9RfLIXp2xqkoQmqHGpLXZQVTeH
ModFO3G5LnnKC307Kc7S1wnJNqA90d/X1+3UXo+cCkp1OsvIq7McofFJTOShlgKV
VlpaXR7oBaYvixDCVC6aUGzn01PAjrQ8p4NgcA5k4joo+0rkrPJQD29hQuQgwtd3
sfsL67QvDlxVvYNTRKapMVeIYqm8DZIRrz+480wumQiMfuWtB6cV3iv85vI/nmJB
OZOCFIq56cQAS0OhMSmpVZ/qscVtboJQ7Kv2Bx1OzoLjOm3yZJMS7VXicKoCF2jB
hh7ke/QtTh1F5ebp5usTkkLnh0kQLVXh7MwpdWwqAjxDIW+RyH2tiF2CtmIh280P
V/HW297TyYOpUzDdBiJkps/YlmO3gbU9CxCsFHPrZzRjxUEoZFtgMX9mTzShIM+1
dHu8QfhZc42j0cB2iHzac42clhFTf7E6L2yW+3erSchgDMMXC6x3Xv/+KEp5JMQI
xU6BwbDrG0y1XwZmi3I90e1eh2KfkmevC/9HB0Pt8pv/IdRBSo2VO64FI9+XpRaW
Yq5iQxZl4YcDsVSMvR5nu9YJ/FNieJdhK4FQKBLK0CNrlzkMyEneMso7LwAid+Qg
8ZlALJpdXpLuxbtR2PcvCV4Gnrm3D7NpHInGSK/QITPLegvNnIcfok32dxMI1qqy
EiyYKFZVxYonsUIC4IKkiH9ncFFl7XY1niWzQ+o9tNHTjulwncdZLvjmQ3p7tx7D
s7IV/Xb9Srt9QBsjc6wiOr65nJa/JGlsilvbql+ojsgbz+iox7lD5nJSHHjYUc6K
BISYEmmJVix8EZoJWdCx0RfCcfNgGJ1TieGq308Lddhvyeq5zsooSxmOuAaPBaL9
4SY94DfRuIgulegc+kNKjFFd16MZ5r+HEGPmcOpU5CjulmUm+90kqkJ7o1rhwoAh
YcD9xABt3kETvv1bdMvERip45IKJfm6MriJYNTq+MS+uXSilL+4TcH/k9ILM24dn
hVV9o6C04kQlKWWjtnttFZldCKQWezTalSoDbPcNt8WIyqTzpl4Wibsxj8xspHIu
W4iIRQ5iiNPVFVX8mvPb2G9TT2XO6L8l08gK2TiSNZSMcKrcJUMlf9MpRHJEDbly
oS8da+KdOZi5mj8PMY0WMlfh2cdo4WI/5OIsBYYVZon/G7AM+M3RHkpFT2Icd7AQ
Q4WWxD8aIjaiabRw3r2udlNAf1QhBFFUrM1bVPti9SZKeSS3anm5DNrA6kBE0CQ1
LKf5Z+DCCt8D+ZsjYD0XXbPT61p/STZytX3tDaDIVMYnPJjfInT29W0egTWdQU4K
b+ghg3ixN7Ru6pSRWP+nTk6wSYIZDHN2UoFjFB5IHPViaQMG856T2imPfgAkFPVe
+KLi69IL+IFRJzQhYyhAg0mIZ1XXIL77hO32XwoUlPZxW8uR1U/fOGuysvsNfRSC
2ISZAELCBL7euh40f0Napcc5RLOLGnx9XYDCPAJ+lNqUlRLL3GjoieUpSx3dLlI/
Fx1RvJFMBnzVBmdGPkkPcnIKTacUjICKzK0+CaY60Jk6IF9CkK3Oz5eR8Bi0vOUT
mqlPXxXY2ARlfEi2J/O4faThhjlyuXVooU8ufTfKwgSUcIu0ahM3KFkpMC5dWY7K
6a2foaUYphQwIznKuYYuHsSVU7apfyo4Ii2c6opFNGHGva8YctC3VujfcPRO/tmW
oDyxbPZe3vxVBUw/LZGSLaJpNZjhvpubZzoaSf5ZwWS8PuTmAfrGftPqrB5AKxBL
ZhgwcEccXVWKPe2GzDs9X/i8C3XdXOn9reTI9Rg/VCPvPmSDIvqZksQjWRp0Uc2L
3qa9L4BLno6du/VDGv+Udk/NWCoXT35nREbtdsCBpTaVQHbavFrdNi/QQ3k0lWO1
FTK8oHktGPng2+arZucCD/Un1VGDSCpSJ2zu5j29YYf9SJFSfDoU+TdwLemJHz2L
sdh1ZiF/J7URSeBf/YpQPUeW5Ba4v2Oz6EtTccNbDSYL7NOOHGDYfQYhruiwWw+0
SQGsoWq+EyO9CXRChVGVX/VM/82a1XYCLdmGVlOLx+xgfMi8lAqi+TxM7CCQGitB
X7B/4j0Y2x5W3jt3JjPWt3pN9HPNC35OnM/1gYZeolCLez7R2uBaNQN8K13A4r3l
Is00tQj0sc+bcBlnOdemKfX0cq0hJjz/s85i0nHZq1bmUnGKiDO18mHo4Il+4PLN
sxGMdhLz1Z16nJmJYdHuyBwS54tFP3qqbCwFwy1AG4CeGF7vG/rCNaYIoineywUr
Byz+TfSTLzZ8tYGV9Ur117BJ/widwwAUp5G0GabBX4tqUtZXL+DGURU7kz4Q2J2/
qD4UE/p0dyyGsFoozFAcijrBzFA6C62EKHLnxIhSYEKVwsxMXqWoFvUC+bCGKeOY
uhkZweTVDnkdlDo3dbUY8BkZ0/1nMYZ84TddcSOBe2OqmjmHhCRoIAWgx7VXw7fh
pvQYDKZmzmC8FElVgg94u7YvPgqEFoh0QBSW61fVeS0Jv8USTRIrJspBJrQ0mNGi
qpagj/enZTQ0W9P28DBL+c+tyGUyNyS/2smEicDkNx8jnQY6kXZ/Pd/QWzxmmvKf
LWFWydNRDqFGnqmtqaic1/EuymlJdjrX0bN3uKf0Tc5ttLjygoKOg7ApcaZFz6/t
gp9DicxsIeBk7NUAZiqB0TGTlkCgOdrYnZ7Ojw/67TBWVj13k2piBqMp91c0oHeg
vWNEGJ6ryD8I/Sv9DjE0J7fd5pX/QJk+wbmtCAWOkUwb4RaHQLC8R8JKK/7m/p+w
co2Fl1fy9Egu5fe46Ceb9Eme5bsjggVe9B4IS7ZcpG1ohMoXSMo37wwOFQYb4TmB
rDJNyan/9aYliekZpLY0PGa+iEStYKahFe9qEVqX98LMHjgygjjVbi7kHh3XHkDF
meQ1L1SAuaKxpJgG/RVIH3rFUa2LM9NaVRTVtRBqBPRwb/uqtrGbvqDCwdi40fCt
bjZcKrhlghGROy7cNgcGHWJbPm1vgeJ554IAeOlDzIRS3xlYeoz9lPvHWWLbGbe3
V1Lu4eR1STpOADPDj8crCh6cRaM9fLAdQcgs/HmM3jdGI8xRHzRsm/GXFYX+7GR+
oPYH9rY+bRaAbrOvzwsVVgQe/uM0LUHv5TB+lSBPLnnGVHxl9jFmAR2ksprMvEjd
dBVw+x6VOofjELRVmMcIB/dhKVwyTMSzecDWsiC/MgkEuRlFaj4AXO8DfRXKL7/V
gZIRlMFZMBzPC7WWMri9fDO6JqR3bdmg9yn60lQcaBvY6VWLqZnJ+5qrwQjSeigE
wECovlQqd93cBA50M1GwhxLeP4C+x36hB5NnoDJFLcSmTFiOSKqb2ChOOBzgalRx
0coXVX1uUKNnc682ZIxRvlcNixw7Jjcm+zkSVrovUKLJYdpo2qq9W3oWwvqHuotJ
0FGZuUQuBQ3Rk2jCnmxP2f06qDV2tJmE8vTmaJXYRdccWtGTe0zj6e+SzWQNx9fP
8KFfCCsCgjZDwrU56HwmKirL5nBgKH0rXWgGWV9YXst102pZOHClauxYmXa75cHW
HJnhOlhH7yvKv9zoOx57CKvb/4KIYNWd3/kKwYDaO0fBkDda1d0haH70NA+eU6Re
e1aDTNBCYYPIEqb2ZEMB2S0jA6s/eQih3u62u8zoOmKtVb8UdhJ+7mWwpSWPxvyk
ovZLVzGd7JmPHmUqFpje8AE+j080lz1PA6CITTWqNnPPAeHvMEXniKE56wIHMsF2
FHmCuhPfZQinO32bJuge/lJBrFzYW3AvNJccPbK3fo96kSNjsrQ1PKt+Mm3/JayR
U7gBNDP0AfQYsqSIPdWekeDsj+X6xzbgIi1eQRf01zsSRhN0azbDSVyoZRFagOF4
bsEPbLrVe1etrE3B4Zi1+p9qi0LoiUEu3jTBr6xZatjP160zx0qItY0apKiSG4uT
z1s3bsfD7NG0zBU6sH5tl0aV1WkqDSTHocYrlTQFrJMhzfk+Kfc2sYD/5J8I9Gkf
y54z4Tv8aSfgOxQWTPp4GrvI3erOjZuYro1pe7iPdY8RZ5KmkNK9yg8+Bpbwx3wz
AHs7m0uI5OUCsh0ajhOBeKDxHBFo1KqFCsm7IQqptK3j01TkENGaeozyAmNHsacF
JvvIsIFS8JNLSI7+exAWZwjp6yy8RcVS9qrcmDxkws4SgDfEi8WGf01XfIPLfm9S
BKwq3gwysX4cwMieNkSiLbl6x0Yaj3QMFRBbhBCBWRUM/KoTyknAezVUjObTk2D4
H+WuEGDoL+kiGxmApuWyGkVhUY146QzEsKx1pd29aHRmoVWO9Ly5YtX+HquU5oqu
gsC3QsqjJPca5mYXpL3AICHO4qrOFfvlzpzZ/qbuNRpaBR5U8fubN9QwtMESHR4u
W/X1VsCvzsiQDrHnAT6yu/a8f+M86gMu/N917f6xRyLhbRdXxsk0eaP494d8VCG1
ukAniV4LH0yUFma8zAOLOymFMg8Odu1SoKKhN/0bXBIvxwINfes7ySSRpfzzt/sI
cSxJIweMDD9L9L4XAwIfLB8lnwNSGRupzcp+WoBQdCy2FGFp5lU+dnHGxhhIfyrp
nheBWiep+5ALI2eFomHxrKIJWiNVG6m8xbtfwU6lGXQ/bIFnCm/uDOFp36jF8kSS
7iSrA7lXWaj03avaqJBApLRMelAjwrcAEQFSEMFpQDnCSH6hn7HiSOvRBZ0gB71V
cxw0b/yOxuoUpzmYOnMS8/no71b6YJCOav9T6BZqyGOhgm8phAeuEvNfT3+K5uYz
Lxs0NWv09qRoWbGrKs1TZqyhmfAbseNtdCbMERZbjj+q48+EkFDwxhMd7948+FZ8
bv7PVEnKdPNTjdt1pmTvx6mz7aPKIoCNcB3E7osjDgRpv6GLTkDihKnb/ksL9vio
HAoV6UjBxu3NxP+f6CGndPh4eMDwxCujG9E7iXgCe/Pt58NthEbja5hDZeLy3NFb
5K8bTtPr8hKdzZdZiD8jkBEo3n4OkkfeRAqHYttdLr/A5MPVmxQ5GeJzuuRBWhyS
UezBAisg90O5CoeOwDOtJ7LtGAcGyL3MkRCCxbWrQ/p+QSfRr60dWJBmXgxmXre3
8avmmcZbzKi9hf7uUsY/RERDFxwJD/RjSLTQc7Fs5W8DNOclEPsoq1xoOrGwsdeX
MBerZn0oGENz1i5A4btgD8fD+oIJpnrzGb80NRjZ0I19z2YtBoFZnXdbmsoGi/p1
BrcIuOEKnhVn4D4GGrTtdT2I6gCicA19dG9D77sGIvRjk8i/XNQmRzCtY5M0Q4ib
x/KPUg1Fq0sui8qLWQMQN17em4DMoTLT34QnucZe7fwWE9Ew2G5+/NboDhLrIomi
JLe0nY/ClY6jTyupjL8kzXfs0cgP65vAH/qlwcW5RkOC3Q53hq8edT94CUQcUoVR
pR8MoZZ1k59MWURK6U1AIYoJz/3+XPhJwCVrK18dSZv/+13fU71yKb14YZHwxtX/
Eey/JDUt6Tya3iBgIBrep/Oal+BsC8KwFpQYWrJ8HXLb0FDG6I9xnYrd+0fRjmbD
rR+lfzqxpA5A00YBUiRz60DI07v24sg1uHomO8+dsO5iqgHqXQ9Peezf22JM5DKk
X+TdagdL6rpaAfQ9QblJnJn7M6iB9cdR1SwoqeyOqted1yjiwHKhC6c9T5rE83C5
hf8qwfFwgx+Jr9J1GKp52dq2L9lUKTLCQD9EKm6gitFdW/G5dKH4nqazI569hKhR
8bQc0cQi36bXb/DO8rM8IPLvZ5zgzZR/prCEGaWnWgEB8STUADKylezH24YZuiQH
n5/1y8stuYjf/KmqVn7+Yi9MlgotZiM9XHaRRLT/ycsyjQJ1RmC9apWTSq/8wPzv
C+iCYJNButo8o0NGRZPq1Y3THEfFkTWyrOoGxUB4bC9jdfQnrhL3SnivPJKmOTMf
gsDyetQnuTw7oz/e+YO0wAkEgogAYdk8v/zQ+FuX+Gw9fHBAeu+K1ttWhRFe/LfY
O8s0U0KO57WiPCtFZ9j6h4/KROC/DV2aCaMWrWIgu2K4OIwZh7+zfAFO3gRkV/Je
Ddo+sNhAPy4hjpUE/azQTOa5f2xdR+/VjW2pPjZQQEYQXe+MM8vNpAEmav246Lse
CWbkoDvOIgG/Ews9hiTLSge/fOTsSlSND+DjN+J5mwL+mhJoVtH+03FT/EdW6A5l
eC919ugu+mCaGLBUcBNsg8KwKcbKnd8ZYSfTXKcsLTjY+XmllsOlN/fgFtrzRIEY
Tfhuwq9N/GTJVjgQNTnEtKA97KH2wQU5GNtuqcZLcMrD4jD9OUqpdKe8XLzSrTaD
TAL37y/RdHrT6UEnzhhxmrbvWMk8KtBFlEBovjnTcEHgsTC42gYVizQJZ/rHvcGs
E1UKc+aGU5BuKf46p2QX5Jm76OelFJH92XaqRRUbmZ3a33yM2BAg1yOHk+e8vANV
lKaKARxhSKJSr8boDPJd2JqAxfkyIas01tTZx7RbOb0d0Zf0UIxrj6lVFsWFgqtZ
nxe+ALwTgRvPSMUCFGWwEQrjDWmA0Y/19fDXUcXy1uer+gUEDiHqLKCzNFEQV270
FnqIwlJGT8YL2nWk3Pk4NY3EIme2rQ80GCdOSlSRB+jZA5u80nPyB3QGz6m5WEEL
Hi4u4aWNtJRga2nnylT914Qmq4fCuVL7qMOw4yioPlIt+51Nrz6PenDkh+qb/w8X
CmVv86FByZVqS217afIqzkVibDv3K9eF4HB+4cSFbIgiG4nVEIeZEKH049rY1Lfp
ohvC9stXam1Dzh4fzooia5C5bt4WnsoqdJzxMWaOLnv5MSeXMFvNtgKACDDg+Rln
jliTHGT5Mg6WTgKoK65vzdng23YQGFS5hBIiBuocFfHlpkR2nY2LFgacqT0aq9O/
4c6foYuN0fmTJpQRHocdKF9DooWNefvicCwtIYj804DNbc3Bs7mSLhE11CL2AFbK
4kDRwKMHt7ZzZciXXRk29XECXcs7IKQRA8zaZOPLeVLQ5iBKK1UimpSSE4eW3PtC
DomiL9i69EnuJ6s3WvXXlQteDWwRqjybmlZjxBCuCZNatmSkBy/U/F4iMAVEaU7H
uTZWb0KzMBrrR1s91xVzAR1AynhCx5ft5KSWcoQe/mC3Okk16SpfVCyLSUD6YH1o
9t4iXRtQfViAYrkKRzPr6l7bMgZYpeOjjbppUHbR4dlXuLC+As/mHGE0CgCrdNN1
7Is4jqOYeZNs2g2XwoZ9FYu1LpUzlYhgu/I59OIoqXRIgyavXeDfhhpDPgLIlzww
6nZVEth/k8rgOGcjbCJ6zTICmeYj0DjHWdn72Qhnhffdn1Ge2XmCzvP++k6NSLdq
4HGC2qLMAyv8OnM+Jc9WlCCZRcimknxISZaBMDErRMOfVNSBW91WKkoISiwtDDAD
bB4CSl5oIrSvG95a+R1gFfgXCfdq5vSUaVc/qqKRyqYa4emcOhi7n2rWJ9T8epNt
ZFCRP5qYWprM/8s9vzmY9vHnoX8ztchWD1RZqkjMk/IS46XAb85saeB5HEE6oHtT
l6D4ziIuHflMqJCAeDDlj1Z/iQ4+cyHxXHQ9QaHDPOXkvzrp+OdmxP/bC39VfFPx
d9+du3dcQjf8zl/SbZCsqh7MFEFbwMH3tzz7A1q5yzyiIdf63PiAHmJ837ea+MXT
8Q+LMIs+SeI+ldbJzgQAZNZCBwzMrCLfFa1r10YfrIdwqY1U7IH87nNSuV6a8FEA
cLOa586Q+83hRsPH0th7Zsi/guf+oJLfYViZ/qSKz4sUav88cVDyIKkijuQnfK7K
NqKrjuvQT6MiOQhuLrZB/BAyxmZ5VZT79eov0nJaKMUJFOrx7ppjJmAkpE7SoeqW
dlUnqhIp5YuGUmgKdxzOpevOrO6xCKKlpZLxnaVLKZwPe8lnWIMHy4BrD9LiMj3E
/80Wr5v6AtaLMkHHesoQTgksdsjcDssIo7mzKcM73C7RPc8TQN9p7ANFKbwoIHP+
96rK6VuPuLfZmS/HqRkCRqdfhB2RyXBL00ZjKYL2dpUxkWx1Ug+bIm5ZwAdCaQwK
n6OS3nqq9VD3C6A8HNIGMPfp4veOwxvpepOsbVCtALEmkiuQ4H5jJvRgBTgEOZsB
RzmiAMAR7ivYd+c5vIv9DZW9BIc90BO+zEaywOEsYyLnBXsgxWtn86TJToZss46g
e0XB8IrxWbXXgy8uaFlNuyv2P9dvikscJYD+tMjLfHYEuE65txgqT8QZdPBOWxxT
CqYZLsa9+FxoEiP7tqijxCZmuIvwY3HSNJ8rZ+9cuZiTWsiYh4QxRcyXrfKLIZ9E
brwgjs+3IjQSf4pLyLozkC6EZ4FWJQImYNsYoEWwFhCAOcd9eZzoYAj4MZjDx1ea
QzO7NR0YUHgGfAcjjqEhMpYp+NLU0P5Il5m9jOuCZ+gQLzI0fzvX7dFUif1gx9ES
ZZJ35SdsIrUfHyZvXMSGrv47EPhs0oUk+fSD4sRipLBk9zVRq02riJfqwOFCHUoq
sSQrCbKeXJwkmxEun7SUgPOFumSpcmky7zsn1iMDxr8QFFck4SLQcDPbw++A6UJj
O961buVq0vQDOyulvHMw1+1ZWhiOCqNgulT/mMNP5lsyalA/6L6+ehOzOcU9odwG
WSugIhIn6+wsSeDRSGTMWZMnGdx2YjojfuV+rBSTPhC7OUEJqNZNTYMwMxkuw4AF
WlTem1Trd6SnDwd4ChEsxpMW4UNR9p0y705MrtOX6Zx5UHa7Uz40WrLg19RLFca6
Zmap9F4+d5UQowCEiYVKjJ5DwquiTfhglAQUSF0hf81DtLOY52OWf/0EXrxVip4x
6Iaz46eRq1zWiuv8AIatTJpslVAnmYFmxue2eqLQq8sqZO4ARpiNcz3GMbCUWjp1
7VchON9GcngtSWjYkU/ySRRu9NlaLQJRgf4REillZ5bt+/+VsZgUGXoE8fXODrrq
SePq9S7b61wCWNhxi41jlRVe5Wyzsi/NFQ+e8lliTrL4kNE/rkFl7EXQOKGV1pmS
r+RPTcJDF//wIU85JbHBaJ3ldQ8m0xC3gtbVfied0yfUDLIhpYYkQXhsv1+MFxCj
PrKwr2R8FO0W9t8hd9RPNGH7wUdq3XSuCij8XqBnSWL4y5GIjr6V8TV6JBGTlbzE
o4/xnisYAYYM/8SY+vhacYrHTNwXdphs+9NOoc/B8tXCUBHCdxLvWlovr2+0zoFc
VwyPZhKivlyBi/l4xPFNwpLEeaBEsnwFjs3gBmLJLRBfqul6Ws3oS4d4oZA2eElZ
mgPlVzcEwx+2GrW41QFQrTDZqZzPKtO0nO3Begxanf1y261uMtabnOSBtJEHKTbw
PGGxHvg7ZdUU6Jy772Ft54+5r0rJqH4u/dlSGGdYUGlEDnmQaC18z4oWK4z6SFaf
4eCU7BG3snX8XwSSPYVNUz2X2xscILiV7URRM1gEs2FlzJn0pwj0KMw0aQbmqe2S
l6MoxFipD1kZHwzN9Dm64+vTyAXqVgK1ltUzYMzBOODtlf2nIvwtvHYuXRJmZOLs
cj/KL6p00irlV3u9FjdG8guM27sH3b9ZpiZObAtAr/X1MKBYil1GXmGhTRAkoqY2
Ba2iQ+vDzxWZWrGgrese/0319foUwm6lwHBGBPOOh3tgePqjEep+2B2c/XaukMp/
cWwcE+Hi3Db1dsqFu6xiNbY8Kxf5I6tQCDqIKZuukQ1Ea1OP0NjGob5kyvKdAtv4
DWKJNfgn37iTvqh2Gh8bqmaSzygJN1hAv5gfxVnakkNpjBxta7NhD05zajLLbioP
gUoHRM0jHOBfv2nl+KfmlotOfGWsTITC4lhDXBsxG+SqAxfWBCbHCEpD9FVnvIeb
khpJicIJf7yLsQIBe8zn5F59ykDLNJwBtXFC1eSrrllfw2rmsatbIwD0MnNMJo8Z
oC+6B14wPx3URRpMMmvL6RVeFtpOosLxzeSyZXOPnIVgtYJYBhNYz7iW2XR5KqcT
HjB5wcigeXXF2DePEnRvZAWnbkq0PCx6GMo4lHFJ1RxDM/gcPALdeDx+YX49A8Jy
tVobEouRtLz/fVGu87TAFPOaX8fMmjiUItCnBy7c4OCv3LhACP2HUm1ttNTAcl58
oIfnQsTlcJlTkGmAKU3mYpaSZeiyXY5cYm8WZ+uNB2v49XRN2OEMNqWebt6guYvU
enrQtmF722SICz1ts/01UifyYvqQjlc7pJzs5+Un6VgpII6NRc1RYAt5R0ljx66P
JQBl0qd6Kno6wG2H+9yLv+4JW3YYDLCgsDSPMU/IOlNdrpaW94+jhotxUjHEEcqY
tlxFnqOiNYaSpOPZlj23ZOE/1UwWzsgZfWpMEO/0Ewp89qffDPIuSYKdWM29NStg
qXym0e9nQxKVXbg/ViIXSoW4Fdf/Mtf8FyHdOmeQm4Ao2X5N6GvsHsXRJBKhEU3/
5HbDTsGAgn9MM88/izch/qKPq2a86WZWAvny45wmW+EB1aC18pmvMJtUg7JHpnxz
821EhHMJElAUZcmQEDDJS7VlXhxkApfHn0FR/A/Bfqldt5hLVkCaN6q/NNHPXz9f
nwcW4snNUx40sizsmJxXYmsbAL5c/RNVErdFYG/qMCOPqXlszdJzCeru3+nXEema
CEQiNFGB785MvLWmY072kCvm9Wi97B3VPHvuk41r0ijRU5ZLPUP2EtgaC7KmqzgI
+ExLnSQ0KPeu6Qqc9gPlLWT91mtNISILNPZ47udibiKbRGAED9fSCFsD6vut3hNU
mXDe75qY8cP++WEdgE89PLdZREK11hdQZxag9qSv2ssiJws32lygWgSqHAx8mXhS
aCHeb8eiqXmR7DvxGZEFfz19jxegBAAJ7IOiaPrGeJgMUkH6OsXetxHLEdZuUG7P
Ckg2ij7ZPRUGn4A8pODYo8wgYbCsnaDh8mBDFIJQQ9F8JIaJVKV0+/cwWa1OdYJw
TSDOmRYiPf1lsDYguNe9ZpGsfjJiL+LY5oA5ATVFiNLHUzSz/hLTQWZY06/CS6/R
E5HLBhAUeDOijqdIvdkQl9F5g3k3bjTjkSIrwu0695v5xY9kjMTxB4U2dTxd6MCC
thl2MnOaLtrzR18pBClctHxPJ4KMx98M4NbqaKC3Fju2392jvc9dlcHHPdYIVDpd
4DyspRAXQ4vzcskYF5aY1jquUDLWDE/+UYdIYb6b+4mkY6/mR163EC0jVF6q67s6
cu5uNYdlcmLKCY1nfbdDfEwpW7V0Rl9y1fc6nJIxqjo+8CQlLUpfYikDUS7LDQS1
3HL8dHG4YwuWP+Op7HNn2h+seln04VAJXrZAlVZEe2P13YL8SF7WSEbcX403E77l
VYAbOqWlpo6tID242myAKKRNw/xDZDfTN2habufOrxVbWxrfEXLZwtK4rqhHJH62
7FULA8+5hV0VbM2EiOhmVDBkJj9eYuUM6uUXToBocvtUNKxjhQ6tP0PufAiD+MmB
hXDcWocPym619R29/Qt7qOleWV72In0j2Uj22vQadvpqDqtV2O3XPGfZhvdGVAyr
hzbq5X5BsGhjiumBOOdmEOJLWQmqWr7hTbgUJNhIyzzyovPE1++LtxCeht3U8Fi4
plvw8lgJtv/OC21HA+Vu1FQN7OFaIkoStHLBLQOUEso6ITNpOLQIDsAGtcVE0dlT
jKZn+SbNQpOqDI5S31iF0MObonNPe4podT2GXOWZi/gzrqeTngXskoI5oxDPLNOS
zqMcwCBc9KQ6RQZezbu7m3qNmg88fWWUPaa7fMdObWue98DE/vvq2JMvHoFrEZIG
KrQleg3/OmeXdo1Y21OxLQP5ATLa1Rmt4wzaUVGsbvQZ2fJwG08DjqjU1j8xX8CA
9/8GIz9T2AVZTHplhQ/QNjl/f2PVH5RoS6AOFt3yHK4ByxLthvaCJUW+ImsV0Tys
ibruW2GmhBen/R78alcyD1e+3yF6Nv6gSZw9l3Eq1N+TshpIIVdAlim0pgsk4l05
7E6+0e/QDkKY5aumoX5QursYTbI/wKh6uoXaVnXZoBiqi7Rv1mwhsXn0phtimLUg
+bXw9QwxD76pGpvAvzPCG/tkq23Lk27P7nSeCH2aiXvwaGsPr8bgbcEyRn3XZrN2
uxp/XHPBZalinM4VMFGZYRTn+lsTbUckQ2H5Y+geFnjch4d63QtLnR0Fg9VtZgIP
CyCxA/gWwKDK2Wfo835a1xxopDds2cbGx5NtHzshxmhHOpd5hyGpAypRzgNOp+dT
/BpN9PHzV961SDiiz/YF34sFQzZW3rB7UkU9Vuq7e6WeblFx0HymRN0ZPfodvHBZ
agqelMa2+qEQaTVRVzefSAc3suCXuUqr7BjjDYXwcDkpUQ/MRExScnPTpfQfB2v+
u1uVogJ9wHZ7SrPgOauWTJuG/AcCNjHQ2uA0nDmKZibSXMxuYBd8eUEnJLSeSo/D
NsuYMbjT1k+YZPQX6PvCEB5DeZYDozL+zZQcRTS4R1kttv9tKfDELIWOUiK5dmB3
nfWC/c3eLBY0nfY8NfOexhC/42sU13KhBo5WVsHppnRu9K6XHtQGL1KHqApq8/yF
wTOwhVOTB6KkSblgYtPZOHrcnRLB8be8TL9w1rhMg2imWd9YfuzjpMQoRfV2YAmk
zmAxUSAJiV6KTTUgtd2jObWEa06qtm/VfFeLfkTStTg72mZk8WyhQYy91b0fJ9p/
AyXQKgp3c+OTIqdg+VCDCqho0rvGYqfuEGGMglcj5SWe3f3aIHK/0+f4/s4H09vw
r9DE8Rtzrwy8wU1Qvjq/LxbUE/8VdOfPaxIKokw/QUKqUrf8kMzPEupzjs+wINFU
PmnWGi5QI81sxsERrPnvtxiTi9VPak2hrnoUol8IWqOOuIarEz+dXLT8cWA9Fea9
aCxQ4stwEqddvKkfRahUSlF2nXIlv0O9RDqZFzN5bGOsgvTvH4Xeynm9dHjZF4n1
2IeWKyKeUquRt4kqJIY/u2D5hiqI8ersk5EQF0+MfrKiVThngXgJFjZj0ZM/ou+e
marLWFY0RlAUei3p4gM3Vslcu1CFHHD5XEJP2+6/YJivFiVCgBxs5qigEWH0JpEX
rISlj+XhvrSNGPQgkBEEI3xqfYnxbL6V4weHiwUD0j8W+ubCt6eIndORxglpYyAt
BU2KJx0rZEv4NWsdS9oyBBd4ypN/UGX9XMclvPrD2zGBRagVpu8DxsUQCMfL9YmS
JNFH9sC6pq2GOCb+blftQ7oYADOI3azra+Bps4x9O6iN84At8cNzK16nD3kEymom
wiOVP3uBgYpZ8DguM6xhtGPfLvbuBA5gasTHnRkwqc2qvDyiySyeAT1d5WkNxhOa
EUq8iBwxfJ5WoZE7Orh1h3l3B+pl7zSTluqMjqJFifM8APILfyXMppGjgiRFxZBl
jILElz0ubueATA4QvFNvI9H53hE7Ll5pkotXscqiLkHTFVyI028nhm0JRF/dK6Oa
NB8JBg0eobTS1xilEJqcEreW71tFH12yDm1RLiqeMHNZZf8a14jVNK6esMCHbakx
dmDZMr5+v1ehnwlzIlte2UCj15+n0vrljVDenjqagu5PnHY6bfnWoHZMXFv0tEhh
5VZmkQk+zVi/iiMQv4h45nv8H9Td4Eegeg+TIrqBY1nNJi2Iyhw3o5ptW7Z3IAas
gzviaFQA0naVpdhb5nrowbKuNPj6brW+YUI9ApjZnxcdO24+MU6coPb8k1IHAqXB
2hELSMFm7iCUq9x4BtoTPW+DbY9MOQlCpTK8Fs3cEGTScUZ9xkcrCZEexkDrlYUx
gyvNdWvWzTIGdtFdpoTmT9yZh0Il8DgOAblAVXCJWf2io8VYycMZIYctwZbOzstl
s1kg3PciHoLXvDp6YfekA1a09ZhvXCmXxuKLPWinBl3B/xli9wkIbA6+/9JrD+lz
MP78ckFuIbTZbEMc/sTWSxvLgGA8Ucc4nfN5zdqTRSO6r0Xq9MNucRfParLekfZ3
vflz7E+BszBI/aTc0Gd5ApLnDwPiigVO8qTGSUJTH3gU5j0TrAEzvFDxJN1vi2E0
Ps/eFKDaJulBmeHf+sVypx5oibN4D/H6xDRsrQ+qixoQyFwkkW08c9UB7l8vldux
WwTNgPnsYzKzKndGNz550HpxJoCKTXCsl4sdI4FCHrEezYv8ld3BZ+/gYSkBrQW1
1umbbh3goDKALbg1rjceiykFqDOmI+2Ny0dHCybtkQZozBPmC/zhBK+j5Fbuw8DW
7Nx3l1lA2KquJW5yLXoIgAHbEwnB2tYVS8KCVeBD3VGl3CsWekREE+LOMq5kZbEt
HJwGmtnezmpm2h/MIwP8D9VeKRXGLfXy0twIux15WpDG3N5zmIabpa1RxZVqXLtB
Sukgy2EYDgjIhNWHBtz2SOJjMMdPNDPfGyhoQT1RfLvtpCIpKi1uvcxNnWPWEYkF
vkGVlEOBCwt2rVI98mKNG0qA1bX7P1Rg3+1FGRkDURK6pIxmMd8/2HVRa8aongDM
Rp21k4UhyrfebaAfBgCM74/GO16qnrTcMb3I0ku50GrR07RRQ/W13/Ucz5dhVFlX
zrFaoiEuk/yQWdn5o3PCzPsj0nDXSW8qJQTUDDckjm03wAVXgQLR4qzF33Jr33Hc
Xt95QGmCD/Uly92ZVf5XU11vdMJ3lYrb7UTt49wf/8l21Y2gsa2FY27a7yE94Alx
V2/C2SNtoPSE2Y1ROYkQ2/mPnjO/kPYazj9LlK2BYIAJOyp1ckKrtYo2W1DaT5c1
J/hb8FY6WesP4QMctf6QVAfYq5qIlK2dadZy6JxEUfVPjAzKmn+W0GzSjCXqf/p9
v2C/7Q/xhUovEZtEi4wrJvLxt00LiwnzAgf/erCV7IUdN/f0o5CjUjKcKLnkCqNB
4I6h89XvX8XPZo3xlOm4sTRb0XJnu2qG9np5ZCj2b503WqI/eJtR/XhUyI5k6qnF
5tTSiIceE6RigOD3JQOVBmpzWOZZSQNcJzxb98Q4XOizaC8qsFUenxTpuqij3IFk
JlnuJYsmCSb39ZqA4Flv1I+lhGhEw0rL04HvFsWHeQrIxdhsSblqVVlpcC4fDk2b
xUv0B+nQFeDNLYbK7tosWRk5vu+zO1QzH1Bh4iCl7bMlGqMyLqXamS1EDmpFEk6n
MMlHFPP6w1Qcb9ca0ghu3KpHJah6vusTPyRBhVVS0G1NxcQZM4nalxdV/74bEd1L
EvFsuZJP454nXT7V8b1W5WrELMyM6RsslCYQHjj2fUH7EezuJxf3IV0HbKUGYRn+
SOZXFZ9aOugOvHmflNfsx40sSwQ5GI0uOhQYRvl8sXjZfuIIS3TazLFWPg9AVzWZ
jBhIsYtQ6poTALGGHcEwBP3AZJ8SVJvLapOSqNEEKiIUhVCsyi+wqa+3g1PG865w
O2nWy8dFHMxqZJUCLDTJeAEfPJJuZkhCUpkxqrUZ/gHwEGYNRYGl3PhaEc7pz8J1
IIBouULYAAzswpbl1SvvjQu5twrflHzECSHGaYjECQzpFHE4+gpPjo+ecCTWSeZg
vZW4xItpqHvn1OHExCKz5H7J0TvrRIHq8k/R4EjlbIJ0XLeZnw9byvEP2vz9IX69
kfjchTk6rWwxe//2E5bZWdadlU6EtWIfUKOl3UsTpbglRAbVfUWuDXFe83Unngxf
dNjSSrPmb5z+atVmAnA/oBTpbhW810D800vR9dABZVXf16kQWkXtr+4DpuW4r9ih
U91D68qK+WB3OjcjUbSRwGyvmrwVPOHksABQZuw0S+JTkwd8tsZHyntwA2sCm0ms
wyBGg3xb9jkDkBEKebPE7AIjwluHmbzeH6XJ02XY6dZmvWWBHAPFCfgwkxq6vLqZ
leRU8npL+DhvwBPh889V29OlfRmT1HA7rW8QGLwdPY6ehyHkueIZ56iyzSYNhLvF
EWwqzEQKQj6HD0a1D2KYjanOmwakrjelk9y/Ju5BqmBzJeZIc8NS+70i5Cm+kyYk
+PxLjnbt4kb/d2zr1cydRes424wQvU+plmesVFUPdxNy+imQdpEL8cAlEhYiMfyu
Wo2hgRjkqNJlG8/h6KqxzBzAlwTxFSppWcuiPSig5eKOMKTnomFdfPeVlhsPhfOm
kXed6XH1OgvQ1iR+SoMI05u7qQyBGMXevouGk8cUEIsCUNmcZCJSLDTIQYBfVZyM
Nb6HFqJ0ihCIbRPj6Cm9pg51yrB/K4575EF5NR296GlOJ7SZZ7Vg/BTw9zwzw4tq
OSwwF83K+LuBp1jWFyCvJj2Ag3plmbUvWGG4os+AAiQXmRAoKln/GC0oWAPcx4Xv
+zqUoJYF4AzK3kbMtsWPYcbbMUMy2m8tLJO8QkgvnuNOkqBLDHuNqYtLlXN+QPzf
59E0GLZoB78oTQU+DBImyN5LdsscbpHnorh7BUwMQIiCF8mLoz1nQnaDIFRCSgPN
WPMInafc1Tz7A3GEOx7BPHPCw59ekHDgc2aoncP3veLNAzHobOwGOkhUsgjJKFfx
9keY9BKXqkSRJmZl9+uQhXMvznRG6CihqMK06LnaLS3NF2kbgZEKgWdgVicqh9oK
Nyc9miD8FIRpOCAJcyRlHWHHrelbe1hVIjEpsfTCCqDLplmhEcuIXCWW+zJUqzZe
q4Hi2A8jYjeckSu9vvaLdSRn/Q9b3WKOiaTF+pkBVKB8a0/SdtXxmFb5hCDFDajD
jGi3ZGM7OK4D9g/ywhiQ8kQOJglqTA1NBbPseXGNJ91Yhlla+M/dHV4IKrpuqYsW
RZ/bvHMqirex+0U0Sa1mfkcgr1U7/sbbaZvj7e8eQOFayPMmLo5wokAymAyxUz9h
Q9pZ3FgEV05OiNasm+qN58CotwabC+rcS0tWAIbmQi/OTeFAOk8e6RTEWms9YGY+
302rIVfRo174Kwh04vY1+dEyjasQFVpFZ3c/6+l4FNvpVM9Y9/CAHTvxUp4kr2jE
RidcQm6dmmIUBQ1S7DxVj05xh+dMnPQLe7v7Ua2QAO8ofwtVEcIsjtl50PCb9FEO
fl+/SHLfHTFQysUNc53QjWSnpFTiudZXFsFIAbtNCWiGIW1e0GTBINz5nfypj4YX
A0HMgd3wbnQsnVo3UFgvPXyJkhlOpDklS6TWGzyvY9F4B09nVkmGKNGGkMsq1nxd
F9Z3IOzPlfbdmF5XyktSQoeo2/49Lr4Lsf6ZR16RHLYUTdXP4CXgvCiwbZuC5wg3
gVKv+oG2W4PKuP+XIIr9YFYdxig8qT087kQ6WL8HCxkrxAUrMKa0bNbtEREBhwI/
JpzoiRpDqaBCkqtaiDrXbItGbv11m/zsTTRrAsxmcDzC+S+NDwm2yYxzv09fSigg
sL781KJUuoi4+I73Wf3GJgnzDBVL6keKq0Xid7cCkhjPRWfez+/fz6uScH27F9ER
Ohgj4Eun/vX7iZrGUSLUdfkPfLp6iD3n9kp7hDEUUg0OjpYH4KE7N31uJszGImTU
0VN5jYHWmEorlAxwHVB0qlNQTpfhgZESv21HL87ZzROYTCixTCq6Cg/Fn2tDzdiv
HrGY4EzrFSNA2bBatHzfkFgQmXgwj+4yw4sZazW7y3QgEDfRxJUi7q71k5qeKQTw
DzfVbbBIJpf0ReM4PtZMuArVxUnAB28Mt0G5umSJVgOZfiv6shkXasI8BsV9YcYE
5NHicTvzlAkYu39lCqq4G4AN0WrVfRj5WGlzjgXkSd2NRM9/dn9xEWwgTbngQt4n
CyMoomnyREd1p81c431Voc0qYBi2dpTSe7oGfG24AQPQ1pndMNSXxEJ8aUoLvIA5
y6gX85ffZnYSzq+MIUIQ1HNWK4+9EXP7AYuCkuTjdVWYcCRi9QfpG9rDztF6RSXH
rBwfJOEc6KUGlrDc7kDihfwsiilfG3l1Aipwl/8DPYY4wCo74P+Vj0yrBu9kbqST
vELSGlF/r+rTy2hglfJ6agiiBqpO55RqUmggcAz6RPaj1OpYsf9egofvamqyNwhU
dH3NdGb2CTyCsXkFk5/TUbF7U7nsCohXioDOnnUAZhUKe4VBO0Z2sdcMCYUXL8x1
Z3YV3K6XDwSDFw4Iy5+CYZ4ipvg1wfSbEUXdMpJ9oV2EJ/0THb5XDGgWrUyXQqU/
U5n/4AnPd6SfRQR8XOO/gQW/DRfTrQcOkorXhe50mcXIyG+cv+5ijxUnD4MwoxWF
Zsik+fy5MWcfp3qUyylPhbNJMZYTPqS5mqfZc+SNJSul6nhLfpf/M0J0PdlPNZ7+
kDRaOB8oih6ASoeiNiIMXNv4UglvSSuzVIJLxrbtJaxIp9g3NuRMJuL2USsykO+g
14+Mj3ZfhNxFZclYdSSiDNEoIqNoE2zjN7Q5XZGUh0IwPFWXmp6cGvso2EpQwR+S
ODQV329yPfFWYasyy6U6C+xvsuSFPZdc8r3Al2ZTFS1ICGEuSlaSHdUYz6qRil9O
jXYxNlGRLiavJrrlo+2wpDwZ+XgkLivsAR8pcqrRP+N/OXpAKysJfQ4FP3AaQzlV
bcbxfJSshUFEtpNubi94V13GNBsf1pLQm/tqZIzuhbcDYxrQwQeFJmbxsc3n705O
UXp6g6ESzkbmc946jCu/ulh489309HN6NxeaHQzWbV4PMmFsPSV9BzHbWgADIDwe
xhScbkAnMkSvI4m5v0p+Fe0+cnuBGYm8ZQG46cmYgmCerqSGnmlTqeVXNTpwFu9U
nPOrhGdOuK/gUyiNVX3wnYx13Trk+/PpXGC77pk9A6as0xqZf15aXiHgDZ3wHqpu
QTSYyMOh4JCl3etMlbrR3ird3j4+jFSMgc2PjTEqHacOasbUJhP0V12nAXqzW4JR
Jhp7j+0t8gEkboL1M9Hf193GKZrWml55dbBU+Qss9pKmtxbxNIYeDFNUg5VDbHmi
Qzres0T5bKaMdO6CFDf2xhCxHvJQd/Wttbp9l0YWx8a8TEPZHCQuaUxkYVEOt5M3
S7WwGAiBj3SpIiZs+XQyeQMKf9CBIfmpdYaxRgoFWfBdb7/k9CREjmQ935Y4x8fM
5DyQ88/IPseNVl6HTJMbGnllzDuuq54G0cx2ibl5s6rh8STGlncURPgJEqhPe+TV
gZJPoPBqSt1sAzr42n28nGs8xgma+M6EI8IrYRxIXFrtAxpHis4LS9cax45TQF5v
pX3rU8TNzJfG+VC5H0iG4uaQM5UYAI16FEWN0CSo5OTpFRyjT74wMqKKgeQEbDpR
eiW1E9uI07epGQo4ZWZL3ebI2SLPdYVSGSJkpEEi16VUms8VMbxov70BknxddbRQ
tmd38+NkW6xjx6joLcWkPaSIGJto1O6TAf7Pk9gAR7iThkc5GYPyDYBX/g+f3yFN
nHsaXSZqDpGH3DMyuWMkOplfYyYHvD0rAcRB7lS9+lAVnwjmcOYmm2OzoavERqJb
AzSMoZg5TfPVUs5vDYzni5wDG9gLDPFceA040lWM69/Yl3N1BJ8Ls1I/lnsakPQp
d2kw/u9072NpooAE/HfRPO2uR6ZFMn87kLkni5TBFcdbepTG1clFayHqMrtUUg9B
WD5txGAtN4y0mscMsjzFntZxwf3R5sYLcHk+56IBBRhM8I16kU5E3XV0p0GtfhXf
nOSZ8Hg84T1W6tjQzMyQvfxdYhOgdbblm6Vn1NltlQE4h8rtPCvQQs4s8CH+5h7H
nR1qPe7H3zgsNCo2Y9fsvgfvGB88B0bMlUUoqwyUdOVM0Zp4FBOFHT/RjvvvmvXG
43fxqHMoC4eu2dUOY+Zq9I2+gSPIHS+LO3gZvo8+cdbT8yQ172P9NgHCDDuBFk0T
0I2HTyCaqT7zpZ8Nkm0kHFhJzWpUoyov4hUOUjH9Mo6X8pWopGja9zb93OhZo/T1
i0cNd2zNWmhjypiGu1kbzhLHjcqrjgY91Fb6WbgrF5PgGjJ6nMqLq+/jOW8aGRNn
fqkpNWe8BSTgPYw/OjJTLtX+655qo5sqUZgq7uIlbWTix4U8Bkyz9U6U7dlymYQU
DPMusCCfFunn8CFlwDdIYpjFPXyKVG9kou8FHbstPNNOA7yPZ9cONBiy4RSfzO6f
FSBpbHQ5Y9oeT4jxBwESkrHDWxSPqg+wHELPtjdDUkAFnhRpzq2a6RLkxwdMqqw8
PWLFMViDSgXAy9JD5JbDmpcqF33Ut6yLUbktMbk6czbiwikqRBb5UVssu6bFsN/e
GFKjxznVmENtDoeLc2QNACgi9u6TmCXw5kDfmFCWhNMTb4Arrt2Bj52hnkrDXRfI
y7pHuOHl3gWkgRAi0UJz8jKu6oErGK/ewagYHQ4yhbF5RjIp98932FbovRS6lzLp
jV0AXgDElbV9c/XcAkkyxhCduYk4WFUBaYV24yiMWkv+WJZUyxQj9SGBnKTae2Ec
uE4Gjq53Gq/gnw19d36JReqwT8y0TJYmZod0kihuaPZqGbcB1mmEK3y05gW1cnA7
zFwQ3SrjqzQ7icg9u3Eb8PHRx0s0tHZ8ApfeHwklKtoaB2n0N6m4tVRcGlAHXzaT
mj5RQPsPoNZO6FQadb10End+Xh3z9tcz9SM/W+nvqDNJ6bjzKtG09vcv/Pt/W8CV
he4LFNLX8fvInIOWJltrW4aOLMAVfv1vd2A3CvwQUvKQGNbfzbEUE8hs4suM9ie3
u3XFXsX3xsZNqQZ0iHUnx3ucB+WuACLJBJpOWL3C7riTyZmPzk1pPC+Wzbd3200Z
d/LCZLKawe8DDtPyNmyhmzAsEAnC8WLgykEla9Jw2W6kwD/Ld8hreRp7V/s6um4G
c0i1e1BMcv17J0J/P+FCLstZ1LXaCGKadqXEv0flQV8YU3OpMl+Glo3aRkw0pXBr
tAT1r4m08iVxDaViF/WGi3+7K0J7efWC6wZzE1hcOPgMhrmG+ytVvZxN5ofIilXs
kMOLfF3W/Wh2M8k05W9ThSAdzqkL1TdWv/diaFoG7JbQCowyh6so6z+KSBnonGdm
dn0eDAiV/9xVLsR9Arwle9Ul35PHujDVNQsx4GUTIlqGlZn0nhSndSnKcRbQoJvu
K1wwfJDmkJxR0WwYqGkZV2GQLhnxNeO110lzU2iEu7vPZjYsoVu80CxM0kFMm0nS
wvks+lO6MyuMYGX8OrzSudplu3d3u9ZjKJb6rlmkzIjlGfloWVqXpzCG3VtL6vGE
8Sr2nxHWfabc+PNuI1SfVnU7CPMbmPgb899YrbYFwqXNlR/VBf46SPB9x7pRUiI7
XP0hy5JUTBOEiBHIzrSOdOjsH9VfcXH2xGWgoAjHWSeviZNZQbjHzpG1Or8S30Xy
4E4u/zb5HcrUm2qmJUDDJE8g0Ht5w4BmacskA7YDfRY5R5EhzZ56j04xrRtnj1GZ
gdh3o6IGPGph00k7gvY7GCEbgzs+hCGfXUswiXmC3ouFopdx6sGilriT7ucYyhUH
g1cbH8MH7Ee7CmvPjDWVgptQZMHE6UswBc3NPJr6kdoO/P5x2Ka1WjqmevzocNNh
fIB/hbNR4GV5WgVKLEZ7Jtx3s0NmTBuLHifuioZiyDiHvK6tNaglqtOLxDngsobl
QYk7n1sLmzkwK1H/dpFi1IW2oKMYaDaujqhZ4ZeiYLARZv381bUDgGzl+diSwpmN
0Lsk56+Skmbg8k/pMn/mVghoLkootC1If5I4/YB8gN1n7STs9NMVn6PIPSHgi/Ol
yMtJbY3BA3zoP/Ij2Ca5MU1XSSyXjK+EUYvufS+QeJHR9aCRK/h75MJ1S/BlfN2W
l/LPu72hJZSB7E6dQE0LSeyiTRj5rcUPFw5lxfMJdKtwNwI9ATkOknC+KRohIRms
GQzXIn/X4nN2xC1QS8XhoAj8IeOE0dUqrgSJvaJBVp3hg49WY5osagd6p98DyZcu
FT26ItxIrIWZTW+72jXJKllZS5Q0OShMmR3EK0Ajqu3JDQoUvyPp2KzwosCboIY2
z1S0vvCFLx5fACVtVkr8beM6mnZKin6BCnBBiabdXsi8rceOZZAhA8olJLFFgw5U
zYSg+KYuIooDNBI44FOdvMRsQ60nW/Qk5+vYGR4DfdL8tOywQh9NZ1Os/0LND05y
VCYB7MD4xxjZ+DAh7IkwKqa+mrjTDiqAKH3Ldd0Np7xCYiDJSQOodQEEFrCemZy/
s2frH76lFvaItyTM6HumIHk895L3st1zB7Tmi+X9RZPd81kHjc2lT2+/kjdWZZwC
0+3uANhbBbeShf8lDRELb0CUn5d1KDP4wXRKcWkIKInk9koRGCY3AJzOFW64NWDd
mWw7s1ydFLqEyFm5VZNfNkyxzCOgyWhLTwvRaZgTho6ldED1Tq6wYw9FNmq5bjUS
DTBtGfrmqV1GvoTy7hjMdw03QBGe7DwrdmlIhE0GVoaAD4ArnZXQTLi6UQUrXhlW
KmB1nwnC1iqXVh2Itjm/+E3PRJMCDtoVh+sNcD/f6QxmDlbPcdm3Ey6e60nIiC6+
fy1VEF0GdCrKL8oIKokp9G93sl9n3vaidm9hibd+x6/vv7sbWwzI0mqmOV3r0TPN
aOp1PfeDQAsitUsyRKHNJagsqCY64JR02d85ELSTUZgXbeEtbRjIdMke3NGJdUQ2
HX2/5I8d8DNZnWXbHRgR7tauDffmWVihCdONI7SzrKI9H9N2uodpbHoWlDu1a70F
IyiJDkQuGX4zGdpABZjl5QzgEUWAovZTLOzIn9NGcO8hQ3/fzlKxAm052qPfDxLK
3w4WGL9UDAT1TwywZ7j4H4p1wYx2apWXnb8D0WIdI36Dpd0L1DetRmlYUjZpBbyy
39OwlULTIAJ1D+kcWRZo9AgoQhdPIkU57nt34EnjzVkI80lj25g478AMziZl1/wE
v/grLUei21HB2p/P6ahqqlHwWrUpOYtnd4DDUjoByi9SHRVOE1n+K46ijuWGaVK0
lXoRciwzN6T0YL5kkeRK4E1SAuLdA5G6iHBy/z5YU00Bq0jGob7pkSGsm/Lzg4oa
+sxL+bE0JSDgF5NlvHE3a7V9Lv7+uF5jT9YdHTGCtOcAxP/ahASpplJaYx0jxlzM
Ag0zT4n7aOUEQzNUSFj5rc/3jD/2IznK2Hlg+0+dO2kieteTzohZzLTiFZa0lZXU
TW3OHdEmydoYdOhTcjdaw7/2ZtiLE39tR68CytHzifof00OUrlz4YV55+tLkPv4v
2t71H5TABahYP5Bx15YJqOE4LC3dzfqMfr+CcLx7uSdFwldz0MuUtK71BMPaDMDC
Ghqq4PwSHR56tedLApiCDUsKTswHEIqjnhKE0d37I6M3FqiVHvoOkhbPKEF5qiSs
dQ3YvwQmL9P3clDPopBMnmARE8JsmYeuVbTPb5BhVNIm1gBTxb8mYs+06k/beVYp
UP7K2kFz01EoD6bUVbcc9NJLlTZJiBt3OxVt9HwGpno0Mxg73bNI9nQtAP1zcv0R
t2Ysyq5rPOd4eO9RsTJX9w/CWYzyOkRzvgF04dtp1NH7hDnVCyIwxzEytl1A3uVy
UgjrXuhGdc9YiiFUTdRDXQUC7jeTvR2CFdVW3HO79R+hOCB+KbNq1PccV/7q4Ecv
xo4Z/k/DIygVUv0Pfv78ntwPnLTdMWQjjocL2mZyZeS07dQdnRr5pfh7tdh60JQJ
JjoWq4eZvIbDUNGDT/QNOYFgzoQDYYS9u9rdP+5yNgjN1YZNT1COjS3NqPT4fHTi
OJcPeGyblt8G95zXUYlEXCErC09atr0dBRVRaZbpZlBapoM32pp2GObY0z+yT4EI
47nqGYNxWarHpF6nufSwZjH4mKt575ppbMJdOc5Yx1pCyipf45S/cAv8C4Xm9gMC
OGRm3QCYD425poPkRqcHbFSOGsG3U2w5uphDculERFMr3M6vEWZ4WTl+xy4/+RyG
zsM3X7xP9sD7VpAQsyk+f0b942qvvyx0TDkboavhShF5OIfPaOzb5R5rxy9jK+0y
kB/7r9QRbCbG9a0s8KKVVaZgexyz1itV1ZvgqtdW9+ov/lKFnbsBJO4w1fwa6q3h
U4lf/q0OQZ/E1Gya1+M7hyc50BfX+Vwi5KKl7sf46HLcBrWktXI7PKgIlDuRj3ax
+0a2bGTHpnBVLV1UWwjCwVnuILIkui8PaC5vetFsHJukdW79Ij27ESmaRTm/KnO7
OLqsCldL6rPH73uo+1C1dG8cvvTOvGYfJNxTvk3yT3d6bdG2rMnCttnJM74q3EGF
ztA/jIKKkNRlk0XXQVqTRXrf6vVUdYcquGS6XHnNYfJqeoYoMTy9ySn7geq7H7Pt
fHmUiK42WacSsHhZpx1r4UCjzNziumIHBQnUcRA+HMRmXtJ5yOmE+NLWd78EXLqD
Uubxy7JWwssWW4Ua4NlP9vyUyacMst07M2ssDy2TavgbKDtUMw3RJ40TosMjUuxJ
jxesgSlCOWSgNvKo/1PHe/rwxYLfRY+xmqfcLDZNxsnkMUPwlLwwk03QB6jSv4II
3k4Wttq9g3530gxTQ90PBJyuZsoCZptJeI3BRlZj0QTku47uaSMyL3/PpGfPDo3z
DGGPV89VZzwVaNxuLpbIWRr2nttXyeovaDeHjRaIQPNAAx7ad5A23iducAqZZJPb
3T+Mhr9FGkEfkaTc7lTNCEt0fYZHereZp/TiZHJcciVcVvwZzpTeIVooxAqZEg/y
O/WSai+GyI4WjamHKAG17ZojLPdKUI0IdZLS8TxqJHRy0Ctzw4s0EA8MwLCQHGFg
nORqBs2NCOmBoNQJ0ZADpIde2+cwVx6k/0TZeuZ+3po5f9frGbAn/qbcPdKkHyYh
xcKdJB6VzquCesw4SGPJo2/o/i+UqXkME41KwXqUyeUIZ4gPz5+hTHwdBdDzV+5i
GapOblpp0hjycP0fJ5Ve7kbyL0K8cNqBdbOd2k7jDWUJEtRwO5p06JhDPRDvnU6P
LVtgtmTyh9K8p1RMtNJA5bLAyNSWLCzZx1DNoxzMbs3sr9tH2pKbmZ0yoZFOe3Jv
GeWL1y2mrQpUDwdkQLFUQvINPyUgjCNYYSvYeYZLYx+tOdtXz2f7wEWWWg5P81FG
7gx3eRIqyN6HlAIZm85fG2YvOLCw6E96OXplGy2cfqEKgfSve5psJrm2f/nC+VUu
2C1Fo0XZ5WnHdq7PnH/iR+PNPAnvGJSEw7qUeV6YPqXGorznmEHTMNsxoSMPxM3y
2/2Eu7nx0NDZTy2WFJSAxro4Qpt4EDZRVdMJmUTAC1dsfg+4deSbdfPmFhAIJfCt
68kH+rs6cjglXmG68zZ/VTwOkN0uDjTYDcyGn9tjWuaNg3Lhuc0g5OWbmiv3+KsF
M6lqA4VoYWER3qMGPbefLUsDqRFi6fr3hIxvGJ4Z2rXHKfTjeJfxI5qQSwvL3QLm
rLj7CHgOiccClnvx5KCOaz0yUssuW9PCuipNNSKEmW2EBnHeEG7HnIAd55MNUO2z
oTAJGpKPgiz2N+8TfyqTfwcrH/qry6PIE8qagVspdmKoX8wqwLPqIowY7/qAACZf
rC3liJpyKo8VZwtVULkBYsmW03c7O+rgi3DL+cO8NEvsA1DAACzd2MSxGWu3HcrP
VJkJR6/mr/azOrvo45q04w7adzo1bEXDooujbXchsC0NjE7VG4fg46XcOkbWV3iJ
Nx2MQKxGdNPGRf2HLsdp+hNdJ4F+aMuRuMLvJx+ihR/UW8+2loj0X/2COqK1CvL+
ZXWqbWoydy8JxKzK7/YgBvFCWwRP/a2hwfnVcm62Y8HADCG4nvub9ydlTRtsb64M
A78scOWsmPE0XY7PC5jD1ZOGyEg0LXPk3MVLuoQHCby1pjjxHPNzCdxOgaAAEt8T
H2yRs93bBoYlY0Omjmdf5n4hsWrTYWIMWDqNV/+ym3vyQox/P4RWNzH8a4bOPU5A
2rnTpYGrDLCKhXLFuL74i2IY3+HiDYeRIjVaGIXgTkxQVHG//BaRvn6qnACXiCz0
/7VLLGdBqWKOMklZjoohakHaSseJ1MEXaXrw1bk1tLO0rbmSlaONqkKNZA8NZlT7
/lRw+umS/t3mYo/bHZAKtinstyjl6KNrYlJq529IQuVfOZOSrmeqDDY0VG/s3oqV
RjI/uWMMVhhtwKGm0M4P8LXxOi2p6nzwKMVJPZhNfFRNcoyJLqLJ38pNPdGfKzw3
F8vWhyu6itmHAP1bc61FkvlDs9FyUpRwptAa+Lyej44PR17arQGKHTj7ZnAp/GDN
00sPlysdbO16c4rqx3kUhZ34F9lPhnf3vY4r+2DJ8GAxllAJjzGI6Lw6YzfdEN+b
ls/zcgaDnmU+5T/6XOA/wqDbb4LKD3QCf2pFgviHab0lyjVz8rQITdP3UgAbq6RQ
cmQ3X4n2Uk2gA7JzcgMw4z/wbBqpWv4w1U0v+uTaQ3xKZ47G6ajQ3G3IZKUgLXvW
FdBvhF7EL6/l9LwP11C974BgU5Px/hJCgWANorkr2lRkyyu9CkUAH6C5P+hstiwk
ovuvW4bP3uoaSX8ljigKfxlp9aCkRhPXnPZGhJPGd42C1Wxd7dlhBh3++Ztd/hUg
1P0d+Nb3mVcwh4kxG4LoiQwr6Xde+bXLjKMnrciEqKuCFSqep4utdTP0iln9D4Ie
cXhzCgSa1s6Kcx4Xk6+POkOugfplHvAek3pc6mmuW+fMJAmtGMGTJAwXVy3XQFep
lG9Z+2Oc6E15z0MbILogRXNJ/LyWf4Td8JJj4adx6CfOLQyHvkJFrEyMeQsd/9FO
17u/LzM8rInBTiKK8FhcPThDbSa9VcrnNAs0UrRRqfNhXvGnA5g4bodo+oVYTG1a
2Tds7qcMO4k9DmXCGl22YwzbHjXlcFCbF2GuoAKtEQr50Roy/NuwquF6SocKd/As
1x8aJRSwNvrDBIE6EX7/KxT/7b1YeKmO6ZElPw99Evceh3yG7TbIKQ50a09pM7ri
v8Hd7qRipJoIro3avC6yRvU1WI0rigRl1JA55pjj+mGmG11ckm8b6zuqTn5v44HO
fSW3J1M11s7yHX7j4K0yfRyTZPjmfDwP6vlGAU5CvRSONQGhb6WTHNlR7dqT7NpU
Hng2LOzKeJnIiY36jKAk4k7EcfDazaNUTsVVguSEsau3IjRxCKTiQQ7prZGxntFR
QZ+tRdJB1fFbC1bLP/OIvO1kfKMgspuEv5lW1BwuL9bfa2fO3B43rTnMLpr+1wj0
5BLc3R1qi31uMuI6WuCd0V//G7BQhz7H00sHiHYrHWlDaAnwdMM7trdIQRnhRRC7
I5qAzhtK7NCYIHj9bbvYhLRZErXn3CMfwXH+ms1shPdtH9n3RQZjcTo2vk1IeSJG
ITWZOAOhRLmvcf6FiPPbIyCT6EPcKlDMMqYHuvTRLfNWHcCD8uIklZXPyZCcEzqo
ROk1G0deJ4wRSGNTqjfZe5fSsGA1/8zRqx8S+y1mqDSvUZDtOfDCiCCwHC0lM6N2
2qB5XYAkUhsxo2t/h/DFLNtNpHpm5Na5/a0hq/9EmQTe60FuxiS3s8EL7NRJlGbu
rNgc+7MlTjQLVd5i4TZxBE9U5iTVV8mLY9SxSuFmis5Do9nEIzOygR+JY5SvIn0c
83oBzX+m2gdWKKHLZuYgqZdSmbJlKIkW+XBy3IKPyo100st4fzh0mpz01tcTIhUi
+YIOZCs5qI4rL6wEj9mpxneqDNiwIjWUu2zXxRyLZ+6YtcARHKD5sPzmCXKixto2
hCNrV27sinqyZtUie8jhOEsmVDHM9yBCvAgoQ/3UlgdDxlFaJQUYlWoSDUwkxUXi
ZAE7ZsVzMdVOKwNzbzcJaSEg7qB6WwoEAWLiWSWUrx+xgqY/rBi+tlk8tTR9Sc5s
LF8saH3VFJYTiCthI+XL3alXO+HXhGBvHFdLSQQMw85fnswEV7DJqs83p+QKXIa5
aBIGD901II1Ai3I2BbMPTlP437jSvlDtanl3srvXBeDoN2eoLy9UwxVud5XJq9b+
eHYO5XX8D97c1C+ACHesI3+80d2hiKKHdjzgZq5gSAYewxgL1GIIahWhyRebVSY7
dmxDSo5IquW7TemzndVrWNH+pQlxwPOyYtMk/o225o6PZR7jsbwieMPf/Ilo5t/W
vnuti/UV78QcW2JyQxt+alrtstDebagNJZAEcZEKle50kJHm5tjB48lBNQQc/z0a
ojEbhx3Spr/3dSru4rC0qICZZNr90CQ8twEBAb13RB/wpFfSIs4KEiIYgPa0RIBN
hOvKPIk54Bo2dDlV+/Kod4VH1bfht6lDszdD7fHAP5JFANsnymFiXcPN0ESdP+IG
L9OEWwpKvhP0sWCghZMYD2alspBE/fviTw5MTgRuylOs6jB1eVBvIjoXfcYyCfJf
7FYikhDECjQr6kkDvyHpAXLRYcWYQ8eHMlCNbT4cbvauGJN4LaG6I9AerBcBpjVn
ZGUWHb/N9fXnHtfvXH1jtKGiwJokICXFY29weHk71hKITikmAdwsWKtF1COIAQ/3
fth4zl8uKfB5qoTM3A+xflt4UQvMX/glUen+TEFlUJeeaD544NDfXZ5m9LEzfsby
EjB/OnYn7zhw0fku9puxL050tHnWbBUXcabJYnvRAQhUCC9Vv4NiBE59baebfWXl
5jE5CL9Dc2+AaojBnvsqEHuIiIBrXq7RZyAatPH1Ctt+U2ebQhnsM6YVseOnuBAy
0OXcyc73c8FdlNgBO4DI3WqGxSQkqgfFaM/9zEfcHfWqC5XGo2chTwSu68MwN1X0
Px0SZ9rVWjd8Mro3EgGP5WZqcgTOwq90ssyCm2Fo2kHfdnpiU2+qkilrSqEtQIyV
xqSB05NsH82t38ePLUKL3N7MQCL8OeQ13Hct70nOaoviK3ymeGb2f/nh3wMXqIIy
QQcbmDLVpbXwg0SeBeZWCp+xE/UjZwwd5mKHEHcywjl2msXKTCADUX4mkLfkyV8T
GJYqnI3X7yupyY8OqjlBEWcLqikMVtzpsnYzsIzNZgdrsMJystciGy6Shwi3+yyB
0nPrwjObrIHnLF20z/Gkk9lOva5Y0Nb1Jc5Z1NirsN0hZ7MS7Sea2zakevL1rV+O
C1KABU0jRYsZneO0AHavCsyMD2OvYqAzq4qnijyubo835ANiP/gooGT3wW2hxEqW
fjNivUg4h1BO3z5CELDfnGojrxyhTUnVyY6GTSY641iW8QMQBLE0VI2T7VkkErlT
FEeEAIMln9eR3h5F1ccWI5nOeHisjVBfmZzcaf3M8kxSbc1pZhy2n/bEbpOEfU5T
T0Je0IlnTMDuFROyZ1+MtmRTwaSky/+fv3n/cDq6hf2kpLLYGrJOenvR4wVfkYiR
FdmjCWfveZjia7W/wVfhHELBSAV2ALIBrO1I3Ya+RKRPmP4RppuQmlAq3fAZ7dt2
b/Of4mcZK3SXxxIhdDK2/Ezly7tDwvekquF49gi66b/2K5cr9+GMAFD8gomckjWE
oXv1LAIgjewTtYmwN96RIMrB35aFjnGBajpZ+cEVxFMZdPqhsgTROW8wkycMWnjt
ECGc1+usQRidajDWGh6YMQioUgvEUHFIg936gzsUqc23/tLN8PzHtER5zMZ50K0O
wI671nn//ge4ZGRvEr036a2cHtcw7RA2aqqyqeQAQ1zHC4Ajm0c3tv0+yPBzK+tE
kWrAuy2/AwSCzJdS9gII0Pwi+w/Q2eXXbk0+vTDykxk8GiYcR3JUlNa/EqIwu1Td
eMIuMD2L7ujx4pJt9LscH04hqfFQNaWsNMMJEpPYoUsoBPQONSAXYQ/rb77vfjIw
udUwoG2GW0aP/Ivj+79Tbr5EL1zOavhh8J6UMZMKq/U+Rk6OJlhEDWHpruERu6BT
NxHczX/KJVL1KAwCqpTEMK6quYZWuTFAjPA3So7z+r5KN2U0+G1IpQ3MCmxXJZJr
Lp8G2X5BOFeTBeY9lpkk20xf2xUm6dChCnySTAUQAZ0Pue3X0Qa4H60bLJklviTM
ORIMzF+g/CMJUkdW9phDkgjXwQVnrGjKRthswjYEwd5VtC/VGupkgDhseInDhkt6
Q25Tws+YanM5Y7h95uywHHi3vpHrog4+r79fee/cgMZPOsH/MXseXTk9eN+DOE/q
vhfZxF1dDC4pbzLy0CRaVgLxQyr0vBlNkNSpLE0G5fAM8HZujpQaiid93XyQunWN
CGl8Sasphn4odHoJQmbBeK4nlDCRBBT+1gd+YqT63A3ki7vvpsxXLCo8uTgWw1a1
ebJurDz5vBqLh/DueRX1sXkzMmwpkXr4mjzw14ZIEfhTbv7/2HvWE2ylWUjjlJCJ
DSoxeQ8Xcpyq9MuMLcPKmRSr2I9bfRXCSGrbD7r8eut+x9Ya0VS+eb/gZGAUL9Sv
ptrv2FM5kYlsQXInIv6jfnW4zaUjl0bN2qJyO8XOG9I0YGmLXNte38bvEXIQUFSd
nDYgUDhFLKb/7GrESxXHabXee62Uuc8/cHGWfs0iISOUWWcYL8sgJCo20eN3GIGY
e0hBjtT1a40yUCQYcs0jscoRAaSV5/r35Lm8cP716pli/a3/0RY9VXAMoasQq4JQ
6ApoTZd15AO7Femqejmqau55EcNqQ8QfPazflWZczUYTLIa+Nmj/4aXwfhc7oZQK
bvV/8Osf92yDXvGawLWEZ3NBdGBTs2MZtOVMzinBMa4KsZVWcs1Mcxqz8ZrbIY1d
kO9w7rjXN10XcFAQHFEUF4aTKbkPB714rHvRnwF1030nRskAEiVI3nctoXUjfP8i
94wvEuF2l55DTeIU7ag1v0HeSPTqxSRBXs3tfMMBJL0W7eJCdN/5PGriTVFcr+Xw
IzEgsjG/4bH2+7UUBwNs8qceE4J94qavxF4JXx5j80Mkl9+yumh6sjHDOCuwJNFR
shGbR47MyQienNEH0s3l4zc3Fl082TEJesPURQ9nq1Bkn08X5Vvw3MJ6pTik5X+3
rUivPnSZAMqeYNqqxdj6wsp3EUG5hCoUBNSi457XRJyeEEtrYSpRiKvkVsamzQqt
Jw3uXzahdWtljYTSSVwoYakfWQn4aSHyJeiNg4H19F68h5vHTY/b0x6jm2Am30az
VYZaKyMzalMrfvM73gyjT4qo6NFEsDknXmMcgMaguqXYmuzrzx+rvOrh7WS3x5ir
wsbzkXUSOienhZgYQnoCT4q/e5iM7wQK+NCuEjsizGD/Qw4piSnYgXq46L/D/OT5
O9kutSC0G4Jz7qEv62kBlknW9Ot3zWA0rfWTXrdz2E8KH97MCws8DH8FDSmXY6nT
gn84iy6LH7MV5DM7NE378xTtLGgVUpEupJLg0/W9JL1Yljjy3VvllajTPCatPyZx
vnBBALsDl4OftEN2LuEBREErGuO83s+dFhL/OarCe01RzPcIEi+qFOe0QlBoOOyr
XWYdHMIUhgJfqiHpToHwJzo8hINYMihJbOEb0/wcckUAkonvl6Bcy6jLVVfECLrn
mpA8a49vm/VDtDUpy02RKNjFL6RWZ5GWq5yparfWtm6AaDCnZ6uWD5jB2B8pI8d7
lhwXVD12rXlhV+6TVC1QWrl4/EgLWv3nIlaR0KAaxl6wrDTTZZakwN25SlMFfv2e
iekpj6RYbjOv6Cp1iGs6cCUrVbdCjAVx/vwseyiMhJdYy32Ooxu5AfaV7qTP5VeI
LLFfAQib0WEVtfnL3slh9zKi8J3xRkHDYBGKrbXzKSxUH1pz1dHTf6A+2S9zE4Wf
mC9Jnwh+5Gv3PUHCrUrMHUJmiVvo4SCN8DBpoz9dYWw8txXKrFnEno6JSfAte5zn
wrRBjYqTVwaYIMMkIgZ79Q38xOXgFUz/3nL5D3sWIjs8yMRmfF8NM06mCIPtvHDU
L7LZQ9bIyT6pbAaZ3yAlafBsKwN2cmFzP8OmWAhUJYRn6uXM8jjPr/Upu19YAEDI
UvoqVBA6g8E+9iYUo5+YKSDvmxwXIE39yXvOr7P/5vrw6a5cUxwZdq32nkzGw+KC
Qu5Hj/YZRa3Mv8I/CS3i48CTOO+BisDbQdVVdnZeuXrhmMAKZb7QbJlwRWrD8MWj
ocqywwROEmhrjbJ5TDlf8/F/uGttEbnbF0k1SAs4CP1xOXIkwVo0FNk5lqhXUwlQ
m5nWEPaennv+TkvejvKBE8CY6SI8zka5sduamM+KGyCTEafhmfHhe/7gYbO330HS
YAL4rYCpz4uOkoYMalq4+cTLpaW3ZFG5kwuuS1kzBp2KHD4L3lD+fVrx/BqTN7it
lHstuTinKjPfuW3R8Bch+dc81X/WpiY5JQ9KhR0tQ4wCE4AR5O0xSOLYPcZTXV9R
UFePW+lX4VjDwX/CyDE+5IjCKlhljU+MMBD4ow+1bXzTsyySzaj29uMEiIllk5Qz
KALL5aceaW2yfq+N4fVtYJR22miSZLKBXqKp7d/vY/Vg/vOO4hwu2xk3gYqTf3k3
xDRuwTlGFNrMc40T1fvGocx3lrLmhp0iaImK5SM+WCeJV5RaDPso5mTc+QI2rf80
I1kevzqZwE+LD3Gzep6cxJewtz63rCSjiJ5ceyRoryeuXokszQnrIVS7ziQTbQLY
D+qKHDqXxZUaehGgA6X5FlGGLD8/8NZpKL5ktZ+5mHrqztTlsZNNCJpF+QD12moD
u1lbUhggseYcqE953+Xi9SfY5v/HIWrW1BdAJUy7adfPow0e8U23cnK+ls4aOlVa
b+vsMlaL1r3PAgCugEi0zte4hccWUbHIOQE4rOpVRdLzCbeN2txkKfovLExZ/JF9
woEBr29G1410TWbaLFydaEvyXIPrFURmf3PFsBiyT1Q6+jKal8XhIeu2TqbgkgfR
IVPZn6hWN7AaAKL3fcF47VlNVddnhW/LV0J2b3Xomwd89UU7peRDSzNFZTmj7WD9
IG6ObpIgFm1Q64OayQCQpL7ml5rDrd3DaOa1EIPEb4hjDluOlRnnF/z9wJJNK98s
RGcTQ/ShRV5Kc7LM1JKoPrmnNCyHg9H8EHYLt4X0BHo5ODaje/dlbBEz2MQV2p+n
/wbhxdPuObrzIym0ds3xyjtLCIqUrXR76nNxNPQj3YJT30AYwALb6sHi4A8aV82b
DFKmkcvQfDX/G9Qcwn+Q+DhPqonZct7HM4wZIeH8K0DFHzDKPOVYmidTvTwcvdE0
hezez3TUi2HxU/zF1Oeu6Q1DkDGQfsY6udz7cIlSEJB8h3gnvIYTJK7H7Nm/N8HV
u3is3KX0Sb5C2mlAgZbdId2/c8STphUL9xAa9Hzld0+iRjXo/6GdTbHph/IYzIJM
MaPKaX5in8FbXlsn+mP7EOZyYG5E8toc6ywrYtv9dTzS9OT3e1ipGV0vEYFEmUdz
0X7//n+P7yNoJfFbv9zio2SKZJRjCogEECc8vtUNZqyBfLICku1I3GBiWqbv5P+/
3QcO4I5Jl3S90xt/OPJAQYkzlEJ7T6GL8wlI+duVB6vRiYWnqdIZ6UBHhZtitiPL
c6aG7K6hXlffu2BgymwpYdyCY/VIzGrmDQdb5a0fYiYSbmTO77lV3FJxZfL5rsCz
jmR4eu1XRxC8IoMUaFKsmNy2feuK3dcR5FE2yyL0NFhJDExUZO9bmUsHdZHghfz6
Ci/MN+3SyB2Rd2Mv6UddfcJO22kvlPZAmG3aUSkdlMvP7wVCkOBvYpwkrzwEMuhK
hUrhWcPxSgsCLGVOmngpzb0OBv3tAO9mBVQNovJVXEeB5xzeFZSiD4xdNrLWxxS2
R8q+zMdQM3oigTk+vsTneZ9ACIIOsdskNPSZwphaxSORvWlCKwuAPm+r/td3Yrfg
ZZ6ZTyKf04mMp8b7aMMpC+RZXHNHgyoM+LgR9OyE6zR5x0bF8U1lxraZtopOKV2L
Z9QMg7TqG38EMXegKRyfY3jJDV0dcjR4skIZkPsbzS4HqnhcML9TITjgjHj191eO
gkx2me3+A9D9brxTEJC54IzUj/jJsryOz0dOHs/o5ruzLOOOwgKY8RogxA7BERWW
tyJZ3sbIeW9ZLbdnTTOOHpJXRf7+VJrsaqIk7qUvCcbWzJg0V6haxjJOW2NC6TZC
cKVdZlrKQG4RlReQSEKfg4W2dO3diWb4hPDAsoSbuTUgBIAOFNIVjROkMWPCu6HA
tq4uLEwQcTiLvWQ9/gsMn0vOqTMJ0SH8HusEUJ0RRIe41avHu9Yd5CbKlOCthh+9
4mSvv8E+FcTV+8UHD30SZf2O2qDOmHujKOY37epUJJ9wl/9kzEuhI1vg0SJJSuQ5
E5q55qUT/vhbztD9SLAMLRYIzNO1Yq6QsPVbAv5c4c8li33xvoAWXDOC0XWFF4Si
JllnDO5tmy/5NQSW94xy3VENkzPu4vf/YQSKuKyZ4aMg4B2jZxPz1YLzKtyZ8kUE
JBohF/u0nYfPTxRz2rMJs41IfRj2T8oIDn6TP1A5vKRpn9UzdjEGseJ1QDu/Ay1t
zWan5WD9/qyoFEpdo5doKazWP/8GaecPgLBNh7TPLURNBqjgA6zZc2P3+yEb4kfc
nheKDrQJPUclKjAdTU2NcuoC3ssjpMvMy8ZSTuSMfiSm+izbMdzCUAtH924HgGoX
I0cFQFEkxhA+zG6euZ+sKz6B4ipIqFg5Mbq+MIDU3ISvkhUfVM76uOeJRX04+ch6
PuWSLIPD6BOKNFb1Y6Uc742s8YHmBFhjzeOUMAOpkX9wGPb+Lw5Bj719tr+aDjxF
YCkmnregq3kf42mtSyg8+9P2K945meCwro2ik6SfgUCS7XO9ZDuiTUCjvZijczhT
oRhdmzl2tMx0lEADx6GP8Zbnekd1c+vAZzxU+TeDBdEOMQXUY0ZjRqYTOAtQ3Wfy
VCN5TBZyuZwovAn/61a2Oa5Y6wyRHhfF4Pa5UqKOiTqvmwVy9FwfvAnC6OM3r6zE
Bmq7P/sLrvrp3s/NkB8G3KIMsFLXXfuJALZuZTChFGsBNnpp5sfHOfGsgUmcf1nv
22cVGGtPuPLGmFfHOtsWyC1LzEy0psShkelS2nDEuYfr7uIYchPwSjcfcHCDWKfu
09NH86vM+hzkzs3Kp8NGD2611UlCHo2RiZLb0oMhaeTQsjkOQvQfEpXQCWJMi3tj
RuB3bmm9S5FXIo0wIzfoNgCF+1VsLd48sYNrELj/cTZr1sr3kf3Qls3b0frraK6R
y2NvdPcS93oJj5ruDjY4hocMIvPQ/0JQwr+8K2AEhjYa0uCA3wsRFeneknJIEwxd
g+Iw/9VUOuzepgWCwzXuO4zBXJPpEYri7Jwu6zb4Z5cq7fvNmHG3s3An10t8x6/p
8dHNsfSTGC18ECEubwB1D6ZA1PFDIumLqWesXXQ6pEheTjG70lGG/ZriNKZ2D8ss
CPd7unDIvJCpB4WByWZnxoGs6uJGfHiD8bcH0xdrQETbsYnbRcK5nJFISSPS4QYU
D7zWyFzjd5JxIC2mmY5ib3E3F5qJJXb9QkxVxuGnbzPARkwx4A36ojoRFfmBamN6
gIO528AMQVqm06IvGWHdRR9fJn93S/B2P4A60kJEgR4b6miGMV8qTr7WxNZJ4nTa
fuZuNInNjKMe1/PSvUgDCLnyvfWBOOuMtZRygkkefQKZmeQovkkl+XSLKTR4xKn4
89vOeYnOOOyqPJFVTheFF8ItJMAo0LI8BGxMDk0QCVi0qju+lLn6DVuim2Ysgxov
jeQ8XesvM5CLmEhj8p8Cm3zOVbP1KESM9lMG48m5Tayt8QX+piQ7R5FMoLnn7+SO
/6R3ape3JD9LxQBBgsrj4xTktd604rydJRPNNm3t0Ncw9pTIXCKySlCTAhdeL2+i
rnmsGl9h7whOWCgyDTG6GE657MEd0DC0NXXe5eXLT2TKwdJFh60OcZMTGdYdngt+
tBGgf4+N5G/RM1GL1oFkRWgfFJyRyJV9YaOhB+K1VQUs3hK7C+ENzMehbeCknLiT
NYIJwJFD6ODIN6l+GWnHPT31Y1WO/Bh/BHFuxMy4PepRmCUEqVZS6SLpOIL1HVBX
0lg++JfGpfhUiOkQ+/BReglfaWo5uFrO4BBOkcCm3lNN0D/75JLa8pgMUQOCIQmL
bBfeKxDk/kge7EseGDWd2VW2cS/7MjWfPdWdbuAVZzbIWe88urdmbuGKdRve8s92
o/dHeInYfYoS6lckla11R6LMo1M6CMTqoZ/KuPQhp54u9GIayNKUvoklYhoTpFLq
7jrxKjwtg4jdT9iN5VrKJnVwko8+jCAvw2paxAh9c9PCZCjAzzsz3ASvXhokQkZ2
YRBq4LehNt2Q8rYQSFWRzuGKQemZ2qnzAJ8H4/R89PJyYXM6lJdfRqHwc7E5cQ4Y
BiAATx1wP6ztD1lewRSl2zk+5n5zOYxhdJOG87ZRwuqT9X2RsJW4h9dsI8F3X+sn
TTyy1pr6O97DVeVxttqUjXZQXZyhU9p4266+zo9xGoQmPZZNKaHHaSrTDean5HWW
lpAG4X0di4qU3h8JXOdgl3QuvIJXT/hylJUZ5FTBi8j7bR+aEi5S+2/i5KV3Ezd+
DDfZ/TGmTnzNnQ383+x8g1T6iG82p7AKpotQIry10KkxxBOLWxUrF2i/dNymY/SX
0ssrrVyKpj4Cc12gfveapsdvhg1PeIXORe8CdeLq90TWtJsJLd3xgxPmMgv/1Gkc
grtIHo/nzssZovTT75s7d4J5Tahv/4aIgfNdTViymRbPxH7BKFJ6eVM8sYvCVaZq
Aq3JbOH5I9lOp48pmHX40W9jUdo2DR/eAKlkl/aehiJdm1A8Jk0ghvo8AWrC9eQE
b6X5tu8MJsZg+b5nRGw8ISSLmPE+tepqpPAum1fAlI8C9fsFFDyq88WQoTbGq4Wg
OI43LB44KiV2Sgr8aTEOB2RAQKUcU65v56bJqrRGgCpj5Fv8X1jCcuSEmEbMARZ/
93UMNRzYuI+x/xWasWSlAOD+mO7AoZNgh3aVPUutbr4WjXX2YXnw/pwrxLEdvDyo
tq3pTEJxvW3WkHmP3A3kFf+p1zSyEV44Gxcx4SWkpUOPW0jEx3CFX/xnPXzyQQ5e
ayAHNRyZ5CyiKvgsMORi4UrzPphdo1DxkrXDiAoKPaXq62RpfyLY+FEfGesmNBsB
wNSpKNC6hS+IO8EyRB3FDS41xQayw0Ov7kDa7mLsjvtt7NPHyvwcQxW/wjq6VkuU
sbGwh/J6B3g0yrAG6W/c0n+AfOHWLuklDLwl4AwU7MV8Zq+Vppy3OUlqP73iWdc4
yXQBytWctbpOo0x5FXRTlV8kNEheTlhYDYdcVKbpQil5d1gEVBpFW0w7/nCzGy3s
ug2Rdh0PZh3VHwkasqVtTb9BAPqNoXL/56cSQzpQNqdBSGeczwtWxKSKpF+tLh4I
v9/OIOrQZINJTey2kTds2BUlkml4bfzvqy1Tj5MyJ0wkNfmAPl6ZfZLexWn4Ct97
i6n6lB+SeOzK6GtsoaHm1UPSoVCzCIS/1fBk+SKYCe4TciLFfQfwqX1NrQ4jfo0x
+twi6YzCmlJ+AxWOSTuBEwwpz3GJdSuMDzBfNWx8rEvm9YMKXmUV3vhJtHiU8w8j
IpE9gRbtGfVlCwZxQZGyYl76W4Suj8BKhft3C2mnTAiZ5IqxkB2c4ZumniQwcAOi
CF4S+37L5WA7qkApUJR0cQJkKNOH7nAz+vor8XNNRTlx8loiCGg2KVNsu3h0G9dF
qo+67KcjrUKTkirY9xgQmxFB0q1A+7CNkFc7IuOZgEEBjCiyykbnCJakhjT4QEZW
tJTcqMulAhlTn1qZEMySKY5rcbrhOQbu8RYL0Yr5CIJa1TJgdupUDR1u17BLInyr
bv6JSEk7UqlhTq0Klmqe0uGSQD3SleLnVsxZ1mgF042KAsaLaM8trv9e0KWKHRJJ
nEjENH8OoLwj/zq1Fj+rp1rLE4zfVR1hLvYwszH0WRVp1Zf7YjyYHXhNoz+ug5aD
MUrr3JAGXIYpv8Yoqlijq999yN9V9yzL3tpUZUdIUcoYTqvhiHnoxQh8ycvDKT8o
p+iOKtIAyZh72FvQGULkYn0EApcIVAoPJ2Hu/mGkRoJQJYe+0+iNkZ7mqaE97mcb
Oo82ZNtDgtBBzTrFwleeNjLmdN7i7hXDUmwSgiY+Ud6CBBaXZjAtVULqGs/cU6UJ
Y9O06KN7W3QJ5G+/a6Zs5y2SsiJvbT9A+UPNyrV9J5310fiLxybpvhdijM9LIMpw
t5x28W5YWoyah+EWLP29UB05GN63n4xkz0AZ/ODVCwUN29xBB/T0Yjjns+AXm0ii
XBwre/BLa5yvufe4TnMqtHPX3O1A1tsFC2VD/OnpyNaSMg2MoVJ8rhY7bV8GKerM
CzMMnWmC1O0RWYkj28jMJhNxzXVrodu2Le3OUB7o0O5tLUN0ZIl2PtwI5YNuKiHk
YNAklRnMCI0QJbGjtfIWfIDSqdtfrLGeMYp1fH/dSTUgn4pLx4MtNwDhYZAUSn/S
6dGlIruI8h9+EO/xCi/itv7V33K1xB1spEJU0Nq8uJ+B5aEMZkSyfYspqEtpoo3s
NaXS0n/5OBQVBh3rgmAvdS7wKnPsIA5lBIXYCDvzesYhavTSxi79xQbXfjbbgI86
5xnnIMtHaarOGHWJV4EdI0bVu2CqrfFlotpvUqUCXOoE0+CtULUsBAvhAqgrU+lG
j/SZ665xmSKnN6JXO6LDtcK7/EYNTr90V6J1lUg0Wx7zCyxEjymcjvFmvsF0NxnV
GhLDF6EQnF5UhzZGfFua744Ed+dxREe1AEV0NNBU+VT3npv/F2pGncXVokHyBe+K
Mb6J7TWX3ygsporjgZ44QFVJNH2Zz+/aHaYkGD53TihADliKH8UPc0senG1rsuk5
X91QwBPM+adSvkGVvFjkofTpZMiGXOG04nA1oEI8XFPEyJ6cAkGIcK+WpsG8zYmf
iPcZv59rUFZu7+LLbpKj/RUdqtF9pqicssqUPIACR/GwcVvvGyNUjMxiA0+vG+Pq
w22pr2b9N5KXcVCFKpO5SF0ohruIUqcA9lyD53kZD8IGK4LDoFka9+jP3R/HjD4h
S6WamRxg4ThWer8Vdmlbf8arxMkBW+oH3kgb36S51Bnkqirg4ZxCFdzxAARpmLnh
ZYGmAycnXbXz8z0A2BIZDoJZjCre5Bnxl5JEbodpD0yLb3Vt02rFgwvHxVgHi0HB
52Z9N//OepoS/jQup3Fvzgz7/I5WG/3twWwl6D2+CfXsXx9TV18u2ALY7mTa2lxx
gzfMhlqcuJlfHaZFUAO+kqTq8xnavRam9QqDHacv8u/8la6qyrWPh4ZikZf4+DZs
oA74c+h40R2xIvlNzu0Q+R5rpM1RxH8YEw2NlHWN10WQxxLTIvDmGYxO0ymi8UUy
wsDLUmvEfoi+FqqGMZ9no6FRV3OIaAihcixfP/zVPtHXz/mxRm0JXL6wA6JAKKtf
4yxilF1Wq3a351AgJT9q9hZYpPedzzTB2OTZ8wgkTdpxvjQFz+K9tf7o8Onk5eAq
LgLj/gp+JEP6Nw9qoP0t/rX7bim38vuBPXtfeD7bx8fMEz7UBeoA3spuc3CnKqaa
bXvIAJ7z702cflSw/XNGog0zK0ZzcvYjfnSuCSWWHZJbbiOFOq5++p0ZfUiU5KUs
b4roqoP1OuaojjoSQLQePFTDQNX2ImjMM9rboaFKCMcrZQSxv9mGXD0aBbKSxqUT
uxUjFtpZgNqEFCVjyFe8VlwF6QK2LwgwUNWRL3ixX9sniV2cIGW1kTmcpaAu6Vep
kRW2OXqjSoWe/faFg9P6klo/bLC9xYNi5n1bjeFZjPUrj6X4mvgNh4sNp/A4tasq
t0jF4HFXySYEaPsBFzktgB7NvRNdQBMIhwKOYF2x7OMhqU9NqqGLhaUnhBUzHZWU
w0TRxzWeIWGAYsBdhFNQgKW+OIvUtQrl4y//0GkOZA+1U6QGPE0ww4IWrlWoL8bJ
AA+CMkLqU48amztiOGtN0flsy+zjnOBlwnpOwF7Sa0UlgcdQfVkGsgtlEPBumYc+
5ZbGwK/A7FO528WcK6iLmcuofelWELsSPewSjTu2jSS5+X1vkcNq1LHmuK4KrqIg
AJh02VGI11P73xVSNn4AfTEbP6eiwVkngVzPXjDHUl1FiRh4yGuM1wLibc1A5htt
TS7FkMPJePUKxlMdLAIqr7beTeVu3JSM3x03rJLlA7VO9ceU2Ho2YlzeeotUlcwA
+2yztJlEvOVowf4FqUzChpcTcAgIghGvQvCGBPX8H7MbowENlbb8A9M6UW4SQe2q
utn/N0+c1Lm6r9hDB1LD2/rG6xYdNnEYmryMJC9bNRPUQmPlL8gMI3C13Q3cpQ51
lnjt6qzDj4Z2eYOcMFVBLP827rJfd2mE9GumCsDG0ajsYusjtlreMpOqpDRCXm/Z
qO1sAMz4hpMsAUYCbpJ6z6uFRMl93Ii/LNmr59bVHJZVFqmWowmIr/sDRiQHR8ny
RvjtsPvj39RTvp49D57P90M5/A8cZEv9UByMVB6l3wDb+l/Go3oij4+XnIJUrK/Y
4z5Tu1RWKM73WAa0oHuDe+LzcdKfzDFylyF8L110f59SbucenmReL7n2qQYmyI+B
iE/Lzd5HSjBudNjdyeboiq4o4wEem6yIWiQq6OFDGAsM0L2GUMbF7PxHZxA2goWr
J9YbwqSPjE7st72UDI5RasPhZ5rqKBZmRyMOXkNf8qhdnz+m4gFrq/UxPc/ocEbB
ws3CPLH/UEeN3vI5swLXqz4mSt9A26VW2SkEFUFPWq3HBfm2b1cGoeFDOcTCufV8
fQYqZJuG+hSf8EVnVVlt0k+RMMFnVvQbPSfKm+M1B3+tGZNeXngYM57mdAIYVk0x
ZPmyHKPoXQDM5Vq/JfUckI6s/AccqeKQanO259MsJVh0yyWyTLtwyunf25XrkU3m
9DNwq4EqemYR0Bl+tKWWftewpB71UdS2gmF/MbcQKCPsYNuc5PMRbxJ3bRiQIqTw
Xg0P112n0aHCctVonQlVzpe8b7LqotL4c+i8sXGIvvKoWMpIliVVK16HRipKGg6H
z0WJZ+8u2h2jAS8KGs2d+9ViNpua7VALCLL76nKY/gdDYDHiFJYWzcWBJRE0lGM6
MY68s9DV2nYQjs5FmdPRlL//wda/t0Mrx0e4tJb9DsSSWzHfwbe2KNuilK59ORtS
5ULBDRnpaiB2faycLIQhyc++vTjLPZe0hifkLrZZRKf8nrAMM/YP7bxeu0gUNp3n
dqqzSWIUzBG/pZZDSFc1goxEPh0NTwBhWnt3X8RciutLjK0BkycYeHIGIeC4hxgm
HNmMKMQsurtl7TUpnbioCN3UV9l9L0wmHGPK/1a+VczQIGo50hEZDl2cn0xI16HK
MMB04dwhjL4xAXlPjS+BQF6yBHnCu3ts4rlpD6WlHPVSOzub2008BvxpA4//MpZs
jNB/ylihYvQXoMcLJN4gn5DbnlBzuDvVjs8X/rjhDQ836dsGG0oCtEg5Iy1U8urG
xkLWRJIJoOU+gtlBJhlkSuXULNzJrHljKOZFsHn5j2WFvxioLAZHyWBeV8SelwyR
mAZS9UDeaDvp8Nf1JFZda8641BHULW19JIrBDW7IJAI0dRf8uhSDDpfM2+7IHpmM
0EqMPbiI7mkzENEQkDRhh6lodIWfJy/VTJIs1F16z5h4mZTZtwqnDA+SWnC9MWmS
DN7dPQW0JDLP0Uo+ZPNOZWpt6dEcok9itnC3ccRsS3zMUwz/YE86YjR5zZGtsonT
1Wf/CNhnDT3Vma2pSQuIqI1x1LYG1WdcfEEIO+84IDdhcph4w5pzLl/lT/qzrXRl
wBfoiys3xkKEpbjhULgXZjjIS6WAtQCTDauK7NSpyQMDY8e9uhilt0xpZK1vmhVS
ZP+4Jkp+glZVF9w79n9smkK7JBNouCjxK6HESM2GYlgqXybJQn0Eu8nehDBardWf
n6deQn5Qm19CIR2z37B0wanUZ6js3R9zGxuXngroaQb2IISME/U4AmwRvA+ppK5M
aRGYjIIfkAgu9Q3yDNWbORyxWuD3y5E6rcVH8Rqt2WgNGoGjnTFE60cJZu2HPtYz
DyMsobhGdu5ia86KCvIk3QTp/aM0lvAVdTVY68SXWxurinQ4c3IePwlxJqhHODff
n4mR94tuRJBz1oG47Q3SnPJznLGO7devYMmOvoV232N1BTJPS/k4+z6zDfD4UtM+
ONuNJ7jWeBSDp8QlXqpPIsXUFWsczWNxwZl4ZwhRiHY01z96qozLx7OL63Dp7mEs
mnEugDbMWjriYHoAdqs4evGO5hcb4FavROaHBYTuYgD5XQaHGGLrGKatN1jXd1kK
JXMTdSFt6fim9olSzr1J8dbXe82ym0Hyu2KjllTsFt/zaBJvHW/65R5WAoS3w/0H
Hi7eeoCoQRnAKcI4bbPZkS82Grq0xl2urHLaK+q6DzwpAuD+BRNUi4M2x9/WNC2N
kEhgqnBqppmPvEshRwaLztzn9uZufWe5ECVb/+K3dsV5drVBRFJ+GPa8uP9K+W2G
F/0TOn8EPNUubPYuHddStsPvzw7jMjXlXRw6Xm1ZlgV9hGrRPt+X5s410R5aVAaf
tMzzrOlbVMahx1QXWA8u14L9HdXs5ZDMb2mTOM/W0OOvn7lKArp2hLwRlav+YKsH
GaakOY8XqNyL/YTGiN10tz0thWTI30FBDC96oMGLlcNUGrCn8fVUNfUq/giuDpCc
InI3z8jsxICOPWNbWB6tGCuLN4qu+UEfRzMNUhRuB6j4CsiV5SD8Rl0tGzsJSsTb
Sft3yfs3aPIUIfVgYyA4lBU7qolPdza+Mp4oPdhIC4u5X0H2m5QHRtDVffLHX+F2
Y2113K3xKTDR5E9xSxnd+gfa3tSGYT5IutAzEnRNHQR5A4VUCICirCw8Ke/Cvo96
826wGJ1koR0+sdyAppwrBzQtnylkT1WiZqApz3XSiVzPo17Eew/6/+c/t7eh6LJ1
o9Hs7PvQM+/2D+DAWSoGc4oWaaQzpTZs4xqi0ntNPAKzmSLCxGuKnWMGhLGGafIS
5tSDwkOrHxi2APLZPCNNF5etLlrzthI56H2E9IrRQ2atFlTm3fjxMCCzHG8oArZr
m8Q89Mji0CotkFJmt4RDqBDBFhaWdiwWjETNeycbtEd9KpoMIGygYlVRKAXrGWq6
4cLF/toRgsOoUZDBvlHzyhJ7GrBLFIfqCniNXzOJEujlOLbSImRio6I/mI/FkL9M
NfyX5Bfx0xcAfJLyINSv1tFQA+dAuIjJ3h0AqsRiEWT+GJeZkXWGqwWA7xLtzWWO
ot3r0GMrxxIHxmVZhsJXzSvK4rHha7RBpnB7S3vfKWV1x+AVI8QUO+BZnOdS9TVW
l49OSl7Aihy8P+ZUbSWa2O0FA72MGVq75d4JTSI8elFdrqzO/zcZEWjFP3EdKp06
CN3hzU2TXSQvpOv+EOdxUzlNjKEP4ltY7Ypu3n7fKP0VFdo6sj6waAqP99T4pRQY
RQtxB1JrXO2RiaY4PedYrooVPMX0lANeXePDBOck2NnA1wD72NxQExAxRPzyVfSY
xKLM5tv/v+iAqDOMjuZMXNU8SCfazGWEUAiRyhkaPOQJNpuiExvEBkDwIoibzKaj
h5XYslnXnYD6GE8p/YzZE33UR7TtmHlVkgRwRbPkJvjsiraz8tTBM6cwDYSSVxEb
LPTMoFm2q8O+Z2chpvTi07I2N9wfmAwAJ014n+VMvwQzS2D4j38/BY4kiJk63xz5
OTS5vPfFRKWCWk4MTn2XRA8S2/yHTIBQ9vnHbOqKIGhvHOP5FaQ0PxURdx7urfUw
i6dM/af20POwjAb2bt7F8367mXuUv0lLY0xIc5ADvu9t7ygZ8rln4fvv3UwLs6xM
iXJOvNxaAMitR+wkJ8ngUSGeH2WxruXM2E8PZe3k1HHfdcTyEHuTGlG7xubvVaUl
fu4glNwQpr4tv8+I+w6rqHKv9hI0J0bxPDzqp0Ujkxz8hKZ+MJxCPTnP47dW/+eU
RWEarZVc0Lh0jMaqfggowK+iKyv01HHDc3lThwQYHpNKg0d3Da+yNVPHSnUGf0NK
/tlYxyqCE2yzH6KJclz+1XQOxZtshHf2N9LQanaTaLXIFOoA/7RTFS5ViRbpxp0N
FcmaA3kkZJ8UBZcK5iUX408IGJtQEi2Q1WFC+NPyHg3vSGB4RUBq/n3vEKxaiuHe
JY/oYjSlW1b9ZUCbHdN6DerFnBU1Z5TZAeLguCEBHxI+WUCENAsBBlDQG8W/yZJG
j3T1Usfc3jW9sXqKimtJQ5j5LS/E4bM7GQG1w1asMV5ioC4pLxSj0aVD9emTR0Vm
LJbbozGa07Mf34xNaKhbQmUF/4YUT2bjC0ataiB3kfKuDcvQn6P1A4nIF2KpY+A1
LdLeT7VSHiHU5AxspGSMC0Y7NvHvmK4e4Op/7+NSstWwJcLs8RVo9+twb+fZ4i2x
GY1CXXnLSf+Vc43Yb3jhZ+PCdFEGG63b0GuyGdKXuJfUsfmPSc5NkNG+hM+YHW/z
+xgAupJ4QN4UoNgRbr/l8y10I1t6+xf/AN4kvLypynRlLiZzlE6kwbnn5285jdlg
aGpdYTJFdivBXmWgbjPKwNeB5WK8KdsCz2a1kAI2EAun0i/5fXI7VUSMksYOqVmv
+kaZ/IrvTSPkBlqopdeHvZgPP9xfTK1lNymvsiwpEa3mqvwk88vIK3x3Qie+uqto
x8eatB6tW0TCGbZh5TvFRbRXesW5UiTbRnTxdp4Lfawd2E1uFPrBNUCLxmAYE+Tc
v2ygk2Sg4NwYkNmU95Z/V6n4Vx91G/ELzeCWML4Jb+szimdJAOyVxEoluJQccH05
cDCYuUfarkeVHsHIkBOrcE1E/4TKS0zdqtu8qw4Y7wbSWnmcoC85pgyGvwFwTFjq
DDT2xUdQuMROFXi9qZNtArmhs6hR3OY1/J1a3auPn60QrLFncbHsXCUvVM45hZo9
oaMohSWKNlbjIPCDrM03JkdgxlCZu0nQdSXhkcbrA9kzo8/BbkdYEyV3R5co+g0Z
lLyU120zMHJk/CJ3xqiXDQO4hb9SGXA4lXVV10yTyzzrfrJReKOtQAkouQKlaVkV
uTOyQuoefAc+pp8risAUYhCbd7tsvugSh5Bu38L2/jLMJaB+AEm6gtn+ABpnCrds
YSVo3+zKhlkTt0g0/wP7g3dcdbWZ9XtkeFOoPBZiPOBAn1Z6c6R5jxDyyFdqDtgB
PQn9XOeoKdKo91UXu5+CPmvm9IdqRPBsrvfeGjlWd2HLXL8mAnaE1DUVhw1WDbpw
nbb6qNi82gHWKI/1tSVHzglbb2T3p6duIjM797pDQmUJvPh6qwk/yLibACmJhmc3
gsh9IXpARkkyM5UJ4PhIJU+7HtW9zJlKAYc8F8+LnYGw02akQIMWCf2GdfqAwSC3
UilFexGCPD9taFMuyr0ROwnJW1spJ8p8lhkMjgjjRMqbN0a8b2f/VKGSh6jBwzoG
qNHfef7W0AkbzNOkf/xitZet+hkRJJ4bRiwMW7KfMj9T9t+B44jxIJHhEAqwqzhg
3WXjfMADHk3/hNcvIAVjxac2wydCVgaWRQjezYCjEVur1TwtlHATs/FBQGd3Iyus
apAL6wR8NFJyry5zU/vL9jGYjaYbNdyvyITQEhdcARADdLdDYatelSkjTbZ5kL/6
pjnE5nSER71i+l++/Z6LlRSnwNM+PwMhn6NZtQvOIJBoNhrO5Y2hOUhEx1s9ui3H
6r4g45P7n7xzM88MzKi7SiWVDlh7z+Q8uUN6cNKgKezW1bGRwNybjBrMmPxSfvm2
NqP1IdJR/YBi4J9OLIFIYFQ/9LvC2+sXM1nYVzofDLI0/m9zbGeO/NO3WAJpJAb3
5V3QRVQyUsjY+0hAtWnlJzyjcUoR/rvhB+kogaQxArXzAn3e/emJIYbKytCSY12b
F7LMwgfyl/SWcv7J2lW6Y+uL7ZSwysy6WpOzm3VLAaBtIKHu3rGyT3rxijNcI/61
zoMeLeSZO0OKVUmkwyeXEusQAkDVtXbk9j0eGsMktaUL6ygTxESsXf6RqOLfpYvZ
gRI3PA5BnUf605oCyR4uEy3ceb+TCamvPhH+nSF17znBQNwUW7yyDvJw9Cq7hwwN
G2St93BexecYgiOeeJNDIrwEWrcudmPduODpkSmb12bEVnthtYso2Ynto/4mbtZK
ooSsXYbJS6fQ6pkvbXnJXHlKCQkkB3xm5tj2nQfsdZlVXwzfccIqa7PnK1TXLJqB
I2YyuV/e8sE2mil77A2ldDnje4iQn3isUK1wZcvzCsmA1Qb+eVjt8Fo6aZO7ARsE
HCa00oyfv0mU3ADZ4LeBbvI9Mb6QyVdyE9QPnLiGgedyO7R7IaFPtGGNwvpVR/gM
ZizHBOwYuSkOfSUhYBEhx45GvPitebhG5zniEW/+IxeeVfxU0hjTFiBmyhf7XMeq
lAC2HYbbYlms87x5QtB7u/C+plFrG4VmeMACWiyaa0ea9bptW3UVD7z2a1m2/x2e
S0o1BfucXtnEckWdk6wRykaqBMqpSOBdqSUV/d3dq5SvfmZLiI3FNZNjYGXKuK6G
SQbU85JLbmn3ykwrqO0L2sOiSuBfjKC1DulaTgmChM8q3YfjGGQuEfE9QzAij3V8
y9kBTi5ksAOuiG7WqxOxsJ+6DLv8No+2yDD2kKM8W90S5gcvQA1TBURTwuc5Jn58
YciPDDKWE/hcp3yMQbz8p9/pRnJmwy0qKBI76gt7dFR8silnqcTTO27k1qtW4hEb
qlor/PUVd1xK2k4EB3M1ArhZQj+7D7PZwuthXQZHiWFtVhJbnHF0BAOBh7zKV2tm
Jk8Yo/Uuq1xKcck6+tD6sWs88NbL9Gt/256VY/n2Wb3kzlxq+zxsNA9yn9a8aaaI
yVnaZpHU3z21wk9i6VlGdG0o2zasY0p/Rp9sGw6ueLHzQmjh7XKczqROjLut0Glr
3OSFDoTUOPu/+7iAREAIDy8owmZ5LZXwxtj4JuLH9MtEfCFZUDm5tmoYYeCBIN39
nlOsFgwIwFs/0yVp0kNCxbJYssHN84PqHa77VDMvKkZdfTjeoheVOeE+MnseAQIh
Q+oXAOWMcPZMO3R0hKJ6yoC5sqYGy3r+yd8uKpJfD/gZCnLsaxYLsC9h/6DIjHei
gyUxH4cOZuqNq2juN5c0iZMRK2wfdDWOqubS+JT7wZdT7YquUR9K112VBaiFxGlx
t5FactV71UhglNW0UHYOoHJf4gvSU1f/55T/kcA9iYV3S98mfd1ShY/6pDEK++sX
FY3EEVsS9RoixVoOKr25AXVtS7S4LmUSjZubKNXy3ftJBQobhAZndgCDxBQV1wH3
sB2S9uo5znFndXY9Rtf2y63BxbcnV4GG1pYKoKlnKU+UzCBbuZ9p385xrYFXZg5q
dnQEu8Ro3s1OWrTlPEMwttEwV7y6Z+ca8g8hF5/Rq6snx/2ccXKgwm+72E/3t+YD
pDLmsNhjMCkD2ZRfuglhE2EJE8iC60UZUVk2peY0kz7/VsNBJZeJfy41n+6Inguw
XHXANaFohjqk5huel1q/LoIpDFSLJmpCJmn09PAU/Qr0oFi9NQZA2NXsSohMZ0nd
2L4TjutOevBSQeurkLmFJomptO2/YkTP4tvRVMYIujYNKBH2vlPGqJ12LOCVfrMZ
e0UlJ2/obcN++Y/X2zTvNSYyJSJUFYCv7viOIHicCG3sW/TbQdEBTlwRfNQmAS30
BsovpQPvXq4yzTzWu7L01fccrKuYFlpBySrX5Y0qs1+/V7NVsamqcxl9YAD4lXGP
AyK6V9wW2BkBN3+dxX4KFwUPXvLV8BE7XJIDfT6xO8d/NMacNJVNzNmG8Pm7EhgB
7/YPzek9oSJ0iiLn8H/32nort3Yk8pbnvx4e3uyKDyPZVD3dPnci4v2uiZS8T5+m
C+m/EYQXuaCNbxANOu5B/hJUOd92A41tCHhGQUDJxGg7QN5AXD6yTFcMFjxgEdOC
2ARLdUAT/xuq8d/sMoqACEhoSVf3KUy5xU3gsDbJ8gJ2NIWOA/eDc/7kL066j88y
pKW32nU6RkrPyEtQsglJJOnXtJEdQtH6GR2TnxD4XmB5rdufYybdVsE5nj90HAi+
wyJszpekvwMH79krtMWahSMVaq2UzwlO7L0r8pr1U9kyMAMtqGzgQUsSSsdKrUdX
L6mjbFb9fFLgDyoe3GQsfktZSfiAwyhiTZ4GTwUbzmjMT1hYQyklfp0kmAH6ttjZ
dgNfMV0NSanjYDeXbhWomtc51YWHW+WTk2aKwuQ83jGUL1FwikbknNMtxntWaFxK
XrRlPlq21GDBOY/9peO5Lfo92EA45w4hhbZcpoMWokTTXKBzvvMBsC3HBI+KuKxF
ReoB+URpBHJRG+dwCSRAY7QwKjra/Uxd0vMfIrJ8LkDbgZVXeHDXKfw6BpiaOPbT
sxyO4MY0qUp4BgY0o1XeKwQ7je6pjIY82UBENAkI7Enb5ACAxz6vQDiAhMNcZScZ
lCv+YxaCThx+soJdVKapHeeHIqB61pQvD0bqMYrT3FGdDsga5arxhEhC/AhVaLq0
eKDWdYrhR8naIMaEjuCkM2ujwfhQ+XNwkpTc5U07H9vA4ogCkNQ4QIDrsZFpdscQ
8TfZzR3fuPuq8eFppC82GB4Nq3qf0sCQeR/2mdnw5E2Vf/F2pzKH0/8fpCZa5UQ0
kZEeGKNAdtkWwll+vDOl9spZS98nOGlcCoUmmaJ2W6zDLfyyayvQCbZiK4aVPHuj
TFz4ZS6CVkCXU63+wV2pvUpzu3O+3Rj46KAcLk3Vi3uQ6NZSWgcWyiG1twi/dkMJ
pWfDYG+8qVwVDVgODg+4myDFH+8UaFLQ8RVwBYTCyHfWYALUcPGmQAwRn44hJQ1e
fsIcHcpYoW+MFbxEG54nGDDSTn9umBsFOf4CikGk8elVRAp5h6Q0ACCg5F78ulHj
y9JcshSwKcCYbJfSZU6jUBWukhPkHG9TS7MJXWk3tQ6CTum8iY8LVUcEzOkT+N+x
AzBmyuWDsvSXGCFzNPG6qys/KWZavrbPz29njhgNX30jDStNQ8ueUNLzkXSen8ip
Cbukq3wKOcXzkVGFwbcWsjj3wf2nE9azsxMv/06EjKrdJdhQ10VeK7qiFdTbL77H
1H5L6k+lXqjUOeEIdrd3lXAwKtkuEYb0cAUeAahckXPRC8KNmnU/iqgTHHl2x6rD
CYZWNUmEZRotoKI8fObeKM/R9cLVFnPb9Qfvj4rjL0cdqG7mlyt1xd1xa7aOwPQg
jR2N3HDhUIECr1QoitIKVod6f2Y3K+bTvoLLtxTzVlooa0Z00AWP3pYH6+fuKuJA
DFDJRIi1dfbaDny03EOyGwkcg1N2OtUcz3YxbvaW8u6ap2RkXQnsLE4slVzjBjd2
/fh10a73Yb0fRD4G8hINWEk7vsCFjDjhqHbAcZG2rSzW0FiXMA+JtXKL+Wc0lJr1
8Bfc5lncYnWNvNdrWZcLP6RGUx1iO3ouZDR1EpYZZqL7q222Gol35ArzeCRjYnPS
rE/78eVc/t4JPbdBM37ZoVvh59hoSoQcHjl4csR98Nw4PTOaZaFwxix+9MOpWe30
8QmaxxOlbCdgSTQBhtcXdoDsSJzaRQ1MDFGJXhyleRFGpYrSArwSqjMXQDrYggaf
D2WsskjN99OHtHE95gj0B9HQta0WLc8ONq7A5jZrTX07H6LCKGeoTiS/MSyY0i0s
9/njAlBkEZ0nrN0HQsFAEEGe4w0d7D3h/sjRqceSfbKRdwgWuPqDRozYH7xGMO12
KEr4VkkXDSXyQ3Mu+gySVu5oOtts+zibWuLrWoYmzBjEBnnPeXStcHkq59YCGjZx
VxWderW79eKNy9QRyR4g/NJQX4TYhiR9CBaE7tthxWSoRKA3OMaaI1Y3YTvNd8Yx
1bybUfIU16fQqyWN5vjtMOaUnzoW71y3nAhT7+r9TKUgWtnNO2RaXE2bao0g6ydd
MNs4XKa9mhWIXqbzQJbLTAtetJwQ3pJj7UBuq2GFEw5PSsrIUbvhLhpUz5Y1nAi3
SppPfoiquE8MzEEl/4xXQBL/lY3p4fGema8C623DOtupFQqFdEIrIZ+7hysOe7z8
nu0RbuNKJcjpSt5Xd3+I2lDBkRVgsfau30W4YTmmBn/rtY8tPrDo16dM/6F0MtbJ
7INboNPJFIh4e8cYvLcN5DvTLUN8qVHAKPaG1IPSp2HxTuWEeki3WJtuNzjEX4E3
Vah9QaSG9lXUFn7/JQcYIzS+3s8V1QtyY+HCqILdTNI76Z6CM2ZAthY+t2Hz8+4O
b8SmT7yTs4jt75RGwHMLTeq60zKN5WjbzFTQWCm161v/FKAwLj9o7kU5259rHfyT
+twtw+cjrxkC+5dDTYdfKp74hq6UsD9zHc6yysSrXslCbMs9uj20jGLInzAFrCgc
623QL4gYh/7OrunodZWGl9erDo4yldAbiAm0VeYwdtRK/Keei7BfYhsJp1L4q/yK
4xhvdlQLEe4Ekija3p2H7YBhCUI4h46dqpetVUzr/UVE/lkY2KxMmVODpYmbnZCq
CKZRoHNRoJLBxjR62w5foalIB83AczqfiLC2E7f+pu1TMpm9DrP24kmsG35CHJmR
FGmfWrXdUhn3VfzP8Bejo3n33tbx9grK2QW86S7ielky4/97ngkxVya+sDHnvCZU
bgR3eTIk7d65n+vMuk6TaDlRtBJFik0tt6r1VfQ/6lipkvtKtRn84opMtrZtUA/K
wsXSDPPSZusvph43FYO+B2alNZFu3XbPa3OClbPwREbKjKbDMYjajGLejO6SKRmU
K04FNH5+fqjmK4aAOELmwo/4d8BCrPOWa9g0oIR2DT3lmZAPUNuIkG1Gzh1pPMHV
mk5fedzi07WLC/8DG1qkLfysqXaq+Hhvc7uyMrVc4lTQi6poSrF2y+cvbXJ+HSlb
2oQFeMq728Qc2pVf06Gy+KJwRpRCYf60El2ayDSSix46y4N/GFsDJvCIBkMTc1un
YcKaeUnMAK27k7X/R2Qntfvn0vOCwu5voMqvoW4XPmMk9OIKY+upicZytGoFV3c3
lbHYMHtcSO7ui795bbWvfZXPYUlrr2GgzSQA1PjLoOw9zLxYNcvbmHQHBAO4pD0x
TfVCYVkFinTlPaD0JVpRkrAm5UiQjklT0nTOQHYLBCWq9iCMn7rIkYMXlzsPKnqc
JJa/W+FEQ1LiXqytHBGgvQUNAE3gH6EBD2EKT4VgvfzneHrP7cwt5J9fkvpAoZt5
Lw8DQv+g69qD8FTXO4dGUn51gG+A0F0GXylBtGaOHoJBTLCwKUdd4zDd2RqxaMI8
Y6jo1oUc4bkqB/rQAZJ32zb0S1zzYuqhchJTt2IWtgxhGU1fp2T9pIhcobz8C/jo
TOyzYpYkOA5Gvucvco2m5hdQHf72um4JkpqrXSSuq2B79MVEB0gnM1CpeSnz38FI
zp4HxktnjXg+ZA1vNWt+tBsoT/lX9NX/zmnSuXW9NGXVVixpz3z2rf6hVHucZ4QQ
8E3ie8jj39V0BZQvwp4lS9rvMwa5YLeyn+enmGeAVS6pZkaN0eZ//TEU2YD45+MP
feZr7FA47ZhiadmMpobnuT/niqMes0qcM9DyMOwytYC4xeIzzWyMQFPdyZ+nT9ZK
u8G3v3ye4SnJozHaOU567dgpWAsL9/fzj3QtfpR4wjOOcVNQ+JUhqpojTCnWLKK7
Jbmt8WtFf0yAgBWoG2QqhIqKp5kSDQhlIemlMkat7qUMvCYtwdSRhER5V2hcV7Pn
P/8oDD9mvglGKsapkeufnAZCx13ByaHJl8DNlM9HoQ37GJ+GJR0RBJ+RiLQbEjMp
9Ypf1U1zpZIjwazzMldm2q4m5MftX7dT0Zb8KAa7cCGYLs4XAxkh0gGzsC/ZMRGG
g0lt3KFME/5Rb5EEe6QPxTtI6fTd+I7UW55yxzcBPrtCKm1TccnEkz/GFdYkUuO3
tYCcrLU6cOebOW6cQdUL2x4ybkIXjBMEHSGCztxOYW7uHjxJJRu6YsiWUoPt5jK/
U61b0DCkWiP7kv36aLpAFdOxAzAh5LDkwpmy+/vtOwwec0dLtP4Ablv5e9qW9MUk
9mUZk5LAhdHwzJETMsxaJ+kgtqRf90YqgYLUCrH1Kc4SyDLXUY/o1TBv/t6QBY9p
nJ73deZt7UuRs2OBmoXdEpegKoaXRIwkNvgpkzZOgRk7HWFuhJ/DfuIQh1R4yA63
yYfkYMbuSxuh02/yWpjh+z01O93LWFmHRHecq3AmLCloUTSs0W85Px8f3pxs4FRt
XhCtxH+gF+aLVQdq6ZPnplcrFklGjxtNZ050JiRzfSpg6NKG9Tw+zwavzesCFcZi
7wFGY21kj6RqxiTjdd9KKdAw6529JkPkwHy+UGec7/tTQx7x6ZUDgvTgmQCyrrq6
EsBbz2SjG0qGhyLGEsqvIXPX+o3981ch4P37SGkoynRdFnwkQCvLNe8P8MZQ3BrN
aVK0tVVJF8kZNJ/2yVgqOxVMJg9ivWyh2vF3Cu63ZsHS5AzqKHf7J8AHRMg1uNIT
euIsNTs7XL63xrjl8DwNR27ZRtpkw8N/K02tB+rDNIQXod+lF2mQoUQtnEBc1Hu2
hnV3zEm7EHFegg6vPpz6e7n8qQC5h3mOnc4EHcuKcrgzWecYYojuzgxsiQq9LYOP
`protect END_PROTECTED
