`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ilLMKPJBmY2g2DfoiI5sCnzZ8IFSgv9tpORRWXyTK8XOBeEcfDcEKW1rLRgW7UkA
pZTSxqnhGJlU+/wQ571m4Fm/IqWVds2l2nLgDTOKLoL60EggvXP/WncyAcOepL4W
bAMp894JV7NiF+Ujomyy7gNTtSojYbtiQz2AmWOcFu4gf+xT0ovT7jQ3+r7ZfmMm
lbrBnBJ+Z/DSkhtwvk9DIal1xGrd155O3QkdIKmy1LcistektNMWfbFjHuxly1kT
pN/kt9jzvqSEundl88WKZilcqb+P+vmj8RVqs4Z0cf1LnoWZiry1Uv2jtULjJw+I
11fkeOGpTa6X7flwwJTSfuN1i7k3bNkSTNvPstDfHrTtnAKXWl7uD1soL7nFtRdF
JcUSpr/We1p/l+7Bo8VjcT/0gVWMhcveJd5l6h034VOqMd38jLlMGgeHfukESkCu
230+vLxZSGZcyT2WG5h2P8n6dIAYmLC0HHulauW1S+p5m69+emR5f9337KL4gpgq
ZRG6cbjfHRzL5BcR64tFBuD0HqSmfrNiqggkcM/P2yN2bbcUWPm/fW15PXpMMztj
cwfq7FOPO0jU/wmdOBuszVnyX7HqZKrXz59azO9e3rs+QSdDSGWBxVEgBzvqa1S1
tpCKd3u+FvTmL0XDTKinP3kzQmN02DQGHmikdp7J9Ps4snIbkzF0cMhjohZCZdAW
1daScI6AslrnkilIz1zIbsPQzalFJARQp3QY8LJO+D/WnAgy4KnjCZd4d/QfzDAm
LEDf/XpEB2J9Go/3ln8fqBlbTIXmYPo7KcWpRg5RCggLtSQogwlvCgZin67cPKf8
vhiB8LianZGhFTAgw0seJREsp9P/zFg4mie+zn6R8qJedMJFRT4QuU7TazznPB+D
/pw9UZ+xSdY5fON2KgWoI4RXzF6i0xWzemshGuMXRMISvuQUD/O4qJpICSdt22Cu
SO3umYzXG/Mey1J96Nd3956TZsdzM4x2j5fpwayLdWfgR650feXenyMlhQP0Pcan
HLxc9xNGj3rSirsZqtgs1wSmdhbwxlejQVqWhRxXtpwzfJILc9YHrnN0HqQNvh1e
B93gi+LF5PQFaoBhnBfWty1J5sR2/cnjwXRFiOV6HU4BoMNJVq+DA18sjx+Oo9ku
AC7N7KcKrbkXCWt44P2TXEAZGoMDkfKql3UzltFScFFNg1cksIVeYg4DbYQh5Bm0
Io3APTuSuAiN5m6Oji1Xa/k9gQ6bhyzGIkt3PApGYn7TVTFK/UROxZkyzxXsryAD
lXOcKcdjxDUEVEuBsfe9q56Tm2j/FR6yzRmEgrDoEklmP4c7nvBL9yX5ljOqcgli
1+faVlZ0/ySpCOTkYWf0lhqTI8MHUAyficm8v/gDDif300Z1h2llIAxojFYrObyU
hZ5sTI3Cuj/Kh38vVCBjChvYbyaxiNINiqrUsikFdMVNnDjRGgFzTnqXo94C/PTr
IYePydeG6B5tKdLomHh7z2GAwNuzR/pbhOTe9ii/uVafmmDEVDx+gZJ5RJmAhGs+
hPBo9da85J0xhy6gUej41spRdnlpSisSDaG0CpN6ctnW3jN/ita+CE4Fl/SPDI7f
3y8fOWYOOGTprLoiVYefEtEgZ59kWWUDaLx/KbgLZTHdwZTW4/KJMjMuWJu9ry10
Vf2a1JzPO/jQf9AsZtigRPiTXgaFHrb99Nx15Qblwknt8K+pKKqsCEGYk52ZIAg8
4t200qh7UJr2SSTKE41LpuqTS53XwJnfc5stgp0z3+dyhi65/gy06U1CYuTRXbRQ
eUuXRHTlJGQ4nhKZqmqgWcT/NlOreniAy8HiUxkWq2KtDWpC0K5smFIUwbmLNOwa
GeKgzRSpML713z7H1hNatQs5GVMVP8ttPUGeHNaBT/Z1FwZPTlpBvzlr2KOM50DG
uVMz1lKgppk7zM4/yTLyAA==
`protect END_PROTECTED
