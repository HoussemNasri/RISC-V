`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIVZMWTrkZgC17V9mizKv/9dAeyusEaoYaNuMeaSYrq3EsEgmYUbVl2SqbLeUn0V
32RWJsIg8YqgAYkQqoGjz3MlfDWfUCg7hMMCBfo9PvSFbJw5ldZzWYfesgHEtSLL
juZ4OIwBq5FDi0DIDb0Rv2qE7ixAFuGJwIybx9Qib1BbQC8FJCfensUfynG6MrLB
q00H7aghMM65tgm/NCwPikJJJmVKqxEolZWJCqc8oGPaY6bfzGwPfzMqykTZlzSz
Ri8KmDtFPYj6pDQ96in+UUlsurx9zbA8F04uo+761cRNnGPDfyskEvbhj9wZACef
W1heS27dXXn4FqtMDUAo600eaeNTx/V5U/N0FTQavuwgur1cSs3w5yrAf7HwHi4M
bRFu8auada4DD8555WJ9D5m13zPj+cEzp5UMKOqOo5RFe8y/ndEZzn0LFVe2evt6
d4a4yG7jmLdtnV87LtZFbWsE9ME4Pxs0hFOQsu67bqTDS1FpQ21kblouf6SBgrRk
4jiRYWcNFWheXBc5o/VWSggVCBEDeUf4lSiKc3jUXK7vRYmidkNDa2oxHuH5t12K
x5uw7qYI0l2zM08S7ElH4UJ+bYMM3y191EVv3v6dlm/ACRVzvR4EBnXlP9mSIE8Q
Azk+kpxqhcOB3Cg8lMDkka3CFI/HflJnvxJ0sNmj5vK+93ZJ0wjGxhBZWnMpPS0j
xe1Kb6wn7IQmbJPCakP/l2Z4l6lD4G8hmaX+pmZsirnb90b8Zixc+4ZnxzrknFIQ
wy2fLguJg3qamIJlPDyaPDjJNunuAEI6bO1InuKzcppTlxlkLR2HZ8opwg4PZ43w
k0fFOoJMRCirKcqkkyt4imAWHeDevddlJ3zDC78gWF9JM+ahLYqUczm0WjRDyNBb
KW24/U03dOcbojRj8uURvj6i9xcyj14tP6jp6CYmEN4RahCnYF59QDJjgUsS5jT5
mLUP7aBZN8r76y6tegZIR9TwjDlnVQEZ7TafOo1d/cSaAPTS24gfqZVawIDbU9GG
rAFVCWjFRKpDltUJTeF0w+celSWdq6rsnI8ADoKMZs9fkkQ5GPyaJnSfxsjAu8Gg
h0A+eR833/rNJFs7DB3W7Bw8zAM+0Rzt4hrN4HcnzLfaLOXiHdyU8A/XGEnbP8eA
UCHrW9m/bVKCqk4o1V3mN/liq4T4zyUUELmb1RC4fnY5IaY2QsInTS91xzxyJqCI
GEHTjk/jNzu6GKcNv2q4bmhIB0Yq8dufL+vAy71rW9QSHIbi5PYZ2lcAaKD2V+lp
`protect END_PROTECTED
