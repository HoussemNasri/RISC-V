`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ngqcSMR6ebGkYCIb0cLCZdex5K8zWxNLOY4cIPnSgkYab7J68eU0TC9xE6ZBgTaX
LZbHFzugTTNkZczsdit/bthSDQWuS9Z7KgSRSOUn5pNS7L+53u8NJnqzcZheMgHP
EKaGJvfaq9cQEdRLsKITeS5vEHHPcfAg6lYcoxsLnzS03adtDpllIET9uOQ5m8Vk
u6FxC7qu+iagg7KnxI++1Sfy/1GHw/t4HhUqwRABYIsBc+kI6azNBVqnEZP491pY
yq8/Pvv/u8ERixxxBx86HoakxrS4+7zwf5l14AJv3bL3/yVJ906dSy5QA5rELK0b
MuEVSiF+bpz7fN5P0/ROlub3ch4+EY760Ce8EfZuaIBTeLSAlJqvnGqe6SDPDl7L
pFZ48vHRONkU6A4c+D+19gqslagco8N0+wUY+XcMuuAYOpPao1pt5ZXf5U9UXOsX
n2+tG0NT/++qL0s0FKrd5xzO1GENIcFZ/uVXmrleMH+RSDtNm59K3W0PrNRw9Zq3
AIIRbnDvz7ls+wx55wFjxU+nUKbFOdswMDnwYAv2xYngD5iay7HiDUMn0hCisKCc
MthVG6UfUJBpwbIYgXwmiWHE9dal+E4Dqayn0eZFY2419/KD0jBiLXOH/N4DQkyY
hDjyEBctDQdHEi9QcpTwvCqqu8qc7f8waolQkDMpBRS2G8IEjhi5vf+vTQC8Ldd3
/AukZDCZ6+qTjWme/dO6frTcy9em1fbSG0mGDfW793yt/Tjs7hgf20Y4IHsg0ZKN
KfT7/oJHXPm7XbhJiULDWp6vuw3GLeCAHuEu+ja3Hj0KLxOdGjbmysUoUyIPgftY
RiArvNdT475QZYbFTtBPMdSbDpu7j41gArrNpDG/t848KVn18jwIOeUKsEFtdze0
Mnm/jcrofkCLyQckFEZdMDD2pGo8hSg2BNmUY8KvIRMaxZ7eyN3bjTOLiSCbVI2D
kInaywnz2gFA0CxtkqlBMjIKseFFWkhHvQ15ZhRfdzKFafGDbKwSedx1stO7OE0z
A588g3m+7Ynmms4OKDMgNUifu4fhZMJeKhkeatUtRfKy2rulUbPvJvlCBc+OtW5Q
pNBFamEzt915I+gO0Xvy/c66f514230XFgYDN0LNgyFnNaJDJXufOEBywFTH4uQY
lvtE4JoslNyWRHalCeSCzGnMSxpalVGkHs6FIv2vM6+838jvGC6a7MU5PCBIZlAO
MRccScx4hrUXkM5mF2+HIbhCiUy43+icOdr6qezi8nxqxhOJUokc9HKnTXOhwqP/
Nw7mAIJ4o7lSLQEeP16bHh5it1r8/ioKmiyl62hme49kfSch0DCmS/aMeeE9b63G
vSVgQyO8BU+or5B+skjxYzxW1W/+rnDg3p353MZm494oA2mQeFb3BowJu4cOc6Uf
+Z2shSWafcuJZ0udFRAMXT3U6UffIVHSiwAalMrsZ+QeLJdsCndcE+9A4tD2yeog
OSWlMb+9B9rvFM0+eWNn5SHzqVY8EQ6mpx5gpLyY3wQjuUHxwORIkma/eUsxm9Zz
S7fVP2r05i1tQO5HA4OPt/ffeTB01iwWvEjqzL9BcqTPuul6fpiqa6MBRQq1IJK/
hXlUzN2fkOQzUh+3/W+hyqMh7RrpoMuScnn01xoG3M9372ulIXgRKD8lEaKvBaec
H1Q1B4Hs8oNrPZhi7Sci603+atIPk1rlSdlYBhBjYN202+QLqRUWyWVikqr4UuJt
qO85Rl00v6XXtg/ax+rJgpfS6I3TCVkUdN05VVey8F8HtN/egQPi2wua8Nm0lyfV
XMhcYRT5q3xQRQ6Efr4cgMpNWktFf0VWg2rowbzUWF2Zzr8qNi5QqYQOxC+oZ2Ca
gX5DCoa7xEtDUi5X0W3L6RbDNrnyrompdM0J+xfZkJS5ZYvHC8OFRzPeiLOxFlmf
azfB4PR94raZz207A1DG10IINrAWC9LDm/zmfKFuxRQfiwIFQPAI5S6DVOndQ0tS
oOpnDpB0Vfco74RHnehxL4CLJ6lJqAJo0zSxWMaf56VTkpmf2wahfVDY7Suc4tmn
JoLL0vpspbHQK7ftziUmrrZhYC3byfNogGh9I6dxbvL9MhAQsmRtJkuRkwcVcRrn
k5ZLbYiNqg6W3Vb8kg+8DRwImft/j3EB960MBhGd+U05Ql67eCWGIWdEI1mIcnrl
k95vBny0AOOdFXv+CfPZQR+hY5a5VadcXOPgvUL1nA7R78RxiHpaBBSvCLwvlY7Z
A+JvLmu2CQc0qpBen6oywLDhI7gCTiDAv4uZJ13WJAK86SdHTNy1CXGrUvsf1eTI
UMV/7v/qLACCCLdx7ZVNn+y1A+vIRzLZziHezILMU00DQrzTT3jJ0YgL2Zj9bHth
+MyrpK+G+sEao5zCemJruzQAGc4cFL38sMmR3HnNfhGAu46aS8pvbtKrsCgXvnDz
PzXc4WXviHLjgdY5qSPTqugJu2rJBLQZX/8IZ8YBoYyOU+6Uek3hPGMkMrSeXm14
VBM0/InkBE5SgRIYDfH9obpJTtVdC4PlyfylH7AW/aiHXPuGtSMzBbWr+rZuvxtj
BdbEYiLyJRbFCcqxdHC4zdbZ2U3E2P7jOFTuHyCp9qsa9GrTQl1DiQQZ+esGh+N4
VQyQ5FfGjZOFXcZ3T/Yhv0xnyQIeV+dWZ0g/FtxHmWyAk2May5QT3HGT7KJnwt62
nwQZf0auRyN4tlFxr55r19k2Tdf8b6zqHPq5h9ENo+w6CAG7KMsm9XjHlV0jRNn7
I6Zf4bm1w4xljdzUj0xI+jhxr70u8ZMQ/as5Jd1QNaOJCSupF/ZQfLLxzuUWpoqT
EktHfg0L2gCvqS2XN59g1rTs6qm9fPOy+sSWNkrMQD4k8VaUWb5F9EfRJZDSGcDv
PavvuvIpr7I62xSQdxBLID3IR2x3XEiYvJgKmcAOZVK7kdi/7ONUzwIz8gZ0E3jQ
DBEnOOOy9O/vPbx0xu7OpESWxnrT44gddqNlZrCFjNjHLkqsOLs6OxhubWqGSIyR
lIaZfSGmaqcYmvCrp1y9pAAF4F/Z39+e1Tu3rTbJPP5D6405Q6POkInguFlVUmt+
2juk2NxMO8uscmH2+9Xz/pWRrDRmssEczynkli8GRB1C0JKCKa+zmSiXe9e3SsZm
kbEB/rBmxjagAKErzkAXj1/C7ZPhhzMzfl3YmYyk8Sq4N97h5BqmzpSAIc9p/bA6
ywm0geUbdQMqNdhwYqtPZEPTzNoApGcnpWub5JK5TQed+LH0Dx5CiVh2Eqf2rx6n
jL5BZFLVJlk1o4lq81e/lvgvrERVoaE4jfsmxw9BBB8j/yuGXULJuxcxAp9Ff2ug
YAWKUgoSScEkHt3jSRlWu8tKCUTE1EmvEOscgCdWGjFveWAtMilmhLqfLsiXylt+
1LSjkPi/WRxitoYuJoOzO3DdNYJ0+LDlVU0B5Z4wOZ9ZKPiaMxi8pWhsPXsxFd5r
Uj6SUrUd62NgdPNAzodSiayD6W1l3e+72HXgXXlnsMWi+zu4yp18Uv9SDVPzsn9X
V9g+Wxc/JSMjjHbltpSlhZzqUnVUKrLKrIuMHTL0uZW3X7xCr1e4J9+z8nMcordj
w5xmqNarchF/QheTu0p1mQvI8dviHBdQeJTTrJS4j+FA0CfiekAshXfZ1gupRnae
JPEBrrkFHpyfAm3oVY3KIJm/A4YjSfGTYbCevoU7pZX0pFLyjaDFw6ZxtFqNgFcn
DFlCjG6SKu8PgBrcvXffn8eW6culTF8MrvedS2TpVlrK1yfTzQlw4LRmqYhF2oKd
cGPb3dreTBfaiN3rq6F13IH7EkWcMfK4I0Efg5KBCwPHmijmlwP6/Vw39rsvZvCC
4lPMMEqpJcBYW6V5AK3Yoy31KP35K3GsbM0ZQkZb+Gbx8NQLR2QsXFdQhgAeCGVy
JXOA4aod0iIiPz333Zp//s+bVm356/R7Bn1YsdwJrMGFFlExk9K/WOTwysaRToqf
Y6A5G/1qIYD84spx5La1uadfn2DBX8+hsJt3PBL5EoEk/dG866IMNHdvk+1Yih2Q
zgKPb2AXZFRmALlhTV5rOIxPgPSRfGDpyDuxLSeh3n8CC1MBqRz0UEi8sP7nMcZY
6p6Qe8UKAABK2VOMXNyTHOG3Ixkax1YQxjIFeQYrI4NFfzbdoPFuHNJGnJnAaBmZ
q0vHj9VvOZgN5ihcs+AqTAi4ng7S61KbGFvYNj5nd3LOElN151lT2c2rCWj6ZyOn
ilYxwqeq7acN+Wm4TRoc4kgaPu6YJ7fUHRZ44uCvNev8EfJRAK0aK9pUbTkCaNUq
MKZVi+NKcpRwamTpU0+yrBm0rzTzjrxEyXbVDZn7x4UiyBtXR1v6wZITxJTVVLNF
8oaAr6l0y7Q010HB2+YIgfQQvWmAxPX/saFXxw2i+wXbBwug3zmqnJ92H2AdGT+o
P0fu/mjs8waknpYEDwiMhR7luSAj/K7rhnMZ+5MWh13C/oZ+vNH4t5ryU18ax1HK
R2CrfVlKBE8LLMg5n2DSVEpkv0nbOgRRusNTJDCN+9QXuJagCwvTjpR0yRz12phr
hOeLfdgrI5EmONBCUP5oUSjRwC5qZ+x360tCitl1CrgAt8GnreJsp83ESHH08/jM
Wx98JSifnv+p4jJj0uGwb/Sy5AUViM9kdmG9cXH5JVFrGw/94OuK65Kf1mdXVM/W
5NO30pCEunqsdOZLAHpPQneBufhcfTGc6Fs/0BE+pzg74mLzWOHsETYBO0BeuiBo
g8tWvDUEll1qvUg8Vsb0lDFRYunIi55RMesLBQjwnqkEk5bR3IUBtwmNt+J04PlR
79oR908fuYOnfooP7kdmLkieaZLM4f9crnIdcaijOmga8ZDl9BMHI4QAP9rqyEv/
94zRPn9miywzfBmQ7bD/hggt/L0YLkraa3JKlXdBFKHXnPyjwnS1KXMZMwRCk0FE
7OPzpPNo9grJQPPtVgNcG+RXlMTxmKn30zGVJ0xD/FmtPYdI5qW1LgftQiBa6S+L
lbFMmxdn/4zIkH/8ZiPIh6IcfKWBgpwhu89q5TtXngxZkclqYKHJiFzgCVcEo2gc
2t5l9bLyvYtNFCnjE6WjkngJXSDxXHMC+w9dsYyJoMavpmICs+d8inJU4awZlRYY
vGG0f+332Z+3V1/wYVHvZaAyyqMKOK5gUR4qnU6DUAo+KclEGGzcL4rm2vgdIN5y
hgfOfh0zSyeC/zqCy7KRBMk+NwMDLpuaUAZSxklBTOiB0eI8j8SvMql0tMkTX2Bi
GfPiE7+WQ9B+qui2uVyqZuo8+X9SgP2uUiUCDWvqhvxSuVBaz2fX2+C0EqUq4v7P
pLfV90Bgy9LaujgFrFXneO+7TaLYBjGekGWXUPVT4N5Zj2fClO7xJPAW7Je/kSFS
9Ys/ctY6UrildSNuwqpQb1OAZDfnEyKG9rAKmaAzGdJSHZhZOgmzjlSjQtk3peW7
A5ZOEesOufLde800UFgsaKviKw7k4oYopFYbf4QJTJjRX99iCbkTD/GqnrzWpd1L
T6vS7O+rbIdBFJRKWHtTrWTigVaD3Rh4BTgyLAJ2AvdiyvQ2WpHUfyn7Cx/xvMhL
obQ8Zn6NhkWS83tl/efGnZANd3/DzdiUX3SpEGOfyhoO8CVjKfjiP47S2Kc4oCLi
olAVRueVvAwaBlmcBPD9S3J0E5Hj4dYyNZse2+4Su2UVbH0HOwi2+HkMhgL1n8ML
FuPnF+TWjlJJTW7jq3jp0zdyTmFx7lCiMU6fTGvYSICqAw6jFXX/U1xM0xAb7k01
gVs441/H5sJoN0XQ8aGTP4DYi3DB0vAJHtDE2BaeyB3Q788B/Pli+NPkApdS7g6V
po8nMiaHjh9Li+myUTbyaoKDdxsuK3/Oed0kvlWkEJXQj62ozTRUPyX0J+o4vAMJ
Z3rfZvBwY6kkGIRQ8H0/rpRvU41RJ5cEh0CNyJ7mcyf+EzvtLi0cEvPY8JiBEXf4
7HUFD9S29rPVBg4aqwrcBkBU9BVdS90u+uk56EIOAezC+wAH86a9HgHzkFQKJS5N
c/09NXeZGB8bgdvSgpsrlCRkofWDqaplFePppQ3ZAWmxaYgjHnsDy1sGwiIR9xFk
GaYuQrMKO5J4l/E+u+zJv5ZJRNQo9l8pQ5G+A/dS5hyiaXigJ9uu9s3AAJxUSoLZ
QU8N1wNqBybvvKsej1ZZAG4IE6dr/nVQCS337Vc/2Yp7lUBG9hCMIyN6Juvy9CO3
eFUbUTEe5Jz7oPGLy0Ip+kElRMxsAukMzbbv1P9f71msUfANOv2EvNT9SgMAfp+h
SW8O9I8z+rsDyk130wCaRCki2gG5ddDSm+EXdL/3T2w7YHE79/vvvR41NnGfaqx+
QN9bIPRCB+ae+K4ehWSW4XnC/SIAael1ZJFCec1ifvAQtCX4ozkkUqmYmSg2MBDG
58vuYh0T1m1s0EZQ0zOmz9wcwSO0fjCOiO46ICr7MFvLhI4lHVViqNgTZ/UiudgJ
mI7ugi//dFi9csb1G8kGzXe4ZiWE2nxzyMu3O+3/CxvyfB6MgGpD4K42FjM6hHmZ
d+f91O89aj4kAqivNRPwGCUBjPr/9d8d+1DdjhHAgdUJMWrncoFZEiwGysSEq4Mb
NmzvXy2FBOAoZd9r+CbRUM/r5bp/ll9FT/BqzZSWDWC1AV3CHzYgNPWVyFgVStwC
+PZ3QvhYaUD7OYMEWYc8OsF6o5YMTZ6uG5K6NZhc0AFryiXYRoyBwiopMSlMLN8P
9pwQOAMSXvxqERxUNCEAt3Xgyvyrb/so/1K3mdEUIfVSkPawXKLGMKE0W2y1gbHc
/FtUa160Z3qTfrRLBfChPQRl2B8y56/KwNCreZAc3AoVF6e4ez+lLSyvicHoPB85
79EhYjkzVKs4icvofpxcPB0wldWewZsEzG0EDPnC+K88ArfIZQOk/gOnZQd32/bZ
+Xvi5+/Cknng9EV5ztfVUbBARDX/R79L4A0TiAiUmy5QoL7orbYt08uA369Qp9ou
6OP46Y83thEuwjxT6fI/TALSxBCRgfSOGLAmD5Aq6r91ANTBfaHhpiyWIFjIto6r
xAoSEX3y/56Xh0aQ2tpFCRW8twahm69AnhYHBAeJ2y5eD/Rki+WewfOShh8dpWcB
BozYULWSUyntyAG7S6B0KopWBk5tGSnnMYi78WZSCbkwlkFLZYx3G1FQfnO1+CU2
lWQBvWk686VPYA2roUa8p6x/OmlcgSeM0EaI56HjWufi0M7M7W7t/137RY2FPvde
bw01LY8ADEvBprkVnnLLACAPam6fG2cBlI5qls5YtNmdyTsZHuPxV98lB9VwUJsW
tlv2pKS8W9USKbaF4hVJkw==
`protect END_PROTECTED
