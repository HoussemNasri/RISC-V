`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lnzja9v+l/M3Fza1zl0p3aY2SZUD9cesqxVR1qDgXlMMc9na8/RNwxICTOr7TVtH
Y00VMEMuupBX7wgne0qEc2XbNIFS7xZWfUzTCCGYoiS0zoGlkJJ7R4izdg86GCWo
hlOzLVtF+thNkGZTePjq+fN3FUKtj10HXJTjtrrDe/eutM4R4r3vzu5/2dusxPFp
ba1Mxk4bN8yDH0XPOu0XPeI47kwKbGGoJnaC0D73wGl61NJt8ec+7RkKOW8F/egZ
be65R7+bPo1eEf4S2/xTtpmQd7FzbgKcM12thNH9MOcu42wP6HbSla6B4CArrko1
Lwilgf+4KrS+tBUXRrv3OsRL72OlduiNQtTrUewTPtGNDK9QAe9eD6REN9YDKVvX
UXcxqOCaTvkUDADeVbT0DcK43z362+aOV4EOBQV+cOBs8G/UZJQRK6dTBx7AVpTX
tnjZaVlPCf1y/Ko8n4V+oBIUjdzwQJL7O4vTIZPECS94/mibLjDPi3WZanKrFGF8
616oOduTtMEh9tiXlXnSkT4xkBvp7oGYEu1udUsVpej/g6mWw0ohIK/lb7RLnHBk
ETRJURT/m1V9EnjL6VDY1Jy2uOr68SWw734/5/QFKRuqwMJOZMgM3PYcxlOoazKB
OHyU1R3tkQ8PDpvAGu6uzyWFgbGnVCLfTMr+3nJI64QunR2W0aeflHbjq/yurEqW
Ul9YmvZ8JpOYI5cYlhNXDUW+m/lGMcVsg6shfZG0END8wpeKLBM8ooQOqpfExcZH
969+RPznEy4L8xkmCqS9ciP7zUR4tnk5PU9nROp0q9icjqMZaL9ONWhk+zU/3VpJ
bQ/Rv/qnPN1Ot9zaPpk60vJ2qwIl3WD2kaa5yH3uSagljukRe7NW9ePfNU/iCT4F
NNrzzlGTqyV8o0ygE5/x+xGnEtp6k4m9zN/l8iSHPazLW+Vu5sOoKgoQ7R1jx52F
K9+dQyrR+LzRd4KtBKqCg34zR2sfyY9RJLB4KpIO6xH9G2Jnnv93AZZxC1+vPefW
PLl6tWJrOjUhBiH22Surs/X4K26c4+SFe//CKleGqAnUyhTkCqm/OGaa2s0zC8tI
pxftPc8oWYt7TtyF0WIzzc6vBt0fvsZSwms/nv1MzElGXRile3J8GyPwoRmg3afT
va1y2GEyFYQ5TIsCSzP/gWaxOqFKWQTCz7Tsn+2i0EC+GTG38CoTTg98NWWnTn7f
9b2FZvYsSJpLV+iIuWuOVwj7ck8Tk7P+rE8W+VtShq6Rf40BK9OOZdE3vsili18j
vC2xFf8YZNrZ/088kTgU86Y/ysxnav78vfK9ZwlXbAAScF9ezhZW2CitcAQQu9pz
dggXKapuxnwRs5MSFTzY8pgI9C9U1J3TyZyjelaZTN20/ecuYSW3ta+gbejq6Sq3
dJ42TENx6MhTwCupoIFijsNJ0kC/cJuUvjZGbx2wLUE3a6ARKOZFgeVUAJ4z6GQm
lIZ8NvC1X7hoQpsebmSECvbqBEHNijY9DOQrdF0hnL3e5gP9vD5FZJ6sYG4YX9fc
FVdNHFhlNhVCl5mpTaRyrQCrNVjC30YmpU+KqAf6HTF26cdc4bKiqIJ/Mrg5eWhc
5KMvqapBFeyf8V2alJZPs/XMQS8VGR2CTgS+ivyxoLvlKSYcUZyOnwdDiEUmnuHW
CKKVPSi3CO7wwLOHEZl+mAfC0EhZvEKf0xaCscxoOFqMwf/+PvEZ+vWahE6IG+OP
ammdtgk5PFZTPcpdq8G8DPCK/C8br38tsmrGd811rAGlcL1zZtEV4iXu68YNx+Io
3HiDIywsoCDcWJcVLooVY0IaovCWbepFHrzeA27cgkM43vUv3U7GNO6T7WwAZJS9
QqXyHOyyuBDwVODEBVO0sIjUT0TzIeCcOg//+/TJ6adxbfqDJ6Bt63NPa1P/6d4R
ca7lOry1meoAj4o5xkq9/eDHBZMoT/7560NOMR6AOBxdsg6OrfMrYWkYtvN2zk4D
HyIqV2FfLbqkqoDeChIJwQKtOXDTBQp8SnbFV4idwxAGLDlMH5uU7ANV/oXAx2sG
+Hq/uiELg9h3IwMRmr7V9ra04TtoBTyPJTIXH6zIPBRrRYuf9kH+GR7iQPdgHV93
x460GMSB3gGvDqKUbE5DhfLPjiGWVtOb+PCvcKmuxJED2WSS8rwKm7mtT15NtYb1
ouR0AlQRZL5vHVccapo2BsthEhCpGBGM7EpzAzlFbpnRGJl860Vl3XtnmW2tcjjU
U6BcjRRIpuivO6pKhgzLbSygsewAMgLM9dWWbnXWRSH5FuRfjFOJ1UUN6kjitbwI
LBj8eABy2e+L81tAMTj+aWmfVRK3+GERXJTXQ/qJzeEdGuGlbczTEBWyjvnggexe
PSb7A2yPG+KWSp+6+8fdXiuGcSRZ03o+vl28872i6GIuD02rIaBlZc6lcOPcgSUQ
XNbRQhQ2ADvRfFXhYvpmt0xtZXLcZbnprd+SaBJNj5+OGtir1iZPHwpPo/pI65Q+
uLGmJkSeTaF9IbgZ3YAbjIqV1f6dv96keT9cr0e7gWnGp/QuVUQQR2IHQqUvObE0
zklU5+tNtX8MA0K63p6hOIFH8LAvkaCsctt4wmSvFuDKYGOktouw9AzpwBxUfceZ
/laTV8Joh087gWXvjQnfdHliB+rZQBL4KnFCnQ8TwhuCJF2utE0iFJAzvYb+hQC5
PWzLGFZs5stdxGGJMa8HNkoHKys85Zf4Kvr82AxrYZxmEsonAiiGGkv2l5Sq+9l4
cuJAoSRYLYFUEzUvl4C9ucNzGO3rnPKn8/CY8RbUVOFxIYYsHVSNh+xO7/ST+D0X
MstLZ7Q0j+beg6b+5cVzJVoxqTlG/C5ThaO09BHXjCYDyyn0MXYvO9Iy9jElcMbK
gjEFmW+EAYSA/baKYXvJe6wphEaAxyMqWBblKLMUFGiVfUSg+OrSv4UjYRS870Rt
xyFuQByxfutkXpCEy0Fp2DU5l1cpUjE7uNb0142aGlPHDj9N+C0iN0KogxpMbSKl
DWceSAjHuwTAmilKwtNHxNyj8JwxX+5MoMDYmQ8WG4wzwGOCAlah5iDVMyyDCTOQ
KkkPjlN1nP/MpTWLpDFeq3lQZMVRoa44DgUDwPT4iX/JaapBXuFcESV0YR+Fount
W0V1fYYRD3PFWdDXSz0aiR1qBK/A5wQY/veXXCbOaBIdBKxJQ8c/ADmuzgBKhAhE
Ojh1V8GltdU+auCWoUGmaNFpTVUBp24DPNirKLWhJ17wkCG+oU7uNw6mK1lZxduN
BzBpnkjnmp4ZsO+VUVw1QtrVTsahlbrgp0ZG2qytydA360TMZ+j1s8CiF2bXBJnI
C1fv4taI3Euug5s/lwrVHKFY9ED7KbdncX+nZ/6EeR1TtowQJF0rC8hHI/BReOiF
ovzjW/qf3nTf/j3Jqt8rksygJAiGh8VOi45g31070l15Qy/rjUkyuLCwA56o6xOA
aEt7Cz+D2B7DIT0hcvXeoU5Uu3cWYcM9AmD7hCljnZ1wHK54i5V86AfCD+HxHoCD
i6eI2owX/psSNsvnVmLchNE36/XKmZBYs4feR/SGclotsCnxsPk2bjCTboJle2Gj
2ZyjjhwYHwo/RGT1vu9mzZRBfcqKdYqAXdYbYVdsG0m1kdi1pf/4u9t/HrWP+o1j
8jJV9MDEWgw34HofDZ9d2SZSrpC9t9S5izNw4ylq8iYzsyI6K52y5MAUOWD6dLaG
eYpHY7j13v6lBGjybZhxSt3gozt4vK97Ee1EBJlWvuKlFZhMt4RgzG0NkmJNHC2b
e37YtjZ2YbFq/SXgjDvyoGFyU1m0a+A0YM8d33Q9EZ/tyoCjTyNIlYADD6Ti/a+2
BJg5UlWpdEL2Xo4URWGWv8aXc8Q/f9BB4Zy6pvvxNy/5EhfL89CGl8tni2HKr6HJ
aJaCpPBhONqQVqibALQ9qYM9fPiTeDjv22Pv2A66jeHCIe43YegWLb6qIWSUiUgk
eHeCNt5Kc8Gkx8++rgB6SG/UJ8D9tor4zscxO9VIzcryJfMFX5ROQvUkVzw7b8+9
4CeqlC/Dwjurxsb/29L0t9fQz09S9Fwfaxxy222Z8Bs5xgb8PqpZQ0BqPxv/175l
3IFwmT44h8T3gNdrZHBsp+Rm6D/BKnryDYJc3KuB6tZ9Wz5eknLAcpttKsA3vdz2
Oh4PoSaCA5yuJ6demJ15/h/YOhApowogIY1wnuWFNBQEcj42UeQX6OJz02kSKNTX
FG5ryFxxv3l2653hIQt5ELrRM6/piYmE86JUC9savKDr7y5S8hUr02xwXrCmTl5I
RX7wdJYR8Um9p6FKMWg1aP9OUEJW3t4irnw5WlcyGsX4O2WR8Pt+3RBqaYXbMIqd
2amadzDG2Br+FxmJM9lyXcOnNVKhaLr61P+s0aiNDNtUg07H/EKWT6UVQKWMMMC6
2aUSO4KIhYKULoYenP4hlW65Mbl/ANJsj+lQSRcFs5HNwxx9x6fRoHMLO6t5uTdO
f0iNbS/xkLblyltb2GjXRVht9LBTZ2s2Lj4X+8ft0d/0APc17qo34HJ7h2kHJbdl
0FupqOcVrb8oDJVLaMG6K6FZ3tY9xRs9VI0PLkd8YHZKVP7GgmsGOWbp4D1j3QxP
p8k947SprOnHsgogdiazWzcUqLujIBQdPwltWw+UkdgyiwE4IBWLXRgN9BSBE9pw
lg8WTZGIuNVXo3+NbtZWeHp59rehPFYrQR2nUxVocA8C2DtKH66RzeKmbxu1t67k
R5JxtLr/L1g67x8r6mxRSgY9aA1H9G1LOK9MBrWiRdgSn+UCSsNVQsOxeVLEYPiF
k86E9Hw16wTObqP5CCvDngLXUPyaeu34VdzmI/OxppzQvcV2n2OVX994IRozt0uh
772zSnbEvqrHN/Wkf34LbUb3RKnxaYo0dvB014waHSx6KH4v5G6mBC3us2FLkJiR
bYRdXVdXusKZ9q38cfhgMZShdW2eZMeOzZlmBpqRotKjjTz7ulNulZU1ZVGA4kRT
VmsJUX5O4SYOW0R8vfs7Z6wFpPbu3QLpxa3ScoKDao4S9DGFeKW8V6lKdnwG9XTj
TEpvZpOG+48L+aIDW9CxFNbnEV/clBbjv4PQgd3Kv2IEuynbG8sMWptwV63SDHNm
JlcE5YNfOviqR0EU4ZWuWuPCOyuofeTbhW++x4ov7wA9Abp1F8mHR9DxnlHY13WC
639ScK9d7dsOm2x8QbVJMV3Duk2sPW9xsKmKUTMwgfdVEF1ES8b5Z6p2lb9dQi50
bwSmGf/sEeIss4M4YvsmP3FZf28TW/uFFGitdafWGn83ZPWpK3EPHCYre7OOERv2
340htcU9sBhK73shFeJLPodVUrgwEotlwvACYvAO4LoGgle/wLna6tia0YhhoRel
2puhdYgO8KI0XwgYfXIejm3Y0iIl0i9tmRtEqev6Cp5Teh4Z1sJq8If4kZdkVKhH
0AN8K+mxeDNTyQwX+AQpUoTknqxUg4J6vLGCMIsIbnqbCZ/rExFotq+qwAhz02wI
ZUWSX3ny4BDT8+NIQAwETfWoCh+Qbe9MJUvjAn5YpeOomM/BPffziQDclTqIT0UL
IV0qvQroa85xA3iZ/y+DEaIEGrqUJlHXR9x9Vt296v+hEPrB6CjJcB+uDVROShnf
O4LGKGU8Ga42c20Feo30XQ==
`protect END_PROTECTED
