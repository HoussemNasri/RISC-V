`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dC2KT9+d3yxzLIc3P92uhf6oCyPJImEdp/yE5TQ5L3v2ATuR1p164z+pxQsdo3cN
VBKZMbABmPIQxd9zhAaGzQe6mWQ/OesxC/StrFDOPY6lseqQaoRUFp87lS7KyrZZ
08fCtb2I7ZdHD4BWbm6esTug3bJwEcioxuBRT3U58EgeOAaon1fs93HrBp97r/3x
iml5ViH7g8miaI/P6a0XlOBoafMVw1ThBZSb6J9mjtARwitzbQfwQTYKvWiS24MP
FBdUb5oqRtx1MvIsq3HFSPoMZrsjlv1uIm/wOeP4uzxUSvlZMEtTihjhDezBT75W
DD+5Xp2uvl/xPyfQJ2gcWfBPAtNkdW5VRBiiXEXK9ZQAJnvRB151LtE6mJrpgUL2
0rmurvQNljW4j9RlMZA4Gly9+Vx7HO+k0Rt484hi+rRKSTGDV7nQ0MnZiYQnQAkO
uf7AElNegs2Xn/su1d0LII9iVf+Ch6AYk9WUy7RzqczqPSa4GX2LGSRpRDGNApNB
ZMLdSQMjUu5cst9pNOhQzynY5xnYk8iqohTyUg+qsEm1QWMAMb0/pzIl9GKk2GDv
mRDdPfz+NqLnifHxqGHi4XTFRzga9NBc4hb4Xzvn7vP6MvuDTF4TsQAx32PK2n41
ZUCURRlVn1uauIi3Y8YwinqLyJLmZQWlgBPV1OEsq9OQp0Tn7jvzP0fWmzfpvs+C
0qUCu83kv9sxN1GgJwnza/02ZO3W6owTmg3t6SG26Bi34zC6a0NVEKz15J4h14Fq
zpz+3qI3OdEZIK0ji/o/lExsOPfTiEmMZwb1SbNRe7JTEaDPDy0fb4LmQy4iZHC4
VnXtD+NF6DRKydhcQ/J8nofjtfGuJo2D7v8Z/ERzAQ/82XT2SuGtATmxLh79yRuR
JcTOpyvd24s0D9fzvOcHBZ55cdHbbXQeQyRDr2YBx8AxAAgNxQUP+MCS/5eHPfLM
tKNbMwxfy62if4QY3uNZ+7BTKj+oFIeqiWeb6tm0a0we9ZcEKJfI3dLBD0GEfj2r
myAbH46jhtr3PjMk1Oc9ADllTfUT/fyyaN/yIst2exf90s5AatWSAD5FoidyWv4b
96ul2IV0gocuT8H37B5FGhd6Hw+Eg7smSQJsGjzJFHoAr9Y6MHJgwMbyj/cgVCKl
08sHC8T5giaaZ9wuuiFnII6ypRImGhlX87FDfT8bdAAiGWM4qf/g0BoEkW3jnagW
2WHNEjbGfDTw9TjBEN9xYDJD7Nxa3vqztSlEhlesZqzyMieRngJLv8WQ6caOjwEa
KkqP/XyRvnqEaf444ErsKllUpmwYtT3r2EdMxpTv71L2dcYGeA/EoiczWScel3Xk
qDztbqkFlk5bdCb+nf4nLOgn2PH+AN181yVQzU2UY3m3o+4ehGdLbm/k1OdYzuRt
sDqtOZxgeEp2KfWcVI4djeL5EwKdM6soKU+RzDdGjG+61I2fZzrrQgBA4q1rX+no
ygNH8IJPRZm1uYjelzZ55SNhfquznabzT4fcOCIeH5HIIAgs53vqIDGJL7K6bkji
sVoVujcVlT2NiPcYntKCxm3CHWlH1CGoeg1llyDfsRZ2vdxP01w8sZTA4G/Z7K95
qqbbw/ZOBaTttfx1aaZODLrut1YQOdJGIrq/+pxIxU2ZGePgsCTJ7ORiB+VyRC80
hkyhcsmWXBZ/atFv8ouiqVGtKHcP8hAlB3ak4Qlo7MyKYwQtHev8DuyJtunFEVv1
c7RzW7NAf5cLw/fGDGgb8iRK5qkqiy2z2fxf2IcOjfusnRzvjuOhrUq8vMByWKfU
`protect END_PROTECTED
