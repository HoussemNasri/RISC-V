`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lgNQBkqgPwh8DQRhG+mgSrvganuJLym+NhEXtX5jPQw9E/YFkYdgQAu/ZPHyD6iT
sDGDGYzcBofSZbc/p23u6xc2bn4bbGiMWdDkyeZMEn6v2BLXVjbohPBi78sbhJQ+
sy4NcCXZhS6N58KgAryNI0HFh3F4BscXx3oRYtx/6LQEQqMV0IfYyXhzMge7I6b0
cdv0gRjrd9fQ2IsN991DxqXjIiox8NUOtkuNpLi1V8HSpnXn4F+CFd72J6i/v4oX
GeKpWflYzSsW6/OoXhOqwIWYhZ5enxG54RFevuSGOlkYm4QAcr9Mutk0/uWKkZQ/
gpWhXLrk75JZPkenYHj/snmEscykgkORXR80kJy0wavailhHZaf2bginwDTddkjK
2EwducPcr8FWAMtGPuuApUBdML6cIsoswUjKfSW5Du8r61JwSv99Ny22vNTmMlrO
+nYGuGRfETDGxI9sStD4E2jfIJkte2iYV/wU4LoRy9E7D9I0KCl8sY5e0I1BP9Z5
R2gMuZ0IQVS3LCPNG72OJ7CG4RCZa8SVu6NCKmQqF4EaLowl68BkNYizhuV3Xmzi
WRYYsAKyuMrYzk6IAav8nZhEohhe8b7gpUSof4qktSiEEvSk1PIJgoLzmCD6/W9n
mi51mYZ2XPgai+eRSTW5+Bk/9QxKZNknZ2kpjhywfmvvpNd0MQ+h2tTBOw9MothP
GJBrOKe3qp/jTHZmQN21VPCsg40Lh8zniok0oSUZiX3t5ilfTxER++xG8p3SaduP
xblP913bXm0f5Rrq/+seuxijPRA1pSLAkSFH4L7k3DGoA1EnpNbGGbgNY19vl5y7
xAOT1fGxbZFu/fQMY7hizpAcjJzHbF/E6dvty7OtnRaXKNM3li2S5UqWoCCmyEGC
CD2VpPMtSU2V4ZA52dX6o1jSkonm1F81qTqyWI5AiDbqeiBwDei/ZaVJuSDpA+YE
a0kBYrsxmTdmJqHU2r57gMUlsiYg93FtZ/bmkF0z2e782RP+EXiyd/9nZRULjTdZ
/H/6g9lndmSNzleNhhMQ1PGG9A32Pkr63vP0ZhQoQuRjTO2d0ytXCWa1iDQhmzj+
I4Ef9IUm/vozX37J5HwtnXfKYtoNMBLJPKR5YOzgKBbS54rjYFKgT67ToBlekBgM
jT5pfyhoZzaNMAsDnCEIpTLGl9+QTXqbyPAISIcZJc21etxq2F279Qi6xq5t6vlV
7kY9XZtunAJowfy8q4Ss4oAZXSWk0IHr0vjVmwKo6DgMBicr3/k4x6RWWAYhVMXN
T0HnOSGQFd6/TnhxeFwa8pnlKM27x/bYroAZ7tTkGmdi5srV+nyHBg3BJeGaZvd0
K2v3VKQLfFGk4x2t4mzqTVjnJ4V4T91ZUg2/I/R58VXpyRtoMDqtZpiflDLs7ZtE
tUkUvQ82oO71u5ee+wJku94Bms3DlEzeXpp+G4ntu+HLnVa9WQkL4W5/58pyeUyP
/HPWypd1T93bqXndrcISO6/Urbhsd7DxoKZ9vrhPKe/aO8wZxHoHpkVXYJn/7Pe9
4wBoVdXTkewhXRMegNMA2mTikzLrzA45sEA3j6oTeHJ0YVtzzfj5fkuUCUDocZf4
VCM8fKrNqL5aQwKquwsGvh5Z35SRm/JzRsCaJeFhFZ54exYu3/zzX75sRlQka8ie
93fIFTmFgkRpwH05gVI6t56sUOaPkxfWuIQjmK84vqi46XAfC5Y8+QHs5+Cb/lIB
vt06pUT5P9QdqSkk2vJFozlqQy7s7/VphQoCwWWez3PgZ/IYXYnZ2Y84ka3AnFjl
35R+roQYM8HG2cfUJaia4IrXub59VVy2zjC6gJVdFieTGIVj8JKUwoUbnZUWoBvw
oxPPSiZIEjqnV5Mt6uH+8w1L9X9jcaIyIHDsJU3RSOoz423AdUxq8WHUxadNblmN
OMy5nzxXtr7kBLFNqBLwOOw+e7yspzPJTbQW+m/wUk6FHcXtfPBnDiBMc4/WSU18
NMlPR6JANtH2tmkfGgLVRMS6fMa7gTtyJ3H4IIc+dAQW0qGHYeyRXJDgva7wK7jw
y2Cs2J+0Wbc3Yg3iI9ucAxErWhT1XKteXnaHqxqFN8VpcSNr/txPY8VpMfsUQ0y0
XFGxPx1vDWOdd76ZCzOu5vB7CUQr2r4HriCD7SwxJnPPChqI6gPgCnz98KqstpTb
fImM1UVqWC0RZzu0O2rO/9U3poevxt9mMIfJ+MdnqKeSOMwqchHQJo9FTzt0H8hz
FuZ6aj0md4HT2cy6tU92kFWt1dqoUEYOndIq4hGTQplC7O5hb67fqoHXoIt9U4+e
qtHqif3CTHlKL2KWdzJ0PybufmwDJPoyqEVg4LTcwryPwAi21o4mPBAYBmOyov9v
ZQTWE5PDCRsbevTTF7W8TsBTnlPSQ7G6DyFOMorRXtSd3cWKuXXdTmK2JaL6Pa2C
615fr8uzp+Lo0rknDHcAxLQiH0jsc1VCfSrfatXIRnnfETs31kh1VSDYGIFJHdz6
vAE0qoXPTraHqHJU0UWwoT/CI29JL2VRWMelZb1VQjtvWcAstdGso8gMdo6LZBcr
ZYFikAHyVN5tUOhq73IgnoxQqWCWSmrlAP+eyhR+5tYIky3DEJs97+d0P7vlJdso
8eu3iDYguJ1N9A3jbPiPSqwDrwJ14r2MUt5eA62zxZT5/t8R9J6lL8UynVXvMrpV
vsnGCYBktj99jZ33Lz9w4CBvccWu1v0232ahdNziLFWqIJPDBKBud5Ts3Ybbr3XU
kOnJYjfaTofqZ5Ncz/pTOoaG4VKd0/3m9MN1FGRh+u3YgjUqKVt8VdHDtofA6So3
aHKOd8iKn3lYgtDDCCKbsD+MVfk2z0PCxcEanVjfbXsuXHMAo5qiv/nF22bnRmOK
KjcX0oqC71R1Ok0yXqdwnkSL2DnCqtO8+CPe8ROidmOHgMlPqT/+y2i7a9r3VzxK
7/Ke+b65xm2CG9urNftxiR3lQmDci4AFz1+KnuAYEivAx1RDByieWjoRiBc5xhNn
HW2JH+8zwmuvNMVqkwUR8AC+komhx7zOlA7AprRpEHIUVQMj1zfSPPCyWUjdRJlC
iUHiSrIf06LxgUEc6GxanNTfESPIbkpLlNSiAAL56tamZuqRPVtcc8medpicklJP
Uji70zRpjcMrQAk0+LCAktHQG7iIBrzZofFO2oIDtWyAmhiXdFS+ipyx1jBQZvGt
oo3R33k3HX+75WceZvm5YW8jrk8G5+vhw47kKQqaKx8JBTrGV6UoaeIk36M7qYPh
y7wWhXfjHQf+8MnxeeuXAAZFCwfGia7KUteinTqeqrWUEXsdZe+Hryfxu4wdyR8W
hBVkwppRtDYVdTx7lS4vpFQFnueK2MZoVJ0pB4MIqUWYqsMSn+XX/HtR11rrq/Qt
90TUC7LvP5cpTGTOHmhJ+L6Bcr1oC/Pr/GHrSw2EwAFx25r4KZpzDCD1e6EH1Ez0
7OCakBTceFLo2o66CW/+MafEQmv3Nn4EDlULSLrLUPOy9LDvhBJeC3rFYSU2fY4d
KZPG40lY6RrfgpcyK5LaLaNj9/Z5CA5Aa/I5yLlgM3+xnWIr3KuRKdupQvWbmMgX
dTv4nPrf7juqygRmkcu03I99tCM3qfUTycj8kgFGg0Q3PJVkjB58pPhZ12S96JmD
21RkieSVb4P6bWR1A/jXZ6rdQg96MGEnY1WC97QvxbA/zzFuO0hvBLQKqg4CE/ss
GsPLcNETjrgMJ1MRfKydsZnzcW2nIeERbuEooDnQ+VBaHlqbaaXVNOb+UEOEAq3/
rvr/PSUTLH2ja3M1ttkXSgTYPv6peBlIq+IMYtNqxriJfTWLopMT1L85qjJcsXu3
28ioosYys36ltbP2n8qXYZWuQOR6s+/jtP664k4nS8u7C5A42hLhPfDFE3dqVA9m
3MzC96mHsAh+VkyT5d3uvErngf4EItPSLEFRivolZUp8t7on1By3BNjnzn2NBmx4
Bw102M8V9TY3DKpbpUK2r4QEy5HQROIRuyLbt1xDlQktlstNJYSf4jcaG4fINrq7
F65w/seI0VDx5XZipwNEbG9bP7WWppFUQn2riwklBAedBhAUmDSLx7aCMokG/eK6
fOtxo80hrGoxqcMP8ttXUcE+jYzJKQ4Flk5esFUyaOx2D5By5tFKuvwyQO8or7+o
wmQzEWm+q4aBlbLU9HWGtq/IGwhSREsgcLyvvNDnDHzKranAc8rL8M1sXquj40mv
uge9w9k03/CMK2oUrR5vpTUxWg+/dTB5JJUSpkZJlh78g8t07ORaF2pBACiEiNxk
Ds+OyNsore1R3PHr72TyEQi7YrPITK191bIScYLM5Owd6NblEyJb9hDJhn+bAPGP
mJ7YrxYqUQhxmz5LHGx4lXZ2indshf52fkOlhM70dmJo1gAlGSI/MoIy4R/DYs+q
EWzDN2SvC+QZQs6y2xzTVpdi1npWDkCCikuOZWkVRsZ/rdQRxVZcQG2RkZjTcZ4j
pooBopyfe7FZK0JWO4REU0DCgBjRxt4GkMB+RsSuMfP2Z46bWfi/TD03ezHQBA1U
LOH681l+vZCyJ9aVPagCOWEzgKcXkHLxZ4pdSTtuen1JvRywdhk6t1ikBKNokuv1
x2EzNONS5lw2GFR5AyKw9vk7j64Iq51VJtPv6r2BBNPfv0TIF2Im2vVQi/oyfAzh
FentrtkHTc7zDXQNH7ITV0ZZQVipGLEXbvnY8ofVGkJI6Ik9zifZDjNSX3d0DxJl
25l1/LWcKKU745VgRNCo15uPdRXh5VFzG59Z42U4WfU36E2x7FB9XlVU/I+vpzU1
GzdPpfhzJ71nbTqIfCl0/v9yGAoDpuo811p/QcN4DscCoe08sE2eK+XApP6/lQ3E
N4PuoVO/tFIZudbx3mXTCb/lfuEJ80WoJTzw4sTc7vgSY8f5HliF313B9l0/DCtK
VWAaFtMwsI3bgbtb0vNFedypPC2c0skSAiFGaVczBHrEtsaojfiWCb8nbrgWhxic
7Qldt3CRE2j4VBWS+LASC2m/qRLVFjUQSHcCrbNO5+uH2X06Hdcis2qI6T1Y228m
vrlFJqsBNgUqBEDtLC29rAchrVgx79T9X7ezLgpZSg0VqEPcddV/yujMscl/p46K
CKNoRZ+hAjgVTlfzOPPIuBs6sRsHkbIJnXvXLWL6uvzgiI+0NADcg85U0I6bY44r
r/9q/x5GaGo33Vh0TgR7ZLHQSEZmGxKy06fm5/iRca6SDalyIwOfpOLYPPIs1582
+ZRbxZArboNfny6V4nEHhUrqJB5BnDzhHckP37DsZelM8UvmbuDm3UnVCjuHVGxt
yIwHyugh2GM+ux++Q8WtxTlwBBFBhcoUddBkSOmVnfRU8DAvejmrQuqwP36tfX2q
dqv8cZ6SxgfzN0xJ6PlUPT0fAvWA9t6Y2QXAdGuk+zIMEyNQM1dSSZBgpJSalnom
42tUR19iWDlY+nP4kIEWEpPAgD/8HTpnMAF4UadW1uoqcA2pBtmnO61+9Q22+mwy
gPSloHiYEWeGZMsWNAjWj7iAmOsNpxfKwdJK6aB8ZJKv6i1BZLMguFbkur4i6kEN
eOnjAXlv053DfylttU3B2iVfyR3mABqk8BhKO3Fjt74lFfnQuP9p16JgubS0WZcA
0nxxhZ3iWBGQ/Obfc7Jx5XzBe+OJSLDs4ifk6p1BNw8nD1Z6m2SrwrKdcNNJz/Kp
AFkHTTOwporEH6mOwPO15VolcFY0jV2mPBzUbRmvGIr4e5CACgT9dy3zBKQFdlJw
fKcv8Q4NK6rfTEMX2Lh7gPJCHQD7685zknNIhiyiBifCwt0ucmMD6PoGe3gOq4le
heL35omAwqhDfqCm0PiYNHNeea4rBTCrzz1t0wehugbqHkrMIB8GYlNISkdZ5+de
oMsDxtXIh8KvGylt+VojdFxmrCHRhvbmpCy9dPsqWT8ZBm+BrAg0Kt7CLyhK6lqE
7lyBQ/v6xLeiTW0Lv1sT36HQXMJ/a+Wpk4wQ+1yyNUVsSnZY+4NwXCy73vnagwnH
5ik8ojDkS8QViX9vgy7KQ1y2C29/BKOeSuJ/GreyiZRtTokb0cNXDAza631YsCJf
HFAA9NnXfJChyRHXPswraO9StZ8XS0qalDi+rvf3unQuwBBCBgPGcVb5o81A79Hp
oEOwxRdqRvmyo0ApORHADE603djczvp1XU4YmqPW+N2owz4zpfm/Jr5Wevb8ID/E
SdHSVZ3NPXPkH4+uxQeSrzxSNumKwOx/HA2S4r4VMS+/1UDnLwqh+jdSW7PBaUEy
Vz2dawvahyn4sqzoTT0GGxpMSXWtaGRmUbjgq6SWm30X1E2Wg4/5w7KK6M/ZHmCE
E23p7NH6bHGBSBJirrlonOE3eHY5xehWW6Rh7FbqYFaWxcTfSxfFKX4xbWcZBvqH
EiYYq2FRuC/X0va6NWTIo+2FZXwMmrpu57mcGO5WuRap+HzAgvT3SbSlXZtuXUoX
+Ue7u2eRv+vpjTsITPQdCJApqSrP++ri/QN/wrhk90k46KlHXBXFuUeEPHH/StUI
twP5/aPc8PNdZgQMzWOSNO8d5/TIUygs8ArwaVqaasZzpHZMPxtYKTEQ1QP8Js7t
ccknhL6CBQcf55EuYoaSP01rQet5IErwz3JpHPe2Sbt2a41xAWKHC8etuIfnQNZ7
+IQv/hjIWBdfynC9DMhU9goKmH2Qo82pxqq6bhnx66imYKSmMsT6oT+KviRijz1+
PowPJPZYkCPAVKUWppQnK5IwKlsbQ4Nu922kVGK9GC84e5w3EcYxLfBipSPiemBd
Y+uTeMZ5pgwyf7BbTbZK36WU8m2rj+EEL95x7WhIUdcAMcwaahHE5GilrgbsfvM2
Ikahvefk3SqWc+xZdP3ubkzZC+nXRaWmC8BB+84pvOVsHR3ZHIV3vLkGPnzJWWaj
6TILCSIf3tIJ/rdgSUvIQ7PmSlQZ2gBadf/RDaxG3ejZI+cWKLtlR2BovZ2HXOSz
KvQXAQKkFXvyhlDxWeCqXLuN7Bq5Cs3VvC50dWcZU/ig/tMWZMMNiI+Nrmsg4YAy
g6HDL9szfdD//zQMIMhGU3Swa6xzc3ReboSb2s3r8GnfqUINB+WSbUoZ2LAYHQyd
SEmRoGMspG8q9Nrps0NPu9my0xfkAOGGsHnKhazJZW4JIhH6uk2VwHaOG1NDXO/d
zzn9W7BfInfn8f5GFQKUjp2qnEXgDfWG0lMuXHnEidvi+0ActdDu7VEFpbBh/l0O
MWhvqxPcMmwCadVOM/PScz18Gybukv4T7DeHZJMJnVz5LuzQNoTa9w/bIRtiLVeM
mAC3Es940/SoPQhjp9a5iXXShD7u9ndg1S73Nc0B+XfKj/UHBroPdBKTRglwqpZ0
mCz0cWvFUVPdB4C2wAaqxv4fIgqfPmLjo0LBoyMtKi1OPAihWmxS8p6R7S9aC7Rb
0skpeeKxv0WsJr+qTnX9RHG/k4it3fPkfckH+ILtrfntK2za+RT9RIiHtD0ssGog
ePcVTX9suMWJRn3Br+bLZ6NxUFdoTqLOjH/Txa7h2UAIOsO5TJfzYDiBgVK+Jf06
web5X6ckVUrJfJ1wl9HfEQesXZfGsvf7yMgLw3oDMp4gYEoRJWaH/FbU/6o9bfix
OqmssvQDC0NmA+Jy0zxzSFoBEjD9fKUI0FkfYCEXhYBwRa6eE5QmoTQBJkmBiidL
OSNpyXwNU+0B917vfzmKuVM2d4Q2UoLiHFls1+/oZouJerbO8RGS/5MH1F0I+Wci
6swkot4RxtgIvHL49qHkC/0tHgZ26xekpKTKTdgeR7UZC0aieTD0Rjc4MKg52pMr
soRjYqEFAN17krYfMfrCEWrtwP+w4uaJ3KO/t/PPqYYJgtzAFmbITpQ2ykcdwm1C
1JhzKLdu1SpDxR3lmJdu+/ke24Jo7+HMOg0bVZidbUXQr0WkTdY26PYG/GEjvX3Q
lw/Qkymedq9GJkBHVuE3vw2DWQf2e1snEs6UYYJxehX6B95mclK/hlB8NWDNHfyT
/Sxj8tD1GxKoRCwHJcNdkhOPehciNEfuCqHbtxkY0RnxXyCrE2ua6WMSqbo8IFsR
t7KlTrOyg4VxrMBv3m9mahM+UirJJOiJ6fzD1hUis6gN49iFeA35vkRb3ma9Qht7
Sn0sH4PMABR8EHhx0cH+Kmi3SfWnWEG7zG7Q1sku2WY1DI6z1jXQBG21wBRcZFuC
8flOkDkiuonGPgdqfoBEKU+aggICE8KSSd290V5/rh5HuTY1QTdCx2xJpRhYDTcu
P7mo1XfeiKEYM0JvOzmdoTuyv4facUJWl9pMeTg9fgvJfHLWNFgze5orU2/BGi2/
PYj7MCOdO2t4o0X1VRvAwYLGHtN+XkfOgNex2/yl4152dIhs+PuNmtfJczd9OMXc
5jWZq/6pFCkSyr36i7W8BORqsp3SsZn6kMnWWWF2CZAS+nzceQ65xGX3RsO3yZvg
P2Hhub0oMJdtTGKOmmmV2+yJhNZBfy4m3Avk6BR+egGDWkFU7zLlJpejgQvKT8OT
umTq+c5fXNA9fg0oQaIip5z5EZTrDq8FQIxOVWcMb5bErP1uq8qfSVS17jBjE20G
x8TBcgsIePTz8NFpGERVj2YCn3aQkOLqTilop1R2iR2tGrA8KsdKoBBLy/ouaQd6
bgYnBrrhpxote+o5O70G1vhppzGPQWJeQl8KqbNlkLGERp9Bxkt4lfd1j7KDUWqj
aGrY6b3qnLpUSlbnObewp43vAxB17ZN9/dbZWkAP/OWwWfQPrSB+DSaubgWiNx9Z
tfVMiT2avGa1qHd0Jmp0tMBwkad+Rsnr3KBbjHlYR2JnpYwaqQ0EIehahJV5f0yG
1SLSij5NnxBlwGQsmIwvMmOC32Br39r/1KFoHPW3fQbIRjj4udYaVZw2n4MwMwK1
RadeBqCxy8CrXxssSPzFXzMOTpTI5goJiORxMqKpacFaGDLXmo0TGoN3mRiARaYs
v94SLHuYUTWJdfya4xuN5MA0IUwh9NhqfkjvlQGJTMO/qJ218PtCxS+XRwbHxUeh
GycEL5AdA4vOujuSONzhUV0Tl6DJhB58SrKHdiWH27qBUM0Ur/O+rIJ3AcU1UBVv
SAg78mJnvxyo1GLmdl3Ka4fUngG8rXiK3IM5SJ8lucye8/1y6pdhHcrW8aP3rzWK
tWyOEaTWfADyDOzf89/YA0pn6OD1xhvEQYCiFVfefPogSpdusGh9Msk+4FO9RSI+
pW8vA6DO3CPG1pG3jcfWRuH+vSUIbF6iIpgEXbCvgiUinyIPqQenZJBEAkGnoUBc
miKIs2zcLIFk/qA6fn0YDJ38xbFUJMopDNtxZ6B7pAW5V+7ek58w1SArp3fvWVD2
anyX4POF6NchhNnDr5wriCfQW9D0LHLrM5NCeMj/EtlkO3SxuA+3/zjZ4PApkYbE
fUbeGpMfQzr3lTd9vr0otxKkluDjmcW9bs3bPWdObyusuE+/ayzX2kxesgLXuO26
1NbzjTGJBbBRldVbjXhsJ0eHqxewFT6q6bTIduBMgSe2k8psd5UvQ2X7EYL48uw7
xqL9FzZ3V/L1TbhohzoLCDsirRYIew/KR0ZMVdmLaooC0YCwPXWbBSEmZ2CIB96S
gVPyN8yRhUIBpmSR+UZiqKYJ22rH1boY8zKkSfVlraF404LBqmaHpDEHehtz6RcL
uAc6kE0Ub9sYwOxyksdLDop6YOSVi6/LzJB8fOjy7sxVCZmtakug8h9dlyO7Ynzo
aRzneH3ELmTtKQ2UZgUVMS7ZD6dMOO0ucAzM4nELv78/rc07xEf4WaSzJltV0kc9
Zkvy8jC5qCAIj6y+AcfsGjIjMi9sY11BuDc/G4OPfYTP/PiYmQ5ccpdDX+pYssEO
FyxYUEPnvMI7Mt+mz5FzZNUkFv+GPIT9s3KvdYkhT9Dqxp29KXCygpF6TO3tGC2d
DYoIOccORlv5nfhjXopFX0ch+Fpoz00FikeVF2nEVPxB49OGDXkYGi9Bee3KLvSj
wwRGLM0R9+qv6BQvvJmit3r+heviwHbLWe0YN2oTljgFXBRIJ/UPNkO2d0fm+2ND
ObmYIkXRMZ8nwsYhj6vVe7GEAfzPhcSg6hiU3Uo2uE3Vmlbf2EBJm98obXEZNV+D
2U803DoTw/V6AA/dDqHG1i2AKeDKMMgUi0Q6DZ4ELGPWRkSckqLHvElJnnsJ1Bly
64BlJCOcf5yU8RCS2nPCYnTbN/aKEfyohbBR+oflwdbdBdalcZz+9obFSS7azFTm
mi7gkDhKVtK10jJuCpRY/AkwOdhkVgWNsGqQiagzwqVV7NuVH7QnOi1sg03S7OtB
piKkGsuj7T384DVK0P6wbXCgO+FrdFiHYtUk5PrELywgOH4/3yU6EMpspyXicGXN
sC3nO5yUBpEKmvB8B2AaFdYnSMehk0d5jOM/KymwC2GyRFdIPNwl7f3iAKAkrV26
X0wDorHIja3EZVSp4uW2i6FFLqJntJ0qGoc38Y4nNgcRP96BTkL/a7VJxL8x/5XF
RVKzgEQVqe7/PHo7VDF2mdNw+sf62ZCG3SESP8HpFtTKdx0GkGuGAs41AuUfvQR4
7x0fR/FnrcZTV4jji6e86DE3ueSfnAdmygXk7g8M1Hc2MD2BBAZ8aLy5oxr0GM4X
1MqaZudoj0pZirLnhzWr1x40uoa95BKv3FcL7QhcvselxtRoQifo17xIPAricTA7
XBYic88WhGXnVxgb0Nh6iqv8GV8CMknqHjxEbG/jUKq5VzZ33Gwmg1AkJmieOrJl
3N3tdl2nPFvj+sgNJT4O31YV9t304sTosILEixuUC7dXw1l55SNnvvGMv2Nu0ZaX
4dohhPnOUvRUDGEhaqnsFTPgLV4Epk9FCrEsAag4T41rqgrufGcQG7/Qr3m3Pwbp
RP7ZCnjmPx+YnNxJDZGSwXKT8BvebT3BEN1uAbG7haQ=
`protect END_PROTECTED
