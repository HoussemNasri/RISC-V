`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qyqqA/iQuTRGwL6iwbmr8uuxMwCmRLLGNGkQz+WCZc+uyeOQOm01WNluZiTjFRHb
lLvIAwXo93tdNJts7GWTRMr871iCRjT8PFtHQ9uu1zSQs75bgXWMCcGwX3ayYgfs
AcVYxrFMt5K86gWc1SJ1E4hcdoF0btqGlOQ0PDRv5ohuCgVYGvo1JPn8wu3B6lDf
Iz04Bggnk9K+i1YBvACY7ef7fPovgFxG3A4PSFr47Io+rno21qFvka4aP/56czJ7
Vv3D6dMmqdwxuO2vJy4IvBbbdLndY8HZ6GIpl5HSRfaZZL6dElzsVlPSU8sBPWDD
kjR+cHgnMg8NgpP52Mi1/WPkIREXCV48qlWy44mOq6Da6oqw4oTKxXiE/DyrVmc1
+RFM9rIyaAjLs32u2UiLqcAoVh1Z7IvqN9H6cIdrG4Jw4CDpdAT/UzSgvWJYrTjF
ZF0UHD2aBIk6sHZcrSrL3mCUGL4arnqqZWhiz6HIKMvuo5bQSNOPMrrOFjgeMJ/t
Q3v0TvS4Y56+IuYrxFP1OaH6v2UEfJDryTYDlt2e2MHZTCfKELMs/q7drrnai9nR
cEwgUiPrPoE6y+na+ukU9O135m7T7RbxV5+kGAPQXq2qVHYFArac+dwZJmxOiUOL
QOVYJXsAjJSS0AXRFXUuDqUi9LiNFNtHDfgjGahYMQiBy1NiHf8uVSFOPQq9ac7p
ldovRH4Sncn1VtCeAPesy7F7poDh/OM6uAG1viyp+Wnu4Z9JnpFP1OxDE2mee/jT
UkwDwF+Gq2hI8SKucn+dxVuMpk7V8tfEh5dJBP+pmqJ8/lYMdtU/Ic6Qu0bdhfCj
l2bj2irrob7+hYfu+s4E35oTbm6sAqUN5qOHVT2uEard2icP9LoYW+RdHQhdt31s
/f2ar943uz+QFZHC4dEto3FnF3AaxVGtHvmk3LA/kRs9uYCPU4farryMQpaL+i+4
67DuuWegIa62MRJhsD/HUjSjhSPuDg5LPxml518Hq5PyCh8BWOciU9zQChH+KY8o
BooOAGSOnRtp9dK3QdZQp6HdJNf0Pk3vEuu01NHowRp3bqOIumnZ99Kz2+RePE0Z
xmZ3gGnFhWg6uyk3qRfdaNHm1+rZDLsiWfnEEq8uYgbJ3Gk57dA0Qn0VrIq1zMzD
qSA/nM/9zvkolyDxIFH7odZLtWZcBALLa5u6+ew2xnARLmHOf+87D9UGQ7qpDzgC
5oZbmGGyviFa8yagEwo+xuSwD7zbfCDnlqP4mnl5c2q4GVMmoNX7OXgMeM1i/Lgk
/0O+YBbQxtRR/EZ4bnYnKwJVIb+kZ1eKlWUd2tn4Nq+uw5AjZ+UsXgc59fORuVQN
Nsm5vEjq1HzxU7DtIczvIdEIG+yqOp3p1Y9INNHHVIcjZR5D/pVSRGIhvlSsx3m9
aGPS3FhDiMoPdz2g8VuMZi9ZONE0f9//tIjW6yDQilQwZ1Z60gc6YkDQluWnj+gE
nwGE4TP6NBByGV3v2jx7LgRMFIaOEMBwgrL15+oAugbCNJe+vKep3X/Pm1K6graL
OY22j+KXRpidGKkQ0gCkJkJUZq30KaE25RU0orW5MZK0k8zEVdSQtNVhdIQzl5R/
79/uXDfFiu7AX3hlD0jEybace7THFtO8IDUm2cmuUcNq9ewwfs1CFMDn+1Jt2ytq
44RDOUnv5dJ1qTHAFrPdoB6vsx61VAimn9sxLCByIXbEKn29c7VcvnMYCVTsEkCw
wYb06xQcib9vYMe2hfoFZuS+D9l+5zCgCwA+D3gNvM2QsG6GzGz8X+jX1Ee41uBY
a16fJn+yherKmt6wm4+3XA==
`protect END_PROTECTED
