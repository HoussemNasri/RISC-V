`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yU8lTAyb1/NUXr+zI0Gb5YR8M93UvOSa++NSb/HpbODh7FkAxMrFdxQkhpyzd2T
kQAnKXaiGJTUxEekjVlYlK+AK3K0fSwh53yaBOGp+3S3vNU0HnTM/kPPnyDfQahH
WKHFfGyPljTc3/mK5f1C68kbYhgsnlx4v/i3x+o+da4CQExT4hM4vBREJHL2gKb+
+6FzX+Of3h6RAOPuoLN3zbxk/GQDS35tKnE3HWq8JEyblkqt8GzqZKSwV+KYyW4J
u5BheTn2gI1pvoQkiEMDNArn9PY3Pj/I/SakQ8+PFMvG5f20UWLREXuTtMYzmfDM
Ppwjivat73oiu+3s3el7l0OPE9jA88gPZxzwcoQJ/lXjkc9v1xkVS/0Jn0usF3Zj
wuVgfLgsTuW1fAn6mSRpm1Ra9yJc1eQERcs2vJjYQz3+eERg5g++SlITCPlUWwA6
tBb82g2uP9NNCCPK6B9WNNBkk1LmGKI6cRs363fG4wtSm4OhA8h7QMIRuAbz7Cy+
zrO3gSFAqNP7oaiIwx+DOXAQOEDt5A5YKyp8fS5cuq8XG+11g1x/Wi+lSttU9Nwp
5S6e/c/fr0fWBvJSpDMqFBjEUGLThKkusQNk1O95fkpuWSAiiodODN5LRea/ooHi
+zxcmqURDu4DU1YV3LzKml8MpIv9FhSmoTt9IG+uusViGyxe15BB8an9aiTbBarD
nqr6DGcNG3Vax0OwLx8i9giPMjxFCCzouzzS5lie+Dh7/lJ1DMUen8PbetXEEcjd
jJFQ4ak+3BY7C0Q7XThvhIfFKaFeeI7hEpb44hFc9fLV8GXq9hCLVNeS7nDyfWKN
65O0mNPyWjZ7MZqcTKAiTgB3JBBdn6TGKIXxV5z3z4vBwxeDelMS5S37IRkI66MK
5aK+A7JX9aGn7mqO2DQGastWTy/iZJ/BibgFhprC+klGXx5/AufCPZrNIdlTNVTq
ezu2SkrY/aK4oOdfppNf/trTaOmXnCXbWoDH06w1RJqCsoSy84bU13d3Rv2q7szN
cgI8IGDC3xfdDo2X7DEMGHiKUpi22TMJlWHuQ8B4RgPFUVog3MwGRy6UwtVmsnSJ
cjFcB1nwIQtYEgmn2wFDkanO/Jpmz6IHRDeEZ6N3BIqcCEJC93ez8I+EBmc8bgkk
va2CdWZ1d0bOVK2CKiQAw8Xq3LFL/D6xzBdiuwajNiJG8yFgIjPkoLF+0I/SMrli
ens7n+r/sC12wQ2De4o2yQKkHemv2ufK71zYP8CxjmjT783Mv9WaEYfxfZTQD4oF
RIvZcKPSZvkzPQkfI0+PkS/fy41uOyM0iDmAKVbKDSQLvOvvqbAxd+vkcxtW1fiP
Zi53vhjOIuyyRGrjT60eqqJx16yLAz+VRLxGa6eQZaAPo01jRaCRnv6BS5+L6/I8
ZzVFLVllDVKa4gqPysQ2Q8S+V8kidmkvHBEwmMLqN0OdKeIjfl+5vSkIH4DrL9JI
lbi+YH3thN5vMvAmvfMivcbHsgwFEgrVLb7UdP7UquMRuVNY9ej81Y9LKL9vS86w
85JORwVDpL9qre0zHLJnwEaiQyjaHI6lGh4pUTftBgWr8Pk3m8HJwOpIyVr5ixRS
eYzD6rkggy+l0gYbC92RfBqCkkvpmSLwS55+c4ASsYvLESio9UEP5mpMeXosbr9n
wt7K1/EFxBLVmng+/ys7A4f6tGmRuB/jDHqOwZ0xE6RrLNrQuDpjbHkzqvstAQKA
XK0As/OeEekRTc1LNW5iqsRfBEKTJpsHuIvTj+Jc9zmcyc3d73i3MoMZQsrDfqSG
d0w0UyIfccFHIIKq1r1na1EndV3SdNXKSL98AIohbeMqfhLjKTJYsHTK3Ne1JnHV
Mc7A3Tsjc5aLtKFhof/+xKMrJ3RC2POW8pGLIAoaiqnGHpflpA2CXrh6P4sIgAe7
QTWd06Cfng6E3GsXVibRFWhcuwVVxvYSwnD5vXVMAG26CkEb7ddrsMwt/KXNeYx5
YGOipUNNsqZ9qWWV960P4xChVKuV6Uxbrn5lvmPt4553fozw4xDkhg6KudfruSFq
AI7Hl2QdLVx56kq7q6BwQAPLL7z7WZRPJU3NzzDxddfhfxtOLh8I8/1jyza9anUA
3DTY5CWqZd21mc//JEZpDfBdHyREAcnJsE3wPzqCpZwD6KaCPsqSv0I8K/CR57Be
x8HvEeJZX73FI/ITmwWqI7votJoe1WHap4mtWS5lS5CXX+Y3lo6nQwR/U7mEMvxU
3EbvedDUxbEZqPDgSqisR041PMMoIUMBCWGcvJMY5sLh+ob846upyObOhWL/FLni
Er6VmevvztseikdhTH+Pijkl/BrQIs4tW+31rvc8bhLbjWRlbPc9yXlx1vC8g3o2
ABqXEJbayFGqtBrZwv5/S8aR3HxbUz0/4Ktnp8uWMGkBgHIEeKkaA10SUXmDdyQB
HjIYBdXk3knb68u8+mwtpXZhUASkHNFM+Dno7ohohGFerbHdcE9/f8HDoZJLiYel
pVcXapJKZ/0bG/G+ApYrkhDI6FumLpQyz6aygUZqG/VnuF38N11Eh5gWZJUY36G7
K+MVWeeYZ+LHOB/1j5bTX422XRvlYxgKgDc/paDXlju4Pcc133/fY/jzlbRNkefb
GeQguW6iRTaCrJtVLJIV5j16hXhSYtYUNKhenSZQjbcBANR0qNPhVBTBJrRLnhv4
rHMEKuD1awNtNK+tWYHpLmxEXgPNVTQxfpJIJz3tSlh239HdxtKcdJe+DIeyhSih
szsUvms1OBA9tGsR4aRpGmaw8C8fo0tN7YFXtHduHQXfrhrG7nFX9MZEB5YMwNPb
eMW3jFnZgwPJDikhjPsRLp4hXLKcHvFUKCb3EFYMDJbBqCQklYi8sfunUEty5P+/
976vdXnXyJf2TO5XanlQbhxd7Je0CNgocMbzUK9ytxF4ZngpXeJbVpISHYPSNTY1
Sv3jJk3KcFdMdOinq9RF5DvhRopk6DvTToBcxCyQKjcBv9T6EXwDFK6cVBE+Sn82
mbSlMolt3jrPlWDEWehdznzvOmid4NyNX8EQDoCtIuZyz07c8DQNIJz8YebrgMbH
ODXUs/DVfMCQOdjFJIusEnFjBetGSmmKt0xJlgPe5vCNMs8ITGTaxKtD+OHm2lPV
JDntFLxmxpyPkzcWp7LnBs7SeTcun1TgTvGn975l6DL1MGiwLYr66MOaKmrmrIKr
q1V1OIvnwzcMVTYEOtKBKG1TStiJ3K1Y/3GwW6pJ8xkNQI0fcGvBqVIYU3V76Nr8
Zp1p1oxAd2+Y6BqikuN/lHRFbfrPpe/UK+l7M9620YHtWGMcRatkpcqkNejQnOQ3
MCeXgrd+QmjCbVe3euJiUcLERliERwbPSbPQi9kG20MdfX/egKWhK5l7eePvN9+F
2fgZYtvN7iVGHqMOAR6wegEhPMc2V6W3i+0JACciREwelDtRjRjlR9o2+5TGBaO6
XmVZ2tKl5JVDduaOCQimWjrT61/ZZ7jz/YJF1Mm5N7GhADSJANgk0LQ23+iWSV9D
lTl43KrRUJ1JmCLty0tPZYZMK/uoFAENMef1ExlCh+XyrpKtP2cfX9ZOItJKFoHx
m8CM4PhkoAYchDnlwhNq0NHpd9uV8fO1ZcPzC5Bv9j+/miRcg59SwW9k1JRc35+W
XyMNOHtXjfhsI6SqIMJHtatvRYgkTW3ACtc9BaV7ScrKsUdI41WVJMTs+L0rPv/s
Au002viJ4oT8Nw5KuI+vv4YYjd12bJLNDzDMa0RPqZMuqV0RVcux4R9ZtD4zg9g3
mqa8wRHDvslZydfylKbp39zKq1SUlNT9gaeXcvd877B0KeTJQ9U068yiB94g6+A4
tERMyz2mBCW+E7JxCCY2gk9zuq+pJ3tgmvSm1ZJ5/ojCRWYlLDSMQ+mSYY2vvN8M
ljN3QxhK3W68ZeQwxB8/3nV71hyHOfm2yaZo7zQ/T9p9AiINMeChvAEB8f8dzwNJ
hCpiiM3rSkqxs1XBbTI+ycxUcKLCCrP3J2MWy1Gf2TDYJMuts7/hJ8+FKvzhwFx5
Juwp9itCXclVA2hFeQG/i1Ta1hHHudrAugFNppIQ+ipHeWi5ESNpCwzzvkCVmN0d
glfbV9Uw11jAooU1DGgi43qP0kaM2Vm7Y0jz4Ts6iR5KZPQQo82f+q05k5zinBHD
SS+p1Kd6fPEJYHC3minD3dMZNd8hng8RR+SpoKGd/piiU8T3tShJa0MAIcfI/eVc
TNSAkahVj1bcGqXT4CjxINYSPtx2O9GRWv8i8tPH0eBBU1mpWpdPo6QZx61a98nc
j8fiE8+mvxdAfKPNIBkanx6Q+Nfbnhqv0qJR3/lTstfxRkRqHY12gzPnIt8QV8O2
aQJxSdZSikMfKAGrgCI93LQX0m3XMmYURG9rU2S65Cu7nfP/cPYiWS/XyVeSTVWf
noUxBHPmpEt7ZVRubFtPmboFuwSBHOTbFOh11EJhfsFo3wNJrFzocQRJ1UzzxNXt
KmiwiNkqFP+9L8Sxn4cyan/LykWiTgn85BjDWr4fwcBJNINsuLynIiXsKTDwhUcV
AWHAVaHc90wPZxduU0l8QLVEdHF2DTcMIwGnhp6JzikMY8LZZ92Nr91xjmeeuK1u
1d9sLA3iokLL9BCJUDqy/IIN+DAJYRzovjkp1OZ6CA6acsIHIfCF2NLcAZ7AHwXm
3RQ/RW75an21Xx8LKrCViAKqcEOYcGLv2Ttq+nRCG2JWZjjbjYy8p8bU9VfRVNd2
c48gdwzbRFvzHgcobL12aOFQ6Kt0ieouv3Jtz+lMpTCj6Lcr9eWf705C9/PVjtF3
cbAS2rimZupXa6j4ODqCNq6AdEcGfn2p3X0yVZxbF7B5TF4+QUhKrauqmVxPZCWg
Mco7zrA/tXMBs82O380k/I2BWxReckhy8priZ3HVNQOXeQGQ/IOwSBBSJw7HjUCY
lAIY43TwdYyG7LhqQWmSeEF5H8lL+TJig06gISpgPhJwPuT8BBEnnkYqBfi8Pc3y
PuZ/joL0k0Nob4k99CLDmTh+XzOLY5Oaq3AhfQ3yM0AhEZQngaMwjerifgvXUrf9
sM50JnR1c8PBaHdCTcFf1XinJRub4UJ07B3hJ+Plz3zpCeMlcQgYHkel5qESpQTC
TYYSaR6v6ficPmcut8+rSdSi5CpYdx1ELz8ux6dy1t2urdGTeQauN3cwC0+Cwwes
EFSH/frPbPwaZiu0yxgnlozY44hYN3s/NkB6boutO92pVqFkeYjBrYc99O4AC6YI
WP+XXuDMczZwCpztGGprpVcUb09vwTEC3wryYGX5b0YGRBBRh2AIdkRshtylIesb
CnHPfwo3pxNfu6HDNCt/ZaRk06tkhmslOutw7aoxtm4jn64g0J6/r/Ou9Dq688bL
SLDdD2b9B9o0zlq3FcK3u6+1xn0a51v+IpltU2FczDAUD+CpSCJ2yjWC91z2Km6D
XoDQS0wZhZkrhDl6xHeG3T0xqoAoaf5tWOI/gh5m659fSQw693IxgwP34fubad9e
+2WkUXFhfFcx8Zzmhmiv2a38bCF80XqB5068JYHG1QCKemdxA4aoKgBjQTkJ17GH
RXmh1VAGetyyiCvFwFWe0LDg/fi2MghNQey1ina7qiAQC+f6rDTckPDkmNFj4nJo
YalmRJtuo7r3hEmxq/JtsDDRLJqYCZpAE0dDiFLIxS1Lr+kvL3L/dVZHzRcLbHMl
HlvMuWDdhp3fp/e5MUW1DjHXRiv5046UjaOaxzX7ATpy7FqT86evCpmsBauUAood
cJgBbTGRY9j3hQOdmcMNjFSg/8JLVFMfRp8ye9jmLeIc1wefOSuUv1OYeHw2pt5y
wP4LQiBiQPm99/djcpU+YUXf77DTdeHPw5/zIqXNnXt9bEJKFvX4+K5M0Ws6RLzo
b0n8kq5RHNuO/K29DzVndRaPlKCFFbLn2iVVDCQOhz1EkPJV/OOIlF/t7/Ef0DT1
h5J7PTYF1WWskayjfzFXpfVjO63yjozYS3P6XKtWsZwlvYuREJohTJAAwRVeLhD/
wHT5A0ENer6g9zgvxHkqc38rgTvnY0rVxo+h/6iPr7jJSJ7U3/qOuX+HFqmH/K+7
QFLyoSL5ucQ+SGtJcxOf2egR2J00V2YbU43+fMGwjQ8kCL8Yyap0GtIe7ks2z0xD
zbzVHi73pYTM03migQTQRWFbXBMFdT2Y7BN56kq65fTdPCQMk6bCzazhTXWtrUi2
/lczAuBxlYqv7W9wwLPEdLCVNyIkGgK2pVzCcTuH35hYw70VnXQkqolLzAYgm+J6
xL8NvXJWQPFIV+N9pJUq07eD0sTzZJoHNrxoEmRHMZD8mf6y84LzGN+dYNxJ/vhQ
NYXQbgpZxIdghDlGtVY0jPKid9YPJQJt8+cAYk2rcjwMqJBzVFUNVLo4Ox/LRfB5
/6p/2M1jTXym2isrQxB2oPay08MlBH7wWsnPdVc97XbYnvY2kG1hyXhMb77s6zX3
aHbUrueZkG5r5IO796CNLYNocyQPPV445+baL4YNpe53+InAXEjUAf0AJ2E2oJLm
q1Eybol1ggnQay0ruF9FQ7DrxFg55ySB8+iW0SCYvC1Fpxe3uNO6T8+cdx5HXzLu
m5OGTS1s0NTnqGBG3iTIVuhTAEglvjVCOKWbhbtuAiYDmYtCXPthKXleRgTFD2vE
255aOxdYBHgLWMgbltvHMG+7SieqvopeydeC7zjAOC7Q8mqgYC8cCctAiNm7fZTv
s1roxm1jhjy3JL0EapAzWK3wRrzmin30hbUvQH7ntgvfCID3Sa2VXQviQS7EhVtd
Xx6sgZRLTXeuRR060JIJGeUvw56PdJAaUIwrNV4s19Efg3qmzTvPI56OzKQGE0rQ
05QGS9hE8HbfJWwjrx2pAfJ/FhhHZNBVD5oC+ktIt1yDanF03SSzA9fw24/th5Gp
DKyAcWOjD/vxfdPWQvx2bkqz1gIN41ezUjb/UiecfhunUHRdmpGX8RUlVeFd2XYl
2Dan2Kw6AvaEVz5fyRQp+mFWDdqVI8jfeMVir8t8GcIFnGT3Bo6WQVhde/C9Q0A8
2eDP/TuGJ7w5QnugWZNc/BuI4aGP+HDtjTl1vD7NF+kpV3/HqHXnEi42qPW1Y63d
VPsYRnMr9KJen6CSr4PAWEz5AlyxYiPTemNF+DDIb3OyIk5bQSys2s5nH+FvtSe3
y7iHE2yQ+NC2T9EWl2Zdm1tXIqRb2MsmLQdUqtu5fJAjVBNqqr6isTOpvMrM1S25
tsjyiVa2WxtfFafmIrg4ze1MOpApnPKnTVhhMCpMp62rteMt6MZj5Gs77tZNDDpu
DYR0DJbul8JRE/YFeFSHRlhJpPxvCX/b3Sc65Ms3lfcD7+DyQpgHPjrvMvyYlIRt
Qd21SAR3r75dEAAArhk5nnkRFJlXGD9ji6hv19AqPwF6iepuIyNPZEM3ZWCuFkYi
wQyefRmRFbNiW1LegQMiHECuYTlUem1ArcAstnewPIQriWUO7sAWIRpivuIX0h0w
N7YHY08bJYrn2mFgmYFBo+NaW+uNgcaOJCwrbOtHNhgyKzplFe4A64CL6i5wnjUv
ZTBIOP02H54i3jxNDA3QOQB2LqUIfoJx3rlriBXgsWoEolAmLJpzrfMOX2rwMVsz
ne/vwD/NkI+evAqftrB4gnFQ6bTn9Rf3sPSfGCmtTkPV/DTqzOfX347LwJFA8cVF
jl0i5uO9j+VUJwAfkC+6eJ7obeCoBEleJkYckdYIfjQLY2PpKFy3O/lUCkLLqyNJ
1y3B83pXI+MW/S9T4gHOcoufw9R7mx9S2mODMRBjUgEwegONn4lJq1Lnv3wYe3Kw
Ghk/gBCfTkvAb/2V4LgkNQVXkPzQb3GZWfjq+PyAK7Mvk101OGTRB1i2AZ/tv6Ft
HBa7B5L3xzv08da26172jl2EsS/BsPwEsWgwpYiAJuO4l+JoLkBcLQx3ZUWoyPwO
H5Mv6EBa9LPZd9JNhw7joT9ncErvQ4VxHLGVVVLr8me/E6jDSFUC28MChqPcTowY
AIPoqVqCAu4Jk0iNHi52dq0+yvdQyjaJAN7CTsXGmFG114qENlxmtjPibLI4bsYN
Vp/cdlW5npeocH/q6usyHN48/59o7ZE7cQmrm2l9srVVRtSen9sFDMCrKqMbThDp
M0jRrIOLFeakQ5MSmN54ozl1kAh2m+bIx34Nb2XbGm5GSPaT+1ZJRjLXUT57caJV
hNK/7I7oY7UBVewGGieYQcz34h/c0OEeikh0/u/qp72G6F0+fEIkZ+xgSxL8X1+r
jGOUIsEqgaVUIlKKeG4p6ehouJifNAzroJora7yeBLW8RCxu9xclSB5t6Qd3yZtZ
U6zYWKqy8ww64StuIBy5I4vt5HvOjGSrirW60FGFGv2IQjemLjPkrL86hOXtJ7Z2
Q/BC0S1HgFHulMAg6NTjgLhtY/i3H8uf2J1nEKhc6z6H3mim3r7grQMB0aVYQA18
Z4U8TGxxW61Ao1MySSQFM6XSWGRTPDqDYL77xKXY3Hpb6fLaIdjCA08uGbNzXYDl
u3fo2SX0zg9Xw0Am7YET5n5W0CByckCNFX6ACKCP7PuRScW3hwdqn4SYDhtHlXlS
nbpmJquZ0BmLjlUKG9ng5g0lcBV4WD8CiNuTJ6LAqLbkgzers8NqeTAzPrUrIjES
TeCE+35CqncOvIuGt9q/UeBAj8kpqpJED/QKFCqLzecxp2BTD/e3pxJAiarNvspy
ur3C2vdcpW0ZZBq3lu0kt8rvc9/onFej6DsJfBM40GZb1nPql92/5JMXjhiJZ3GI
ztabwLhdBcYvvTHPXmEgXDsM9tt0xBRaDjvW9Ra1tiuRU1qy8tDkNO8XG9QQCBxG
LaEGbC8k2AWv/7i8t+ekBGvYyvJMa5L7cV5OkdvXNt8FyacI9q/ucDYi4J3raKu5
Z+yTtXwzcRzknv6mAmniAN6NpbaO1q8g1ix9gpeKPL/dj5lSxtHW/8N6b/4tINap
aqAN61B8SvJKGbZ9YfNnrwtCvHpReKfZXkJMiVQ6Fs+03Ty7FFFgtwBPzisx8Jrj
XvQc66ku4tVFEhcP7ePRmVNI6LMwTfF1fn3vWmdhjVS8x7MamZewGmzypmI8/5DB
IPgOm1yeJZSLxUesaUnYxXH4Ma92YQj0mgl+phOiYzX6fchPX6LYDT/6eHZgq9Ct
NP+q44q1x/8E/dmwNC4SpEXElwwWMSbZlbLwpjbWysBlUkFwMz7jF+ECcFzdREvR
AX6selB9MII9oVH47cFNyHNFyucgEENF+d3FKeJK7li/+hcJ2aUDzLXBJI5cCDDW
Ju/b2j7SXAfoyoitc2p58uwFZVr7qXvnaJSXfg29pQj4pF/vviyooxILSoGzoSYj
t4e0fIjQkcpGKHhui4VFeDWqoN8pLR1gvKnC/+tneqN8RZbBhKPL1w0n3GKjNdkZ
vDIOgnCIz8OOh0CAty0s7yKUaRGfn8yL/i+zVN3fGeeQaDQoRcSpbu6LiMBe9S1C
sCKyomALmbXGK+M6x/22cOkuVGe4u2nqboOBXozy9W1HOjsHGbxnJQftGwv/fC6X
3ME7T4KSkzhfY291lG30mHTCN0H7boacxlKRhDVViT+ThQXPueJn0L8sJQFjGPbT
Sh+6F9TW03MirtWlJ9+IUbRWffebR4AeuhfxSWC50WMKZ483ZuCWIsyhYnOTieGQ
F3IJBBpFq1+ZSs94JtXKnW1WBY4HE5kGzJSQs/Y/z7EuFpy3zNNS7JXEfsvE/v+y
c0zp/l9rZ7dJl2LNW9OdB192GtyqUeRo6f0dzP3cZr0cLQ1bubUAKheIfiEsP8JJ
CbqvIOZLtJsexcE2wiZmQ42/deDOHf5vS2tuSZDUyxr/i+TttI5ByBiIbgXcatPY
MqUYAbg0yh1tLatCavkC/vK1OXwLIQ5LXv36wgLiAT9MlfDNCR3FQ4X9dT2ocDKI
R07KlAWpfUJGd8MQFjROCD1aEDTGLlqfpitqyIJ/A4hXojd5Db47N3CWXhqTDCh/
DI4UG18yMGZGbSZNqdrqWs0pUr7cRIESzYBDe6QO8kZbNvff7ElBkMObyZlGvwRn
AhiZ+HnNH1qKjHeyPlP0fQrz3+u3tjMw/l/vb6bRVUTm9dlOaqFoWvhkoHKU67oo
REMXPjCv79s2VJVCJeesrSjnBP0I+4Rokd9+UpUyrujOOte6F7ghFrXrlJ3nMxtz
8BBNhAUs4dXTr83RKUclUbzX4vCYMcg23I0dxtKoVWfFFNWyoE/JiWp9I2kfnLcu
giK/7XaXLPEztjKgMBWBpmOf7eZoKmJchCJbb65wwbBgb5lWkkfYU2YHFIjmX+/K
WoOkr9pA0KQBJBPZnXpxvWinmQI1rB/sm8Bbaf0FG2MqpctMMJHDjhm+k85A+J1c
/dqwAmrG0/MhKJg9f2aR/YJPqRnI+le4eKKxb8UqBTaMRTbLAPmOe4fzfF9v7z+h
xxg9SlpE+NhK7kfgZAN6ERIVeP6nigmF+wiCz2i6xJ5Bl0iJkVicLMB6A1H9eyaK
RzgxTUoNg7JiOWiE4JdbvjF/qdglOyGaXhmRRdv45GheZTb2oKcfsAkUrMQNSMuX
wDaRrbd//6mxYWhtf+7lcUEJ9YHgYHF288WaQ/bhgmzP3rZsN57ldfWDNfv3ktTZ
tW7H0xFu9DVbVSZHOEC/3YLYdkQe62iPrY4ixCSAhBtC1zLVlVm8R0g/cs29mcnY
P2oVryE9TOBQNw9Fhvsv/rhPev2DQoIp/zH7dfM1cBOmjMM7bUuBR9lZ5jbDRpDN
B0M1nRUw5AsvBz5J2Qut3vdY7XRbf2e3ZtPz90WLa8vEhWCUybrpfK3wDwKy4kEe
qgldtbT/unwzYJQpW7Q2FdWBrND8ODeRl9QNcnoFvrSmzZtkgSUoK14XRFMnraXl
UhrWyoXUAtcq9Er4Oi/jIN5MtT/UWjKJd3RcPhCXNhkz/1P8Kvs+F8nNxbq1NYL0
7+QZkr0Jw9i6wesHlliHmhJYOTaKTUKI5+vS7TxDyHDdsZBIvjgUwrmcQNPuGbde
0XfpzmI3yrGj+lfxk7oynt3ftCyaoMJPfiKl0n51PYm3WT9owYJAaFjn5f7wJbv6
xsWOj0F4zsVCKL14RUQt7raSK0EfQHfnOn4w/hETPiABxEPGxvO2yPoQjWuoIayc
1p1WjKww1LyljlVQWccS+h2CIZ7W7AF7h/j7hpSFELwsJ2abOPw520TBt3up1K5y
FCZMVMTu138E7vE/ovCSQYTsHN5JrEP892vaqYO/QWRF7sP8ALNH7qUhmJoIFnsp
vBf4Psb5Lr1HguKBFz1QjFKlbMe0hObUrCeV3Q9p5eJEEdslDGv9KNZZnwsOTK0Y
c2lx84UEwmdH8+uHd22Z6p0vW6f+ETh1GGd4S6cr3CzsAfV6Q0W99oXkJuRD1Ca4
Mm/E88LwtN1uEqz6O717AxDprHKmDqOcHahaTQ02wRe2fzUffsOIFHQbL4WkCWvw
UeE0luRBShoh/8LxJ+QsIVUHTX/0T2Mc2jYSGpSK15KkDnxeWB8PuoI7QP3IRs89
UWapa+D+3kgozw8uKIVp41GD1UvGEwPn9X4hQEtHZe79bPs/413Xr60eyDPB+YYO
HTmFmEzYba9Ak53GtBKATLdVln8DT49VKBIRV4SxIV/sQXXl8etO2VXPbmgFe8pu
tgaEmvvXAmB2cXPFQpEL1tRPWQiOD/72Zwwjss0y+Zfvmis2xBAlG4W7p1AKRQbx
CjmNMOdVTqGnLE0sDTZ3I6UqdxvRLa5KhdozLySwTjMFsCPV04OSr2ECr3WXe+mc
6AZRUwfoBJdn8eRHbHkrGykyRUqdR7QiMviQJjXozLfwPc1FKOHWUr1Pfe/rWxTF
3aXZX+Q3AiP8rdBvdt4WdRbDnApCx3kVcdtGgh7GJJssbSRCLV8cW7HH08NdYagk
DzMZXdrzKKxTpf421C3dzMWSgBvvODRzsdpzjLN4xtiynmRD6DBJbSnhZA60bdM2
kFaBYBLo13IxSpV46ErGTeoLjMMZwhDEaOS0kr70mYIzaa5UzG3Mblv2SdZJs8cO
en1rT76HQKaFSQ3cof43bQHFfE3v77v26TEIPPW8K6TGbjL3Y7DBxjmZzpN2pchI
kl56kX2LfXBRvwKRT0XmqEZB7iVzqmqVtuEhHs7cR3f+QYKxak81433PMDS3qch1
kFdnjBIH2BK2tcAvjfN1DaVCwZ9SdumlWFZcicDSpT/0vum6UtAUiVUZu1nZn5Eb
OluotPFezXDHbT3kI+3EOOA9YSka6tShBfuQ9sfuNxx2nWuNCwi0FQg5scfklVK2
v0qRjAuRRoJxG4bsVvqYThNx37KiVgdBlhODZkiWrDq0hDl1k+DM8vkb+bljPhLM
GsSX2EfTjgxeaMBKKhgYI4Thx8n1cBwEpgEI5C7wXdCmbojI29mXA0v1zZsDGBid
Bal/pKGY/ivHUmr4w/QohwoqSYMu4hHuiqcAHlki7ToKlHRMUUMPMNPNezS+IcYI
onQGJ6UKHiTVVpjVtqyOAAP4O8OUS/198JnrCyGQO1LlHzgLvaZHsPA06+6XHOy1
k9aLGCLoais9dddfRn++PqtosXHMBnxb1NrPU2MeG/SGwweTp7UTBAmrzOCvH9YE
mYcnEbmgxGAy9sctYKXCumqXQg9RRhTB/vxunYaG03Am1n0sOHTVT6wcQnEbu8UY
2XumSlIz7Q0WtelnY6qMoG6wVLlF90jEKBqPAsHMeOgRPxfl6yn7fCg/D5hckM0L
Gl0+Gv08gel1YqDnFgUOEVp+pK01rM+qkRSeGHllte5hEhj9RQ2HA3LXf+S5bFBG
2M0hksoufobJ2pXXmaU8PYY6YaxWaaRyJTaUSzeljiiikPns4+VkQB6XWpaXLifY
Msm2oIbnJGxqDxH7MykXGcQNt7b/d8mepm2rpW11fv1q0KHYEsK+VwcYqbGj6brS
k0UaJwAH/qv2zwi8ygawVDMbJr58N/SMHTHDOwjw6/xgQppYg+7V+z3s7PUW7g06
nKcedDiTGF2JvAjjiXLOdfbpt16BbTNcEHnm7bDiRlEwSq4k6Q8C6p7wTJpx7pII
E31fWhzK07BxzGLTZgT6Cj+E8O6WS89frHIh7L9KgLzdf1WMM8SawOW0ArV3CgbU
YI8aWH/jZzBJVx03OZWTqN6ANIFim2w5FTBcx1/4yJOrTRUnrQGioaAi+tPGiTo/
ZeSV09Wv2B0trXi6ZwytzZdDr4ZB8+MbPZY+ylKKUkujL7wnJeZc1ZbquaP2o05b
4TL3XmiITrMq9fl+HZ3QLGP09T+am5dwGlmNkmRGdpZAlklM+rK7amh15faU0yMR
xsppm6aIpSbImXqDBPhJBVfWaw1gPcB8OD2JHya5Ue1EKCm01o35fQF64JN++IgY
dmLCihVaoZAgSdlaReBLtGFzdrJzTlsDgj39VMfhGIkxkj+PdbH5KBD9e3GFKFI3
KM986LlTr1V+d18CoC9D5PiEQhgsUMLxICycrSx123ZMiJwdHxu3l7eipp4bOXCS
qnP3wMgf70ub8JRoB/nmObSOnC6OxULyefnbYSSFb4b7JzuOC51aJkQsDWJlhZM1
OkPZEqCnWfdUMZfR8DKYjGjoDCk1drHWzBPLNTvex/1uITCRwdCWJzWnpCKPw15x
zt5GzW6jpS/1DPjyb9QLc6v9nub09cDGPf7PbLkrQSU2PPSNaWvp0RM0sbAHAY6w
IG4B4sjpqTYf8xKQAMNzvNLtD87WHlWM1Tm0UuPS6yTJLVwNp+pxaZWZM7TjDBeP
7FLHOw9ofY2JfCUEEFrLh0ZMvJo8IeqTQlGpe0S2D7WqVIms0uIZk3qs4A5qPEpg
mGWwpTy/qm7T5idDLYAYe9kP8dsOctCm1bsJiuZ+PkxsYkSVmyKuhG3t4SDbGZgu
TfZGpvwE/kwNbZZsg6df8D6QOrIEqJkbaael8x15Vrd+KlNQUnCSFNT5YA/562+B
lQaJK+o1Y0xgp17nygsORwzcQfzqirF79IRJH9d+RaEZGym6MHUhL0Kb8AmSWsn3
p3rVvXHkQRJzxzW12m9lUWkk4svLOXqDsVgq6leRH/MDSx6NnNV+xdYd65Ua9J6v
WkBnHGkkUFIJB5vKaP0TUeyY01sZ6RmIM3ms3TGNumJibhVideGPny0LSlzcTniQ
WG9Ur3Du2wboH5biIFttjm90SVB384BroRrrWeBeSnQP0S1Y9zrHkw/z8+mo62Fj
ePB1z/gamxltsQRa/ErEYnUMORJFqXUTp9qbhb2dQfOGK0IoOan+qUggz5Umf9xp
cMBC4XZukv9u+C6hYt5FFfX0UfAqMaY1kQUcrHt/RHyNrka1Bi+/PZDtXsortTJd
pbeOE/D1DE0Hc9Y0DbyEB3XqCcJ7nTGQmfXtPU1eNMbH6EnP1PkC8FUFhTgq1bqX
KtwkRFmaS4kzTy9dI/zVAv+BgAAHSejxjJ3F+STELzojRyfhfn8CJvtBBx8hqpF/
bJTpltpJaciN79KQtMtzQDYcQb/Tqyo5c+QCd8EqEAyCVAe7BBeN7WY0H8MRvjWB
pBF0PED0TQy6Jm7QLpRtfrTuaM1hfh5xhqT8U93NYyAze1wEsAZxIm1fXEggOXIB
DN6vn3koLr0j6DvZ0ZjqHvJ8MA9iJypIiiT0T8/f7KmPSAzDOmkFN6sRVd/aNseV
InBbO+R3xiQ9565Dw5hVK7J7n/tOm2gJEanZErRUeBEnGoI/98d1aR9Ue1wud+vp
F5zksSsnv4fb1vZ5rkeDZO/v0oGtnWfXKrmTtcdNGXYXoJQ1s1/js/BwX9ek+2oM
nv93XME6CSnvzbiOoXQh771bt+4IfE/ytZ9FLa83SplUCK9ZmLPsK7dc+opElll8
oC6IvmydRGohicnMXMuQvYCj/5EZKiyGz83LtefpVvDXLWZqMj4th+ONAqS/BZxt
zs0w0d/MUGiIwXUkWgMBb3FgG8GncMvnL5NvCzta6Bg7psXHR0oJaTmJHuiTsYuk
az5GdWE2PmU0kuCUYQcLMlw4G7/zCnil/YQMJK+khA+iyoVt+6aYF+Ea/lQvR7z6
wPxnn43dS79jWmhvgofcwIE4IrUKZ0QpHQNAwVvTBXJcDKzvJBWCU4MZgibgOkpD
vsWzbgRbGjE0SYPYFLIoMSWfZb3eU6HlcutEyjZ2m0GRgI/xiuOFvUCsSpPNFhV7
2/LGGC5FAT2hkBggtU+gykY11J+pZEXilNEdpwFjnLyWycTKTObdB1Kz/AYamD+1
6SX0QMTnKLzifY18fCyGEXC+Cnsr4uC0hboJwrYtyKr9vhVxspYDtdfmL8QG96XX
hyGeYFc795AGsIC5HAkV9vl9jGfNv2lv18S+a5KcIljpyZxzwgjFGNhOK1SR16XV
csliJAYkuB/HCPLoo1Jve3UVc5voBBta0PfP7LPO9+TElErEookgdu33yxnDvHwQ
/fn/Db6FBRYyeMPLeg/6lTyar5t4krq2VwdrlYGUHmPD4VTWpmqcB1xXwsncXNdW
lMN52+dGpJGInYUS4Qqbm1P5LNHmiOm/utcidg/vSPwTyRDq9F+O7y7UaKOqswYy
+90GXZoA4EkO11BiwvcFAaGW9efc4f2+rZ/tz4am9wQUwFJ82tVPCH3A1GMeKvrY
nvkb0gI4m6x9s02tTLh03ktP0osEVNDMWIWGQpcSjbwHcWTnP2/RCtnRkGVT2I0N
fPdUepcz0hXMUhxFA4Qs7PlU91KYCdfiY126TDvtFLzbXYhBGvLXLX4ODRPB4v2F
aumQrX+yRqYh+5GDFBRkDmUgOHZkZiV/40Ghp4mHjpvVBlsE8P+Ses+rayjqot8a
/RQJdVVwQfbSrCJ7jrMOqa4LAZsKF4zK7xhDEEBpcajCB5b1dS3+qCgM4m4/6gp6
tLnpyXNKxiSpCN4Ej2VhNvtWHP1uJlDStDD8w6XYuO/u5zskuzgoy2tsFg/2fIas
vf2156LhHUyZXnn2azOTt6v8PIpMLOpYQ0GCHNLBoO6tuivnTgbQdsOQ2lCpMNPv
wCzIyLnCXfFjQIdTPlZdZSMqIO7LR8yeB1g5ejY0sdj3ZBIhVsytApxS3dnXbwp/
T0gWsdkAbc2ME8JZUbUVUeu4+C3mgSSHJkgWW1aa7hDtEnMrSEp4gWllqdo29x9r
IfG+qBR76ukJ9taa+qbRqPdP3cs5NoOIwYBUiUeXxmXb1Bao5fue7rT4Be4p6Qug
oZ2NIF8jgWMea1I5/172edkyq5Z/XwCdAPqp8KdCEr2HaEH6QIHPufMzmhgw4Ejw
8b2hjoIR/xUJUWO2cKxlvyxbe0wCm0w0leYtwnQdu8iKOtij2u0WiDUZtI0NW1ZA
+ZOyNmwarvIla/jS6gI7+PNH1Sys1yWYkwMPw4t4BTAoJAt1IlHhUJT/qk5Z6OmO
U3TVlE8YjrC8YKspPA8naueXcDEYJiu/psztUrMMntJUCYGLA0L3Ub1WRCPuYPld
TgoFpJt7ihy09DxUm/MSi6omRh8oftZ8ysG1jy8yo3euv5FmpsvXxSjWwz4/LCCb
8OokK2zc9vCxTYfwxqwBIxZdBfYNJBkVRv4NtYTBXvmsIMPk0keSiF+9MjiUjfkK
XX9kELywG2Ci1ociTF2RTpjn0o4Dv1ZARADhZlCdsokybQWQq5QWJD6zZYDO2mE7
GsPHmmoHLYaxs5jP+Gz3KVnrmNdS3yLQgfE362Diz+zrK5/2XR0LQhHzS/CZBghH
WTsSRiQsrgnuNyUBYZ4b33ZRqBCksnRy7Qj9ZH/qcFAiIbSAyhPh54bCiFzkj/Rm
hTqksHfcQyx60jqJUqDCJpD6sbLe1Hn7Ex+KW7JLkFc0ROqIOQ6X1RpLRjdmjAKU
7//jEfCRSFc2VypdmOU4PNMQJAXz/cEV3d8Cs/AePSssARwuRUqrcy09DeitXhEC
fkqRLFPDNTPosUZC0X/ASxfUh8opnx73PeXCW25NIitlacr8r4kfDb1ZLFy8w+3m
Os6asGaVNmW51jHqN5MI1Mee4Sqr8UzXST9bvllqFN3rTgiVs7arHfEfjlcs7OT0
8grVu21tATE7W2bb3zqvsTLTbHN7YqTxvqMCOaObAojfP33Gs4MT4p5jVZEkvdGk
zashXshxL6DaTsXKtHgwAP+ieIyoA8E393zRVBP7Rpg7IDzb4PnBhgO8oS6FnfiH
BQa6lc4NGKCHR9n7fzyXa/Wrv5iJahgntay/HFM8GD2T7Y/CKzwnP0I+Kh5ojFAS
DU7fk7L20y8o86SNL4Kslz6zkYV54psA9X++cBrVeRtiFZcBsD+ABGFNc5to/DiF
0F6jdjxFcoAqfyDvACO7Q7xUkgYHlULFoyirf/4pZSKHDBujKGHnN69uA+p4tR/p
HvAtgjb7cxnzonWJFYwKqAsehdgqWzxTNhgPR6bp6FPvMU/lQkpvypW0/r4lFJEz
O/JIV17R/Sif1Hr0ednoYbdRtYQo9ufyZxvAVNY3tMN8paYJV4tyIJFdjSM9cawe
wKkeWfL3/OsdgNSQjmf/aEvgbQVg/HIg1UD6b5TzmgfTnwXKi7zy98JAA2jEjHbk
wBjMx9mNyAfr7V0BnUCFkh7lzU7Fbh7BJ013EQvJlZMraLBvmJzUMsWjiQbooPSC
F5V7vAnygZW7JfGnyK+MTm/1Q2IOcFVp/qIEJJOb8ZhVOVAYb0BLPfoLAVbi/xFH
PXaGXKfneMpSIettiK/Pvbt5gcvZcqS7eOKEFXvTB1ffRNwy+x3lFm+wWnLUYty3
NIfTuPedPuI2/NaHP7oy+mk3XI9AvcPFLbcfqYoQY2z2gYK+x7bGtWQDdgjGnOGm
Cp6nkGRN8e7SgY4jkzcayHgJu871zzRJ9LDJ8CgIHjILi6L2Lif/8etePmlv00Wd
qJssHbNXYuxHz69pQw3THrSqV+DkjCbedGncFQRrKZ9Q1MDSc8q3Ql9UYBlJgkAU
m7uEudJVvgsbYEPNuCq/VVr8z8ZXuph9UAnIKYaRUtMLaNdmPd9FY8yeWabGY2kK
trOTT6ZTrREQ2nRgM905lQebMlm/qpQhulPM01qJXSvIn2HjJ1bCZnVRcMOhRpDx
au6aD5uDRJbWEnblotRbl1Y2MSbg+rSf4f/zaH4D6iufXDXtvP1m6synadrDv479
cT6mPgiUtDiqZ7bs5uC+YomxXvxzt03xRzj+5b33tlYx9Fx+ZE0wbgA1u1XRddAV
oN7rUT475fMsU6fhU7Q0kXVR6D4i9yfUfi6pxl4x65pxkAtyK88JfwwPhyzr+cnV
zJpgJW9sxSIxXoBRhoaHrvFNjnK/wJjlQm2OAqnRNqmm5pAkhAPFKdMbLmlMMWUw
oPquSQ7Wcg8zBSvyO+KCCkzlnUC993u/axBuVUCC59WFsYy5tquxAqJt4cwDwfA7
0uDGtjaZ0WHtfQKZRxZ9ZlB5DI/uXeBqAXauC1WKzP1I96dwfcoyZk3Dj/L9bg2A
UEBMUP7oTOiFWx3JHd0IWuk+jlGfoqZeT8ChBFpjJ0rfpzZ35LChbOvnHWUrQYrV
6ZoMhIcVUuziFuSfgmPc9W3jB+7JIPK10Uv5Rjjs+tB4t3FbZVoijvLPiq3QSoeA
An8otcqyAognch+ZMevdT0gIQCRph057uvKHPbCpJiOHm98N6FIcPCrk0JhaJl7R
LHFFeWCfqkH7zfQuHsHuR7A7Vt99nsGEnpAGEV+qNKb4dBl6ITUgKTdsGqnAREoQ
lWDbpMe15bIyJ2tAxK0l4drDBRi0t2mdr1zosk5f5w67/cGv73geOf00ZHG50p52
UyLaWfvczPi9xPT8CPezP0OQ/SzSGPeGEZYjuA/j++Jy6gbjnwJmuFc7yxes8GO9
T3IuggDrSWILO4JFNfmqFgLvkr1h23OlSE/9kHUYYD8iamA1Szw31mzpEuq5AgBn
BMP7yE9nKvhEr9GCosmQFIxP7qYprcqZmscTKheRydonL50GdOr2Qfs7Gk4bAJ2b
lxZBHOUA0868EYkzb9m9ER/WiXysh7oftrguLoqCvlvMAlrN5HRpXMEfnuE+q+WS
nKzIskSQuxyb0osrRkYXEdj6g/9yDOY+XengE3DkKS0GPjbCQMeKwZibAau9gNC2
AoL6HTvSLnDzP6yfVIn71J0XLwp4c55pwP9AsHhdn1XLFF+QgbkKfjUOb/dnsHF1
AVg+c996WEYCRhjhoJ6bU04/aUP8R29wRDcZYA1MG5gnBWewCjOrkMkRu0hRWtFA
m9zzHg1DcAFiNn6T68mFG6p1NtgYMsMYAi8zQg8aZC7hHOvTCC3Zv/FfEqBAABaJ
Th4Jrg2d4R1/wo2OU7ZfnFvExXUkfGwW0Leo0v1q2vGRfOK0FIxD21mTpJC/K6OO
VO3zvn4/Q2NynHcEu5s0ChplMdRdF0Mf+pL8lNHQF20KDeG0N9yvqlOZvuwojfKK
wZiiLJCrO3eyE7TWjsyLYYt+ZdgAPyZnQHCWV+uA3dAyGSHrwYE6BvBO+YkmqI4d
4cfrjKJQpm3unT5sUM8vp3Y4w7jKVT0jFs+r/x2I++PFyTs+Om3vQE8ZpybWB1le
OLsLqiUsihjL0Jl4cmiVR/da3rEbmieKGzuBKCNulFv6P2bj1iHvECDiO+ZojuGr
UZ1rOmfC4zI7fIIBYIG8Qrz5dHijdjWGNinXPM4FZdJ0QnCrGkTjDpq3qbPDAKwR
6Jox9efgE8Aqq2X1IZJF2/uVVJBDquRALMIjxuYI3970ZyDj5N6rSMSUIYP2QbN8
oc9eq2JrKZcvsMUM6kSfeXRFKssrzy4+ntIOUlr9fX7TaAlvPBKMOsu90q18m3cz
hpAiK+E8EDRYuxz83zj4PEZgZikkz9EzEbKkOICIFXRl/pY8e2bbI9J1tXGCGZjq
rIiflLa5Lgg22k3OKpLMsFPAQyhFe8PadIZHcOD/VMQe7/y4l0V/aspZCYYwiJtg
TYZ8nzmoYZjEmmmvM2HisTqD+YoSAsk76ibOY2GUXzimWxm2NH3WNR6uX3VxNcXT
RF/HamMc0FiQ/dQ9QlUTFibQJa1N7MIWuQ94sYH46Q8YX+dGInBtyCpVGdxWXsv0
qmgRNx8CYlGgwKaN32eA3nPopdvUsKPCYU2Ioa/b5eicDONUy4rl2v+8HwG1dZ0P
VGWbeGIpdVVXBTd4YPwkGEXXpre99Ci8cu4VeW3j3B80pchempUJIz/Q4BvtP/1d
vt471MTRKj9NULB5qFppzRzZmxIgZxv0sW7uEVmxawwnUyXhltGF7ljXJbTg5O5s
m38nfvYUoAPWGMwyoCOtMAWSsf3lf3y5hyitrODDS0bd1IwBYz0DvwWD5p3HLxgg
TX+rd5hAylZB0WvTnZtur1H/QnV3LlcHSaWFYJ0u1ghfgrOVdV/mr2Ag12ABB1Q4
0UX1+XIGKqDQ4nreP9Wb9Hpqs13s2GH+Qxp/nmUfaiN3erPMv9AUso1r9xT6SrL0
3BdPU3lqxQLMbMNylDq04wvWKIE0JKbWFTe5XB8/lnFPqZpsExtu0TmYPll9JixV
YhBkjr66xU5Hdn2fuXgEfyOlZFJ2Tmk88KzXSf2cNgNS4RkZUGy0jh4pXmYvdhO4
a4PAVA076+IRAJfljFjaKJPtlE1c2Xdl9p6CVfPk7xVvcvswd7cAez8FhFZnKIxe
Sd6XU1Y/u9S7Nw5u9HLSszpJiAXHckcu36oJaESmyNSAKak8aKMnO7xrgQpWInyr
PJ2Yp3TFIOOi+2AEaAJEqy/ixkUa8hVvn18E+KZkBNwX0ZMLaG9fZtO1a6hqZa/0
IJebugtMltSa/bY6SapAMOEPzOADFx37iizUMauksL122JpkYo45tjFYqcj2y6UN
bMClpJqdtI95BXotAvC4F1MS9Pi06VbpyW1YG7AoNfaqc9cFHChwbqArKa1qGyYN
kcwu5MOlBcgU0NLeppFipMdKtksGW7fS8lBLIIrEs2nrNczHB9O4B10Ur+qqKr9J
j3/QAK+HA8mGuGeyBnqnRDlnAJPTeZtz50h4AEQspx1iTZa1FZZlUMVYlGNrdMvR
PTzwkAQlMYRr1ys1lfoSyQKW5/VQ3qyyhKTXgpjii4xub/NCaOIBCEKJqDpajloi
peDz4QypQGrVbtNU1y6bBB7gJKqWusaw0csjcE+E6bsXgykYRJEGP2ym7F5yJUd7
itxriuHWa80DT/NdigI3BXY5v2E7WqDKB7b3i8tUoyFxnqBTib2RjwuA+cY8GhBa
7ailncy7/xn1VDo3wv+6iV7L6hiaOyb/jX7wtBROQqaIm8jiDtgRWtoUqAfaufWH
56ClUbO+8pw3OkrhkcuOu21foPuWPUGi///Z5w14BjqhElJZwe8pMpl0zUrrmbP+
8X1QS/m9ggcUBw66MJL1kbWU3klR04ISUB46Ce6Ohv8HNsf3RfFg3rVm8HZUQ+7D
27Q8UWRhSwZ+Kub+cDp1MHvLl2JU5922KGwEAbiQGNj+wduZAHaMsCWwPnZKAGXL
Jv/aA4lPc9FH0hNYGv3d5WQfPv7u29gK7sjzUzSJuwxBnMPYl7a9C93ICAaLeShw
mtW2Rvg47sw8m9r0y/HdivNmhW95De5uvzZPpm7CcgrR4vWLk4v4wdGAoV5AXe6c
h6nwswi2gVmOR2MZl0PpUYudDSQVBWuDVPpf8y/AWImsnH1cZjgYfMiViR4jfKYO
bQZ1te085gpEqN+G+ZuhTQ1FNkuTgqVsMuK+e2Lik1kVAsAgY5aMOgesvvSdoFxh
WxCY57r54rxV6AqN6HK/YxFQR3wT9dKGQUNCxtC6jMGKgnWmGp2nNg/UqJZbyFjX
PXOu3FOOH65te0lVv8gEdDzKSSIk/+UCVD7W54xhqBvWU0zzXD9/UYVh+idEzinM
qCS7Lc8+d2rGzohMN/yVppTmmGd1+v28WXCFSVPkmn5ZWOmMDamyj/yQ3xrZtobq
6zpq90kWZWcu4kVca6zEPA2aR9C1oK+pMLxHqsaXQOn6ijJuioVxRdYUAOGVkZ+B
H0RqK6T02GHxech+4+IFr/6Joq8W8gOO/eUgBpHxb18dubM80EXN54qQumo0y3ay
iBd7I7YbsWwgqu+uJ/B88NJGeFTLVK5KcBjfYJbFTx/B9ez9Mt/KU0upTdRrkGWb
gWR3WPftwFUN+Lpg3GPciUwxxxlCFCrmsRp5N0d3kuSS5cyKDmqn53LzV3YWclGk
jFaGcrfRKB1API/YQ7h93Y1IAppMd33o04KwE5sEceCOn3NPcwQv+0tJZZ8aLw0l
ColICwzkosk/mzGnF5jH/qcTjrNn6hIZAY4ImQjR8nsVrvE54IV9nZkAeVzlzWxj
GVkv1Z3BAipNP/NI8+nh+x4p4+0U6ZXmvmFBrdxNSy7znpLrP3bRGXNJM+S/+SEr
zf5tH+13wi/ah03WwkBsp1d1Z8rWWGrSWvFv0zRe3L3DfuH6Vprvz5ML68oI1iTd
XqYUmZwl+I5G2oMfjkArOSqP0fUZaxgs+5Klc4aQwq27f4+Nas+ZLNPxzkhzuiM1
Lcid9V8h3t9AJ9yVRz2HJtzz8u0Qe9JXWNnTswEmNd61hnmRWLcKp+xgAoMYmvno
Rn0VXYj1GgmZc3bQZwYZEZ83+kJU/a9+yM2uiLMP3dWe2eda7wcC9aBZ6KbtKJ+W
dhOUTuikM5/B7rLyMP/tktcVkA/PfyozEYdBtef+GEjHBw4bcP8mIV7vuRgD6DlI
5LDE6Rodj22BKhCAK8RbD6kRvlIUZVt361pr/vftqmxhoLw87ZjJXaHNjL+Evvk0
ckG2oT8gyK3+OUInbP6anWwMde59AYNIhiLPen1pZrBJghN0a9HzkGsZyr0+2JIS
AsAgZhpu4IYM7z29ECxHe6v2Ea0jnTCO2LlcudGuMFBFQdA6YG/81GNdeJxetXv8
6xur5JHam0+VKCxz72uhO4fPrBMTe1V3mDX1cqFlEyqV6/GKZvl+Wdj9wKClKZ4f
N93JWKb3qLdGwIKHJmEcWV1y7ZFWFXDPrt1btdhW4tvI/39N1XJgJ+0GQ1LykMx3
t8aNtzHazDK/dqOL16qNPkGEGwkt6PsoEfI9HOEPq5CLoHUdHKggUGxOprgf6U9z
RJjjvUdZoX4XkqcV9DOnqliEo7lowKeiuE1z7TdM9tQHdzNH2oISrKJt46Ud+iQY
y0t+7LC+ePWLNSRBfgvH9ny+1posVzhIJ/H72tlpQG6ffKE8GZTQiKQhFecVHZR5
cG487P+aWoNZCmU+8k04xlVCA0w/BgIBfVSFD2CayCR+j30HHQVyiejLrEW48PHX
DeDY+zLj5EqpwOKSWALgk8cnVaUPxz0SbxKKM9gmn/DsfkgTbSB0T/Y3hstMD9gI
rDZyAX3Njyl8KZehZGVbtzVBUKvEWf292vh9WV556I7SM+io+63xEzL6nrR01mP8
xwBo9TGQm8zs5MrffIdb+p0Llu6UXbUXKRMWxak6q7UxRAcI/1bwZWIW2K0N/+T1
KztTZkn/PP/QZ+7XEi+3e/CWYBHLLT/QZJlTqQMxO2pXzt3cvFta0sMNjr9bOCeZ
w33hdXXAzHRnW8ori1S+fo72KsZScnCByNDldN4qu5V9gQu3iEBs1rG03TH0RObu
78KCFzDtuS+LJXErFXckW2/YRADfmVoIloWIABDWJA3os982piZWNXxqWCECtvAO
fS47y6uQBLyS1wQOPxSDDDcBtliBKHai4MCLwjQmRx9/HSKBjkXM6C7Cv+wInAbD
P6S7Y9DUvWu87kTaywiHBiStZgEX1SgGEqaAmYTro/2p1KbW/K3QUdA/Klw6f1s2
pp4HrVG2ETqoutBp1jD12pr16UEg6bwajEBWx4OrWqQj/Q9bh/NVIgVc1j2qWJiB
boJwWRpvLw/iCWGtmOtVdJpp7VYwhx1/1b8L8Vw3l+zg/u6JXiV6MKoYmnUJh2QH
d2ye6KiZB4/d98pRZZKWnBXNGphc6EhF+7difi2C9FotLxZP9lLeHarpKCNDzEYn
ubQaHB9DjddnFwSOtMhq+elU/4irTPiGZlCOUiy104fYFTraDEDhBJtm5qgwI9j5
GaVPHmyQYaNO4S+6RKg87l+A3dd6kBo3bVZzFiBneAOyN04FjO29VYq/MXF/zuoP
w8uD66xQeOL0q6AIqaV+ze72PFrDELbgXQuPQYJ5wqWaSyXpHOhjC1ERQCFJ09Pp
1BZ4sFyX3iXc0AVNvRd7Uau/PDOTKQrLW3WVwqpSFbfJKCtu1R9QkUUlXSPs22si
6FTXyxnSjJF2salNFw/QC8FdczbXbfv3KRvNLFTE1Oy3GZb5W7LkK0aBKKV7l2aR
Dn6k4RLDbn4HUplXeDJsFJA2MINTb6G88QSQEMpXJyXnV4cwQrIFNY5xt4NNacwb
pNsGGMJn9hHMAlcsl3j4KzgT5JoHmQ8qT9J1acy1X6TskmKZy+a++EQVL/1mKUhz
JkfgOrlG5WV5yGeGYmaSnKoAjouDENg+bJAAt4bBW2ibZzUsaPynI2N5RfD1xBWG
kiCzIsnu81kobhpIUw9BvS08nOhe59S+eBEj6P+uPnNFVxoR/Dh9BK9zqYA1LOIh
2uRj+O8ryxNoq0GwdIcPSuwyfkMsM7+S7rOTT4SGxZnGIHzxGxE6EjBZDWjV4YRO
WB/EfkAU5hmnecHX3XqJ/zuqrq2Gr5NZU5tMsFecI0Sf1sIjZebuQhBIjeUrOrpV
UT8yW6E9E+XNHJeI2C73VheZ5Ghl0fswfd/JYlJb2PByy7e6Fc3o92wHLs09p79C
CXvMEDSP96oLC/hHrsmR/s/DCeK4HniwtwMYq/Wc22mvtTQVOBipYneJTEoYvuq9
9sKVVli7gH2QpupY4ZWQLCffMQGEJ+A7V8TDx/JvO6s0Ugo4RDBxO8DaDHStot6j
sXzlKjDxYWkJJKFiObeCS2K4ipeP3eqTj8xshQdjiN16PQG6/Tjd3tqM4G0G1NUX
tjl6Bv0YAm4yZ07SaV6U+957IUg4Cs5KGvdjY+ZP6MYJxgXpIU6diQWuCZtiRd/y
tETH6Cx2TGxIcrasbJwuyvwqpPERFRjyWi6Rc4gDSDVo6BKso7k0En0mNG3O+bcN
0IvzlX2NMdAlChZI2dy/oqY8Eiy25D82X+HzOXz/LEy0SvJvsZ+YJkU6+uAZk2bY
WVGkqrtskzox23mplw4JMIXz6yPPpRFrPtN2VN27L+WGqwKkx7YURFxs82mJjNRF
8XJV2q7QRUjxUKatsj8T0fHXU7gCj3VhJEUpCCk+uge5KcIsObf8jxdc0j0t6uGa
Pp/3C4g0Pvj3wzH4w/5KklfC327iuImW2IhXTVz6zfdTxZANvtVBYEHfFGXv0OYO
D6jO4Rt0KBX4mjHdwc1dGdEVfpM/2xv8J2Mvwuhn8vH8KlnXsr5f6OSOGrjaa/qE
I40kyIS9LUHc2Lln/Ok3nbtyoNP+nwFmG4n+oawhdGNUr5HtG6ULmpPlICZVHzMk
jhsTlwTdSv4aZ1To1G1Pmq2cHdluRkdaJgd8qJk880Jw+JbCK9IAARhE7pnAp2kL
luGO7wrIKGCopwnG1eLU7adbABlhoc1bpLK82Px59C1bBXOKzk0cWOWfzP1IgZL5
QVOW+K50tssBPBJhEmVg40D6D+B0BL8AhWljjbVcPEwld79WXlDK/xQbKQMN7a58
iagUn8l9oSqqbEOxY3DTUhoF4wwfUz611B+GjZnuRZmNN5qtE1C6Q9xbZcUho+IZ
paWmo1eOwm4jaxS6+U7ptK0BylL2FSmPmfWe70I+l7O3eMFR1N7NgGg/7os9zeZc
YsnrJNXAklZSudU20oB6qEo1udEPvGReNCb7k5ZGVYUI2ZDxr2+74GhURTjodB8v
GPrbAvpFenMkRsg2jebxvhHMoFeVpI0+PrgIBjgUvwFXj5ByHt2SOEJpQErMAEwX
3i3pDq22pIjirnSWgQh8NkrhUnpIG3HZ+sVwDBTS8wgsyLSx7n9GyBTDYVQwUdPy
7pUTPRgxFUzmJBDbyHn9PuXtYWBmBI6CPIPrDlL9ZJRc76sOT2Kq/Xm0nyTBQof0
mWDC3AjVpqx5DtfFw9zguE32K6mk2IM4i5Iz28xudNBGZxMLGizvRhM35glhBABe
vIoK5JV4x1yDOvMFMr+oM83ZfMvO24f2J6VPxsy+DpbsPZXDY4oTZeUP21E1eCfl
BkVKB3D+YNlXWBhiRp1Tc1WpsICYUgsbu5NtTd5uwSHli1kC49WYFRYRvOVQ9YpS
94wLAHycotHK8DXo1jtFsmgYxhqiAYGguFTrikqvVF9spdZfy6Rkp4z4hu83qoFJ
qsqb6G0fYVaYXcb6PRMyKzNo0rg6Rxi6ivpDbT3jnOqzp+E3X7lAoq48Phmh4vTl
MthKR+yaHITI4B3qUAf5TuTDB5YEGZpFhpphReuyD0JRDodisEu2IOmnuGbu8jaf
X50wX9tElJ/r+/WdCM5KMN7tpyLPO9MUHBEjEQ6dk2v2lA0wsfRUu5cq+R4FXw9S
jnfE9KJPDL0dPfDHhf4XFL9jbwwZYidYFeTC2NHNGhBpTiX5y8RRte63kUkKdKwF
pxgERW3alhIjuRisW/317xPbLdBPiVTTEdsgL3U7EMQd7M5PUnLWRHU804DqZSJM
sCRdd292zE4sBG9w1qwdY+O6K+2H8FCIPvWF9hZeSillnkpPWzWMUhbzjsaohO2d
33mEwS3qAeEZ+8elTGU0MfootCI91ME9zMi+o3HpQW65N2S+9XawEmInyO0w8ai2
aa8/nD3Sx4lF+U2+iDLLeECvEZWmNFbrV3iChBVFkSgYdcekCso6jiQVPmpSV1XR
gSo/y14HLg0rzdLUqSOQ8qOaIDUgP+u/Yu0wRpv9QRFrm+PhQXop39DC9wJzWY6i
n1yYavf6VOgkF5hiUjE8S1mCnG30ivTGnhUrlgCBe04d3WhHnHLSRglBEpxCyeXo
7F8xbTODXJ+LlH8+qm0K5ry7wt/IryEOK9t47P0qfDT9Y5A45Y0Y4NSitGov5GYr
qDFHMOjM9vN7fiZgVuYt2AuZgMKY4QI5GUyx2C+Rc4WJYmKXglgJ0dx26EUjLoTA
p/UQUHYCxjccJfHZ0pR3CH8JQdkwNKnKgYYHmdLA0Zyp63vpoxQ0aPfrUTeQGmVg
LKliuanoJLygANrsKQrE1LaR7vJmDVoP9nPKdYFTT8Cu8yzAO6pmXq51bnM48bpt
okgXaPdwsFPSsOOTOM7ghSa4VOuqG29N3J4LfSqJRd4jvobgT2vPKRGe6RRDKCh5
hoqnYfdP68eDWLCVH7sh0UOSXLBwSizyzBjpmJwopKw+Kkbd3hXX0rKaJDziIDrj
XKoPakBbAYkXF1cqHCZW3cycwO3AmZuKtO1cmsiYYG3iZmxoMAj3lj2tSjLDYVHK
XSrleRjBtXPBHDUjzHluyll6BYepyx/V1c1Lh0Jw56XO85ZvgygNuslyOPgwX0aT
ZYXR4xg5G8xcPoNXILVINKr0nSBDAovFuz7asKS1pnLxyjrw8MmJVggBR4kAx6v+
QgSdS8om+PAxzu7k6x8C6UF6gqu03Wjlp4Ga5ZyKoX5c+xaxVq48jcNznqbiSVQz
SUuFA/FbmNxAvSzUtyWxUnpLlTxh+99P+eaGhmRMzRodKqhOiB8r7moACL3F7y1/
WnH846iO1GtXOOQqf1XKDWl8J/zWOrws1In1PoIgQKMq+cdNntpxKI3b6oseaY4s
cl3j4oHdxFtwWj987IZC5pJJ/c/tmrhQJyF2K52fLzbSLCf2uukSc3dZjyNPhK8T
b6f+duO69gaJ2+NU3xHhVhbKamCLYyjMHiSznnRYimUgq9NHBhpS00A3a/BCkK3a
2/O2XaTPnNBqU9HWRMpGxlDb4NKH859oXl3hCLhddIwYARGNUG6+WEbni3AQZIe9
Qxa90ObPGC6ho3Ul+InfedLDN0zfXYN04Bxj6Sslgf9jNNHBPBnwQOnOAWyZjp2o
0+J476PyCDZrj1iyFcyx19hjfe7qXq56nGem9JOpyF/NFMsK9QFgLL+/CJ+p7eeA
0fUCusiugVlROUovfMIAowKcSYt/OmP/g6oR33EaVCiu0aIB8lvGC2WnYJAdpLhc
K/6FkZF4hjan6GwIu1MS0wfv4c4GR7BnSKTyhB1Ol7/lbiqPWJK9CKqmRIMfGUwL
T6xhjaJzCgSZ+JgXAoeWW2lGg+oassZMMWtkogbNGUwkVrkjUrTL04TZasHva8g4
VJKLypRKk60yct57NT1HnOINCNFAwaYCe1nAci9Uvcq43eEg3u3jpPXbcaRiu6gO
5FKC7bHZfRN7hjmNhbCtcrK9ru0AYVC3hd9q93z9UpfeQmxVQGk0nZ1u1H1lYQwd
X49Py0iIWO6amxvC7ptgyamjOnTkNotJBwNLd0htqaKcUwxyo2Qp6nrNxIhDH/Ye
k2SGIP2SXuoCOTTVILIdVFMOL3KFgup8eqm5bryOu0x3wbvBt2YDfKJ82TMcA34h
COru1VOgwWYheArnWFGCE7AsDR8a5qA/0AypcMJT4j4Hi4MVp9Mr/qUiXpqmblrG
ARu6zdJyiH1RHFcW3DoBwN6kNeDKl4gt3GyLv1TcK2cTAmz+uAcRsOCl3Zl/B1HE
SW1NL/57Zw3C4Z1U0dKNnxAqh6FUrO63k8c6we/8Xv0vdrnB0om9tzFje4A+RQNm
SBFikMFyEHImjHkMRTZuUWD7uFNMY3tfXtOgid4M29fmgPjRusanuJIfFiEWyh4K
voJUukeIVJ9g3nN9yGCCycxkjT7ejyQzHW7YlZoycZJ3JOENlHYhGFwzRDSaMa/8
ZVMXf9hdP6V+Kk5o19nAH4MW2+NgKsWtDldKYUK2G7tyq/wp+z+ei4xAnARuFZjQ
f9SDXcFUq6jQKXQcaDcdGtD3Xb9ua7nIMYgHmB2TJDVsJdDw/kpdX/nSyjr7X2w2
AetI7jzN1iMlL1GG8eJhp+WykeAXhoHY5arNVdmnb+uxktO+oUfeq/J1bbe+R8X4
j2Y0rDCQKpsxf5037f5GsVT8+eKySO9ZTjkm5v14zkrAPKWeDebP5hQuaeMWkm2f
Kmx+MUwhElRGXSQAIPteNKjwW2BSYpJJJkYrfl6CReIMWQQqYNalIUMbydu4PDze
qfOZuc5t41vOcBk1V73f6CG6YG1f5/zXqgEUSXySGo4Tu7g0jAoEWXQhm1y4/XD9
UZz16r+AZg3G/uMofakci9Fuox82RClFqbFLYOLJlnsVrGQb0K/+u0ZwXzAPupkg
LxBpr7sm2kKdIQf4cwxR2CUuMqJ6FhrOTxJqOj0LMVr7TGDjkQuAOvoAX+Sk6k8M
RP7LiYC+zlg9Ba7OwX1Qn7T6u8jNz7ToVQgW3pJolkDwws0IYJXbLLo37UWYONIi
crPMhk/FNOHsFqgAG0Y8Ppvv6TVhHhd9ZHtN2e0kQnpMfy4H8YSH0kBB7uXA4egH
2tdSd9xXT2qMXzKWop5SuRmrCKxZ46nKG3ZCEuHPBL8jwFKUqhPm6fG6MO5bkHLu
CYpczZQJwoy8OjYHcrAWRvi7FlxMZIUiJmtv8WUcvLyV1iqovJiRvVHdvsaDr9JB
74CINPA8O6aLOZGGEM/3mKZfbePDCr7cA549uW03BTlZj/qCEzVuCjwT6meEcVyW
gjJT+6pJde+O8Euq7XKYiTI7Z21lJU9J121xGLJsbG9SSOvOnFJ/XCw/Xy2qMkDX
IA8DDLYYVPuCQqF+Gp9Zu9CmwHKrSZRMyWCV1zD3qPL8o64Kt+nnCCb7J0A6Rimv
0do2VhzAzvKGwCGJYTVRfDBeeZiAuo6g709GfGvtQ67nouG+Nf7Awf4xXP0S/VQx
jozb59o5paJYL9WHjxjirVMW41tEC+dzhXONjoDRkZto76hmgRmdGvuxX5HqpZU+
gfoKClin873nH8uXt1AGCLM+L7q6qcpCs5LZG4SYzIeagQvEhrJfmffBgGu1cORi
jZSPCE/IoBP32y9GBb04yU9oC7qET6+I0/Ksj3xHMxBxdsHYwC91w6BZA4JZ0f5x
Qi8GM7BnhPpxNuLqJ/gaxUOg6NVg5CgZi1r2DUMtOvb/EuBe8aWd93MVj/geBj5E
lfyAHuZF75GpeMl8N498mYfaII0vGdxpDBnktGssWyuzBWDbKAhUbzJZPwG67w1v
8e7tmFnVLR/5Q7qTea/PNTTkHZ9tyXsx6W7ORIMLVXfReRox59yFcVc9n0Tpo9me
SDx1pNMHxX+nyLLFGwfM642h0cEbkyf9b17wPCV/rOTVMCAw6buzhPXt/r8XGNsd
aGQ/iFqAJ56H6TTn/w/rpnYlMosW1CabkLMAe/sdStkFzgiJK37jGHW9I/33RKIg
fTQoo9h9rbPqV2RBgPUW6O1WZlwTFyjpapA2wjkB3xd+a2TDkscqMLDAQZAheCK4
8CwfImWJW7zabdDdgfrqGXoi6204TaH+ZjimfrX58HmZjjzoMiFxlWNUPeZmrbyC
nmjUwwKS9C+qVz4OWhOYdNxgWk1nLQVYkCsAHOPWMzBSUAgdb1eM/dXVQORlU7dZ
gAxpaSfR8r6RMEjeV+jvi04HUaqerhcauJYuNbsrVTNPmGEZqsxwulQWxHS0udvQ
xxYTp8vSri62VcStnmAC96uwuhfMdt0u1bmAOZlEva17ZJDRKRuf2QVz3drt/1JQ
z1S1X1WP9rPvku8bkMJv2eOuDWNWGyhXgH4k6JuGn1l03Xfxwuf3tcLv1CFRynsC
zIPYNrMcn2/4BFB5X9j2yJHdOHuWHPmk6DedXLRakOczwDVCX4pohZ+xuRWooCkM
DQDjkDKiEGu2882n/xGH9ZhDUhLNPD9H9xTicQbRGhtn0LEZM/bnaiazIme3eDQP
jKN4SuESxv4pOxVKm6sn1mXiKBklqe+ZvnwpmZQkSxG7SH21jZRUghwuHYPYApdO
ACUrkd44PIs4rpg220E7ocNPjvhzjcWZ5fBFHdW0aYFoof8FXMeXhDR5gHo5gSH9
h35BIoZJY0tLGxlVS+co1o/OhTDNuYNSLy3vgmFa3rQlPCbTHIGkc8BWTTiNZWns
QFrIxOHrC2NB84OfxhtHL+CaR3gVWIyRHCEpFEnnn/Vzysw0TeYCLdMzeQ/xRdoC
Ur2GabNRQLz87pQEno58mfJvdawiAqEAB7yDP7yAq8KdQj6trC75NcR+Hb2mV+Gd
QtC2ST5w92gZOsNwtkk4kjto14YFAQyZTX3ENOsdi5sOwHEFVnPCr0vTa2BzSipg
HaC27ufYou6oMS/8UEHGTTHxZ5lyupOcPLz3jgEB9YzsKdQLE2rJG0nL86SGg1Fe
inwMh2RsIJc31yrdcIYvhR9lusUt1dXqAiAbw2sa8HerV67oJvh9/PP3dqHgRoe8
mIgn2UBGcqCsHKKZ/8g3R+SRSpILV0xi9GMSdfHQ97u0hUeSD40+7rPRpnjeN55R
tuKly8gbu3H3fcpEsnJpKlf+j/VWZKGbNphzGTWTdX3WoLWUkRkzVzOG/bUscqF0
bEca/kC6wU3XkEsbS4H6w4FBczGDYO5y/Bm9lDOSyaU29G0NY1KcvL566uMf3rEl
h2s+VZd1U1+5TruEY3ahTQbmEm5RbXs4GzEQVIL2KqxxRRr3U5+OF8Fl9LKlwxZT
XYvg5jTU77dZx/KtSU3uIIb6Cyd+eY/PoetJZv1SmbUhiXAkSbH/kp8hrjLjbGgG
N0AKOw4VcoyRR/ZdSiPlb1K3pX2hSR30MJ82Gd2j4Rm14F4hPodSdgVy9O6Ut6Bi
0TbKQjPs/35tH00k9r3K3b+2Y0095giePgHrDz8qGEJf2KLAf0LYNE6QlYDtBKZP
MSWhb5DUoDfpllss3mUAqVOS9AViRkr5YJkZcKVM5N3YXKU+h4ZgstLMkVAPD0RE
lnN+ougYOwjA0RmYt5/VGhj9jcL4sNqJKUYrCqfvMuhBBcqkybnKGQAmSjg6Vv93
Dmqkd+rceu61bhTljlNLmu60kC2sf+jTpbUbDwNSSloGnvdVyhqosM103kqS4IEF
gBuUAAkK4IRO71FZyqQr16IZqJjsbIlbovZOv9KE5kz1dL19TjuJxwRamYLOLpZo
5IKG6srEu1mAb3N2JPMfkpb9sJh6wHBVpVOhsXR4IgUi9M3NXx7SeRzHjciqlO3u
lbyJ+RuXgmIKyP1zaGU+0W8vv91F39ePV30TWE036VF3iz0m3A0p+qeE8NC1HUxV
EPnPGle6BVcldyvChAZRVylrvZJAKWUtYgvtRr5ki2bStauxuf145xE7WtOVl7hX
xS+IbixoJPG3yucyGJ6xziyejUUkKywoBsAbvkl0x0UIlurNfucbv/+kOWkb/M+Y
Y+5fjYpryrUyG3QIRp9eLlRgkP8T2zG2rund2tLxMTyHs5eqzQJBtluZhMIXTBqd
zy7sniFcBJvIjPzOzHwhe5jypunT1mgmJ9xOeA/x4zKZ92uM/HLt1QnvlBvGs8XG
QLwC57cCzwKaMAqBXiALH8JNvCCGzaEJhJ0sgn9gDB4p5/Z8gHVqLbXKmPwh67nD
+qZ4CDTMK37431mI/BF/9Q4bf6CXdPulxsFM21M4s1Mvy7iYjbiWcqUVElNcPB9E
tgScm/H39560SwrKRaUwSDE6m/rze2uv+fERKesXVeL195q9kWkSKqLvPl6Y9HoV
xEV4a+C+/J7gEJVZYZFUqIMQVB6nHPbv9251XmQE1kr/4v0FogD1OPHPR0klmqj8
O7+Zj9onP32XT1SnQamoNkmDohuzBGz9oSrpgvCe5gevEfzlyl0DqxrJvzaQNXYx
o4X1o0B66RiOIHAYZAFLs1kcWGRmWC5R/nPLx7mgkIdfILAdHrj4DPSf+wZyZPyG
22XqkdZjQ0osa45Hk/1NNhrUpPOFcClFrQYzTrhI1G6hAPSc8NkvQJJfBgCWg9Zb
ivIlAqfBjY+hMqxzAEIOvdM0Tz+MXV/eRA2hUS0PfEO35sYa9WKkcZzEX8jG6dHS
xSu60iJIxfq84rMWN7EafMJju7ucZHhFrMXKRSha75ZY/hXPTIIIqkRnbJnpTRQu
jiXIyC4rY2urPQrENzsFDEm/3fu/UYO9ZWEjq0ULoT1ABFnqdOdnRUYTsbSFQQ7N
azwOJll5oIpDlMbxX6iPsOS/QGBq0R6SjGWErAJNyjQtf0i9EqcO49m0CsWQbgQ+
8m+8VM1igQRQHUGhKRU2DrJcKdwsIuATjHdAbdm8sD3O7VR/wDlQPVKX3OlY+taF
iu3gzHNVT64+V3SQRO2DpJDAE8uph3ZFvB+rPoNxW0FxTvXqGL0Yl9HvihHnSIW2
mrPHyLS6QLg2xBefVCsvZYelOggLqFQtYYN63uUWCOHRU8uuUF7wXT3s9LC7w4ec
VHM0htG9RLa5DqFNl3NX0gVH8xuzLDW9F2kgBGoR9LQ5iq4n7VHfW2wY02iqlg+t
yGnSnA7wtRqmkdtwNujUfiHishfESaywEF40FLb2VSR1v1Rft6Phz0X9ll0Kusyf
rSMBUvcK5IC0vZz4M5maJ800X4ycQihwJFcnyLxo0AKaqNq5YlEo+HmW/nRfWLsR
A6wmfwJxy8ZKi/VUSxquyyc2vbFF+jpvBOp5Yd/XfAmbejzl7QzDSkC+BAVOB1H0
hougC0+sF4acxkISPe0CF8SRa89Zk2ZSn2RBWUXqqito2u0zBSoRfgWeYQMFJ6Wd
cpW/R1RQMm5R5uSXzA6PCDLoWSyPQS6pKuT9nfI/09rS9XraYXveBUH9eZFhvjb0
0B0/RM6OltYbCetdTZWDdLlfoyVTA6tQlU//aM7MAtQ/aFewy/rUmLI0/CkdeQpX
sh8+5yM5p6ltWIF2XB4EU59m1YO6oAsccPpN60jLTqifMHpNi1C1GaKvEw30bQ/3
Dgi/c/eu1YJ8/xXRv/clylLjeLrjbZDPnoWyBRDdeKWevb7RhXV5dTQifZ9Q/JU1
L7Eef1MmHE+1m+OR9xUv9e+YKNEzEv7NFsCclt5cQk2Mwz2M4lY2geS2a5V5POot
Zwv3OHCXLrm1Zo82dMa/C0vLlx91m1pAML7J7vQeL1KIqXjb9aEOSZ6/n89eVeYU
yeOkyuuIYUc5wcgSSKmrMZWt5be5uf7oi40o0POV3ETdbmWm7Inw8XMp4IsFG/Wc
8BzGyt02pMscH1ZFfA75gUVf2cfmmioO2p/OzdEab179Umc807KiH702UHEm3tA5
tOu2Rbc0U0P7RbiBayo4hc8arsQJ0DPs+j+15jgosCYs+8QlcxlZy01KbfX3+5UJ
wfo0mRDMm22dEiGiGEK1KLqmh6j9bqCr5GUkdE80v47d53fFeV3ZK6i3uQpt930t
RnN3jhD8EUQyl2f00BtYJ5sKi+8dnK6pZs2Nnv4b3qEnDz70pyShgPsAef0biSrf
L1ubm+R/GVmqyvUORUq4oaauJ+pGe3k8VQ+3LL3L2ZYP6v1IyPqayNvi5wNalYms
GfkMsSL9mbTDI8V7Nb4QhF1vWq81k9KFGB9XfbYPPvCt7f2AMy3yHvWoQ6NVh0bo
EHjMbnWV09FNFwkJE36SqmHHWfLZHIF5U1X0Md8AvODQ+o6tDTrVtKDFx9ZY6AW9
uP4fhtnz92zSm/rQuqLoo4K2AQEdeIHAaGFTgO3PuY7VXp0SBuC6PoCM16gXDHvR
bDI/HhuqTXT8EgAb5MO7nsq7u8toZs3qiwGt37G7oTBU3ehfNDedvijiQ+qNpIXx
Tpd6QJ/G/OnDICeSbyGEF6PdIs+5DOR3G6FLOGK4EAylCj4UK6ZnQ7cSN7oezg4l
2tHKq9q+IVa7P+1ZINlemvwBRqe64+pM4149tIk6LtM1b/e9IshYHzd66GTDy3GW
wVa8bbP4CmPM43fttvBNGzOYSaVqlFVUMjE/PLd/8D5Haj4nn9fze0GJ/sAInll4
fOBHS2dpBqpzGZwMB+r9WChvK8G5Mg56+miecJnP/10G2/gHy0aUXUOjf4ptpGio
NpRWXpd2Yt8lhH7aBAuR1tkjmGEONstWZV6fXS7ODc/S3zqldYfYlEZaA7NMUnWn
xp8fwMLt/Z2XU/y+fbr5i3qOrQ1UHc2mu+mhUASL4f8Q17uSo6tmVtG5G84q154U
RYA3KnTnQ45s1jJi3UqVh2cAGKe3e4QjdA/Hg55InHrrShbLEgnRSx6yPrs+gmUt
zm4imxp6pMavd9vIF70RI3mGCLQXOyC8a6tcT0uN+XDwX+fpheYVujz8hkFMxrc+
8t57W8Ubm7dOqccy6tNnMJF6RcvVDo4cdJqtGiSsbCAHmEXV+0zl5DNhNgeHuMku
RCaoAJWChasHp+wXmt5flggnKk0jigW8Ufr3UurnLZZXwc5XG1F8zQpEZREoZ9jy
f9/fgOV1WxYO1VCHZ6xjivvKkevY48ffsQqTvuTRUnnR+9g8OrM/0vTWCSVn27Iv
jgB3KEMfaLoTPrtdutul9rC0juN9xho+nsH8C3eYEZFQ+62wWJtUqhGgN5Kgx3i8
oEUnvIEX6MlcHwcYoWlW9+78cgVG+Av7DE6n2coENE8LezCX8JepevU6eguGKCTy
NbjT9ZJgC7HHB3ewvqZGQjeKwouZdxhXt8yldVmddf+e8kAZ687q8xENsh2Pe+WD
u+JIMzteNiUKktUnRxRybwy41Zk3Ub9U8IK6eiLXmvi7L84D46/O4TEICQgOxXiS
6e5wjhtqVUwSDsrZFrULstGVjXOJ9ogg5RupeqWeAm2PsNdROti3q52Ln7L4ehm5
B2WMPO1tHnERDstDUX1Wb6ld4mlGCsaei5iNH3c/t4GmQtaBsQ3SxXIWmhaYs12W
7z4uwPkOUQDYaqGzFIl+Ycm2bjAMmr/OYY6RT3O2E1Ee0M/isq/po9NhGueAX05y
ofidcXGPW41IZa5qCGv86zHNJIcsGb0a3cbO5+O7irGN3NbFagF37ibZBXbD3kwq
d1VXOjxCX/C6zBvrHE0RufTHlr97nqxcUQQHokDfYXAL3d81Xp0w1eCH3giSksPd
6m1IaHxG4dvOVWa5tkR1dZFcQku90zaXCCCcsLFPz9xOumPdv4mbEFpXinAlphIl
sbon8W9g4sbn5J9Q2VH6xj7NCcjgygRU45FUUrjzq486hNuLrMdXzGmIThqa/LOC
GGzsPDHt3jGTDJr1pSPObI0Xr1Q9P8MPEbsZfB2D/UXfGwCOm1y99X41Lmd9ahE0
nX8mLiM7+aGFv2JiFKgMeBEl/h+TrZaTyLowAALZZV8cEV9NCB0xqxivzyePbMfw
iilKozTHcywnspiYWmY5IXgrN3cZIivXB4fL36O/KiFqpTnJgDii0DFwkyN+BqEA
bF1qVWUdoRqct2T7xuXrvawWlKYsnNUTmoT6fIcWmPKZQNZvQRGuZCVvJ+iGgWTO
9ar2mmkwhqgLYj89EucaffBj5Qp5yukRzvRys/QlBx6a4dlelKLPM0Fsls1rmUMY
sCEKO8jce93v6SVP7OZgQQV9zLS1dw7xGkQ6qycJ+zmbT18V9yQ9WyXXKGECwuux
4CvF/5ai2+nFZK3H+SO8YfW/0JQjXSXEGuyjtbaT34iEawv+R/VdZ1MfdOCZuTFu
xze9MbvtXgIueRdzQ6xmPNHh1r7GbbqwZL3lbNoC2h2rbArvZe3MdiHOHRLhBOF6
zD+BfFnY+4Z6cL+i1TI/WsWWjVDqEnj3DNR44e2APXI/ja4ssi+l7bZUm1QzBcVC
5kFp/An8q1u7hyA5NDjTd1ph6J3lCMblES1tKf+g5YWhw8mT5WHVbV70Q38i4mx1
hH+q+VGyeCoibO4vEOEEUxCGVFrFpipt07Nk2H7SsJb3ku3OpHKgFMog1cBQhiDo
W2ZBkEIueaBfWc+LHgQd2cG5FaEAyVKtIBGv8NVf54ZvGnSPQEmcE8In4X1/nPB/
RBEomLlo15JxBdBi+Tu/NqneXdH2tbgeH+V6pQszIBBDdU8jTyBmXRKUOel68PSo
95ZRzOif3cVCHLtaSu28cDnbsStaUAndcMAbdQBRsTsTENonNapIoFFGq3tpY4VS
M3qBFAQr5MniHCF2lQlpt6CFpuzymWPNhKfuOyhCKEG9NFfmY8L8W8HVOk16VFSi
+16OuMKKvq1r8/FrerK8Ovu5sNhtApA1E6B3IyrJhUs6cLgJQleoWUoBnqukCLhb
voe+9b7Ao6ZbxfsyDvLUs17sA8Ct29EXEX7kZmwpO/Gyq64LFpMtzXsMXL3z6g5E
PDnw7eTRNwxyKK2Sr7SqW/F5Vpx3Yh/fImZVCd9lgF4fMUWdU0U8SnBEoEHwzVos
s4J8JykIJiVeqORIzxb12+4Q4y45g8uDZiv43aKPOgQX+mmGjLJgFbfCvnzYm3+g
2w7rdJ/mQnSV6sq32FJOCHW1nqXIVUjEkuChuTXWUPucnAXL6oH0I7pLFMx1QbOR
HENBWlAWv+UNGYBJuojMbj3BgbhjEEGtRxAKEXqmTbNCKJfjEIMmqdLrfpN5XGQN
50yywSE5MO2R9/JPWAuSN7Sy1dTZ5VU4UTzKYU47gj4zIhU1enWPUhoEgJAB5o/3
T9WE7p3OYzZG5R1UDIrKh6h1uoTrWC0NxgXMklXO0/IkZN3ZdUFIAm4todj2hqG2
A3XWu1VTWoiKEFNXuaqxCHK/sNJ4EXxL0ZMb8XnCgoIKEoWt/JEfaZ3thHd3h5yl
3juSzRZGbcybtqerpj0bsC9CMMtYMNdAIG/6/QWNOJL09tysIQ9OM6prNpdJN4m8
QAKnjtiwYfZkDbiWscBU62by3ZwXtxjtABLMlFP5lkv27CwSWNIIMGAX71xOa1Hw
OxBVjOJmXtFsGP3rBkl63PrB9yUJYzh5eci7QCH7HdgqIJ8uamraglt7sN9z12j7
4EU05RvMd5Wv4Q5aN1FTnjuc+qQpcOSFx+fPVCBvS7LXzbbJZrQmPR9ZlES99uck
wvCVUSMgTyna1/7R6K+g7RLajxKEjN8Uh/lC34Vw61PlyvhTqxRmJXZqbqwK+iqG
SbEMJMTLpmRKwBg+n5UhbRd7mHlLwypuPBLuYLUbKuV/ptdM7gVzFAOGoTAH4HmG
4x16asMx9BHZCfFvaMULvD95A0nsq77ugPEJf6LRNqjDG93Gsh1DRgYSUm1XW7NC
qy5ShmOS+Mu559+c758E91npGZiz4cnKlAdmCjXwyobSi7hfegaPtGiG0/e+aDQS
t8mTE5t4fFJgLvIHO58KHiQp0Q5dcYNjQ23nC00sG4erW9F4SvuhqPeTenKN0tYw
U0WJaaSX3vHjDV2yqdtGVL3Q+enrN1LANWWT2QjHzysQkRwqFCHyzHoXwtvYFp7q
BQ6hlCHd3h73GtTHIJwJyaAG1lz9iC//iORVftlfN6rFrnkX5i0AQtCSnf2yMs4T
pPfbhSFiCep/f40bOCS2/x+wKkEFH4aIKkc9X/SL1iVmb5zsxtXxpPVzGC8gCBNi
Ca0l9ifg9j5j989qrHvfEvLaZMpz2+Tou+FfPaqTU9hdw3Wr5D0sZoQKNxxo/8Lf
RAjBLLpMQvRJ6cwjGnZHEgXa92+lLwZcjoPx+wluSHdehN5pAXza2Z8rwN+sOx8W
7wEGmvzX42+0hjO9FzYlNCu//mD42fJ8ptFbJGQaDNSoXSdDJo8WhHaIKekFp7rf
vn+zv2s32nRAlG1MneeI9kWiPRIMh457WyvQEg76mLLBjtD3LnCxtwHy9f7fLSN5
HZcUSuwQ9PrcO1DmBCZsdiKE0PeDg/cTRZ6TfVtrA38tfukunN1Ig+9b8nAA2E2Y
x9FG+QGwIhLr2VEJKS7KZ0WFbpCbpJtT5tMHDTAK35QvNzkS+V26skoQHBDGVMkS
uG81N+J/j2i+dGmkKQZ40X0UQyAwE9RVQaFeML9BQb9B3ykpP89KNsHh1IMjBpgc
VQaujl4z/326Fm364oMr411lAWd6oLk0p4GWuawQl4p9pCju5d8Jmsg9A0pvwr+v
5BwJyoNMIQh6fZTYGy9Y0+f52cJgqbxx2QrTHq7ICd3kHaJOnicHnJZQS5ldTT4n
tYCGiQ67fzl1rIx/3OKtkBQQ7rxmkzO4mw2CH0GcCvbzjnldZ29hNsHwcB9ERYK4
3qMVJ3X1BkARX15LWdWkZc+gPnWNIpIhlyFhLQv8OAn6AjtmVF9VRH4ddnIZ1dEx
XejAzxDtbMkM9UmR6uL3Nn4QWwivPTAOoDWWocvJSIQco2g4l32SavUllbrWyQAC
Wb0LMX2Ygg5tF4vtpPZDr6uR1zHV5Ye2iyKjym7012Yybf8rcMA6sUBbVjErUpYj
WDq2m6s2RTCAbAwyNdn2yfHODTSVYVOnOVJTKRamJm8fujHDwrYIb/Mxj+oOjZzl
v/7EUUzNALikY3dRiDFRQd3CHkN5WlzfULaVwn/8a8XCqG/tZNsmKTju09kusJGp
0pfv6K8GXERojRO6fXf2I9R3lPRVAkowAMMi8LCm/E+WgyMByGyv6Vyo10pjfUyq
ZHnbrirjTeBRDbKthPbZ+ErwpALZVL3JTy3ydyARVyj7UtLGjiTfpIzAPzQLevau
hBmkMhMLKc7xOUUP1aUneIJXRk8ZiBxmUO84dJOwSV0uOWifzilo7XKJvwWZNZN3
R/z1Z8RAEdWQDdd6EQJUnOE9n8e6XvuVzLiUqQhjlEbzePQcjqRMBj8CYR1efe81
WoPzU7fUek+Sq0xx8fC0CQQ6wwX+2bHrXH+2M3+xUYSydy2T4/mIqaPnO6ambade
4HSuGhAXpiZ8glpWQP19HYtweVr2zXJ9wcqhsB1uNJ5Noqvzs+u/Cx9Y84NXDKl7
JNaLIjy7Ch0cbetlGT8FEZgsMt4THFP1B2kK/tGzInyd1b9idT12N9r2bipqqzOr
33NEZOm+21ydtlWGN/OW0f2ybfVL7u767Q38YnbfIHbGHgk6S/ApjkWIuU6GgNF1
iCZVOm2GlLkRcDvIOBC+CY5OxM3xO+KhGYjDCGEPjZnxA2WdL8wcuGXBb1gnpqPz
p/bIqAHQcrTCNl+Mb/XTHCsioWR0oTlnTtW2SC/pqastXV5qrkbHrx4md5O/P6zz
cPkye6gLrmMbsKqkoqibQacg2uN0WjjoSqqvuEDpcbUamrunxmeIF3w7IauJBN6J
tochUk+GIotfRgG6Bl9okVnbQQcCWsX/T/feWz5wyUk3X7CrYizBJsz/yeEpvTpS
+oIvM5YwvcO+y9BBuhOIaVXuREu53pgaGP3ruqAS3LlemvthuVZn9VlwFZK3dYAH
2kpPEb0B4fr+8G36NiF/NQc/uLdKbxUa8kSK3S3oNzLJjC3Gk+unSC6uMNNSzKmh
caPEz2JdCZYXARTTvEQGedZcJ1rs68WvP4NxL66bF6+ksfJ/Z14nNvrKzdwNY6b3
L8i+skXGqn39WMEbrv8iTFcXaTQ1VN7KGu/5GnZx+NNwVK6YpASCMB5drMJZvZjG
c0g/yumZO6DQywDrzBKlPHKFWB+94f3TIlMB8E5u6gvfXmptWUHMkD1wd+XLBJ+e
XS4ujHZ/COUcY2zbjWwoR1idPlYFAIhPhSZrBKjiUZMlSk1VzGm37ow6OLe6kgTh
3l7wXfrjyIdO5qTttxIbENsjj/dwjYfYDyt2b5cv79j7k3KphCZIVWTJLrcHqdKf
SQIT3BN5KQYyH0+9v/IwVP64h9XNDLdfAMiVhrxFp2jibUXQKPev9/RmMsVfFRnW
qZE6KElic84rHpbwzjbePMVlDcQobX5ip42KPk+mtHA4aeyWXSOwJ/Il8ogc39xt
9Ljo89oDCohUvgZqYhizNEYgqBWMltHIxu6HLNY7u8LQUiO/TvD2HT+YlkY00OEu
B/zGbAhs4bIaOSDLs/80hJ1FPaDU6Tg/UxUbbKVhJ86vSMZMJ1kn2HquWScvmWBy
ShtU8E35hRQZcJ46NLYd8ER9y78UQDmx2pPCMGPz7YvnJjWDNNDj1QMQ+bVcXb8K
lMQTy3MIULAGsPHd4vMvtTxXsT49cS5u5WC4+D7hA+jZQDBVzTSMl4TflmOZ5Zt5
7lsVQgYALpSNGoMfjzBCyr597mYioO2jYQd6RssrRAiccJ9XDg+S8mJC2rtTrEjk
EhR0HFD0BF2SM+xgCKt42HzIsCfN+D+9Oi9pGunwr35cxqoUVMO6oAUdPWyx2zd5
2ZMk0HAfurb307P4e0kDdXBtN8wysNE/gDLtIrbU4N2NADIhOJR/U+XjQMmtiPyV
d/qvYwSC1gis2R8GxFhCw1atnAXYzINX/3zs3cOjCiLnweieos9lb93JASihNtqJ
eBalAK+Nkwdsin/ZpYTF6naJtUr5n/NTwFKXp4XI1kE6QBG1KIAthfjAG1hWFjqi
tv9PujgltcYJYZG5ZglESzB+Lgf8/f+XOTutdyyT7rClnBy2uo4vTL8V4ITmGO6f
L4rPRsAOh+GZCVrkmStfbdjZRYBcIBHs9tht7ep5EXaK/qzqzRc2ZnfE0SwQmhZf
x2nJXB3S2xcviVZ3SpwqR8OYlJin1653rZ4lNaQRqEN+l/0hHq5AjQ8EgqAEHO+e
3LhK0bRpliatadxENpvm/kj7axC+U7Wt3IMzMVIcTuEp2q8q+vui2udtLQzLdZSl
tnlLvLq8T4t80dlxNJgMmtRTucLbh2XcrJF+dJ10pEPG2noUN6UHOLJZWbmV2p+s
TDNbvntuPk+wUTAnlsD/X8s6Vv1VCCrDHscimSPywCk4W2otTgBXTCSyTkeuRnAS
xlOdMrjLyIHTuyPGlx30EVoe0GIy+MHdnQPpnfGx8E4vNSEyHz8PsbPB8GdrZ/AE
7RmqZWBmgy/BriVNRclYJnhBhRA5g2kLM7DrCw+YCZSNZSCSeFsAQLZGKlBZqQWy
Q3Bux0K73OfJnJF8Yv08P0J1Im9ync2axTupMSlYJkGheapvMI3C5VKhADPPTKxO
9lLSB0iL9FmIZs+Xi8x02cqg2Tuwbo7V3ZO/kisBOgULJdbTn12lV03lu6Xq6dvB
nHzfN174yZVXp4hKmJNZOG+ZatZBPGw+waK6ICdD62Cd4dHZSuohy2xGGATDKC3F
AXjkIX7thzHqsG/tIFmBZ2lFtSj62dYgaYt4qENnJdDzTE/y1vvvRTnI1GT62sGc
F0qHlfhuDL9SdIsZV2oNEQie2HiPYImf4gHeYjISlG7KGMqIv3MMTL4vaaFp3cUQ
SFhAPmlpdifI+fmAe2+QlYTN3dB4toS/cbVXncTtI7yMgOXjIYj/Wi+eU1WU3Azk
Za09V8kTQa2STn38SNZLyQ2Bo+cQgt7wJowTwfvk7jWXro4q8dg4A9l0KS84WLOD
OIbIcr4PTt49HyKSQPUaX4H850ayafhMSNr6ZqgPTawzxKa9ixd4XjL+d8PlXtYM
1TbSU5KN4FP7wZ/FaplNWKk6V1bUQm7OrvhoFYDkybyGeh4oaC5EQy9IX4/GOtug
GSFQZ6aAN0e2c0zFQMjM0jsYxj5Hfh9R2sEM23ElwZ4bnRYzZ+NY2+SKkTW0PgBw
4gcmmG+IRqmCZZ/ttUuiW3eYlc9q5xIIqKUPaT/cgITzrV12ldZkatmu9LSVGqJw
JP6JzULzB5X3EMRBQcUj/yjOFPSPg1NATo2VbQ4718sw/degFUOpMjJrxb95BOHl
/rsNWytpDVGMFOw/+NgpHK/V2ar+eaU9kKfBWQQ7LM4aBeRMD7GD3X9VMUZkVqbO
iKIM7co9QfircMntcc/d4Waq5c2mlR91mjuQJtnpuQOZSWWQOt1fXaMdMKlvPz3L
3nUHdnTlGWd9bepnJVr2nOAnImwoRqxtfDPhVrOWOHmZJvUsG/VdylsoXIbGiHRf
Yhq4ORmWjinoB4C2svuv/vLAyRSXlieOxhqz4FxkzZ2SWqs3xxT/cxhk/1IQ9jZo
INWPeGRmATgmq1NB/7Cv9OGcDt243O6BxZg5huQ0kBwIopjlx6iwu3jGwLkkXeY9
jVdDHD6fTiKvlEivVuWNM8F6YEtYCh297IH1V2WeKkIVytCV4tHrI0lnfZJA0zdc
G0mS+kfOX7WkYuPnJxjOA1f6N/ubyWEQ0lGnpy092Ot/UksCZkm5nytiHRecsEMO
fVgDuXKSO8CfO+tzN2L6D9oKEhvCZvN4aSbKb8sQp3oq8A+zH0UBH53wXnrVXiAJ
AFj/KXSxsRGCdDRXK+UH53V/TycD14SqS+hCPFTnj9KLU6+4QXuoOLrlnUxOWQpX
9lZrYepsCCF8GKp4k7z/TXuj4z9/IWBdOeAkQjk3indEAYx+mq/WV1qfwD2/9w46
GhxVMoueA37qQVpLD2nQcjs2+SkYTYmVqiyB41uwmXqV8+Pls4uCfU/aOJ08UxGy
udLEC9in6Gi3d1hGwrU1HVtw23dElEk6afXclh6t4hUSWkLSAD4b96ko0ONf+3HZ
VbF4Y9wALRy0rI81uG5Pd7hWQAWGxKf4OnYej3qRhTWytYjzIk3qzwL/Hv2+NLAo
UsuTa6DQbh6ATAGRxALGRM+YwF0KsbN47TAerT8+J1loHClp9v3dIIz9dMZFVh18
9oYUcCJ4u0+11dtqqYfqgC4esPytCdhRLAj7+cej+1fW+NERAYsgZJ/8A0OxXkpa
/QBWd3G7DoeJatwiYiJRwTvvEwhKPbL3DSTpQkdY0Ca0nRFXXIyp34bFRPNjDIP2
MtEKS06aM2fBoy0bPHrqdeFupd2Lb7UH13ItOnuNFD/pIo45kf4WJAevZ6FX9har
S6YEz3RNoz7lVvoLd/XfTHgoECKgZuavUC2mFuKGLo8PjuURlNtVvL99/aLspsv8
El3c+U+JQARL3u0bPe/oyMLFzM9EuTY/jYr1Fm/YFSRpWEm9vd/P3HWT18jQ+d/d
aoty8hY+ZH2PyHMhgFlznnAMFQFmNvhrbXLxnHyBeYrmbf8zZFVoESpm8zWwNQP+
znu7Qp6HcNQoARFeFDoq7Tq7yyhYVL5+ksSgLE1gltSBe78cbLJdckleoJ4ubaYf
/QsVnmLM1zTkL+DKYgMknSD/Qo0AIW9rYcPOX5+jWTxbpJxumtpBozCljjFHb0nI
24p8g4aU6k4R7uUxspSSd/JiYbYsjNzVpYv7pBUCr8JFNPWalGaqovJzuoLMVm/4
j/7Qzx9S4dBs8hWY0Ay/SwCk8XpR91Ee6uFwShrC2z4g9hlQej2JP2ZIMA+HzNZD
b7kQvxHTTWi8UPdqipA9nSWHPa4/no0keIf/weXPXMnb+6I+Fp3PUsO3O4GnowjL
z0PCGzyTAS2OqjRFtHZNkoPaiQe2k+sX3rpOMkKJrqSrbIarN0Bctga6RH/wTifd
y2Y6MeYiyivJebf0s7xcI32IuWe6rT1G0a7Pc5+QGiwR2HPbk5W3HkBs25nK24+o
P5nAORAy26QnmUEx2C/QdAJ6Su5XHlVUKeWHoZq4BFa1Lb6N6VvdUqXS9wGO+DNz
eV9tCmH8wimN8kvwq8VLcjAJctmq3Md/s9GxBys2aTRQHCp5I4h1vAS8+LlHfmV7
nQ54/uIFGZ3QGELL3zj3nD4A9EbP2CujCQkpPehr6W9qvmoLB9BUlbwVsy9hmhFq
2DtDxWzsUIg0NqWc4yJMBAch/pfSqhvbkSsf8PKpIMv1/PIjUIAV9tZn2Wsw4G/O
IUbNk8IB2BShStWLjWbbkbFOpLj3jXsHnPqpkxp76VUuejaxUDnldCoP1bNPUwKV
6q2dupNa230Z+UeLLHGUT8KDoDKanCtlTr0yUeiQ9vaPOUC5LZ4pdN9zsjJqg87p
Nm1fJ0AKma98uBKJ5AfjH1oiDun4KpAqK8ugLLJHdp/5/qaFaSg4whFtCHmNP8k5
OVvuRqqB+J6I+pBWbRtufUHFiXcqwg0LBL6jNUK9rfTkVojSeQ59NnoIFZE4cw5S
aBx3YXnC5V+Br2tTTby/2tEXx1YEykzV8Kkv3AW95r2hTpi39hutrA9a7hHkpxCK
f/dOkLflZZKznYFI4ICtY/yFASB3/vDNp0ixJmOMmjiSD2YWzBkKiGauOp55pS6+
u8R/IuwS5+Om4dSvzpUs1xs0JglAzruqycdcGb8y1wJ8+awJ6JowAPWUXIdSJjtE
2/V2RBWswFhJtE3qhIOf0Ju80cidnktrOjpHOnUiPaxl7bhyR4JdKE2eQDp9qwal
g4t9TpEeqlBtum6ETs3dzl7yH3GA/CyORQNn2F2TYZJ2a7h3rnO/8sKNXjtrfdaF
lT3TvCD0jSEHiKe3yp85Kudb8Riqm26Yy04kCOtOsi9SQ7rriHjmUgsSGgd0d0NQ
m1XOMoyFi7TaXBiETxOg/vOM2Vq9mEkA76ETrWxf6lOZ0Nv9a/UdiemJmab7kxJF
4PSc1QH3EOdaTOw/bzVNqBs0Uuej7XRLM1rDR/ecVD8TUI6wmZUIItyQyoj5Y5sl
thAlXyob+0vN19+kArAVzD6VQonhkxyqmdGO4FOFqC087xJ2Ln8iUR02r/RA/obT
/+mcPOATxNf8Uz0N9gsTDsq7G8ekrfowmiFmEhYspNHQyApZ3LHON2jm54xZm9Tg
T4FOjXS3mQA5HQUVqWFshi09hCHkX6WfzzsajcMHb7S6KfBiIfSk8GOxd7LOwFLW
0Ppao1lGx6gyBrEGW7D9BkhYAOGN3+5/g0gnEWAzQE6fgCXS2cco8l2RaGCNGOUI
hncdR2lXZLziP7vF5bblkRDb0aLZ2fatfFmAFrWo1No27gPEYwHrGkxa0ywxirF5
wi/DCowWlx7QsHI+LtZBW2YLA9jqdpqQKbYfGwMYMqUbiL7PQntFDJ+IBQyDsr/y
Z2WIyWRNwRO4Ueq8ShMslWsTs42yiA13GwM2lzndgkKEcPvTIrc28mIbymmO17YW
2pGmr3KCfbKeYoYARigEGsb18n+dV0TQavh5AGa/Jrs/1Tqful2oi5pi1fhTXYAR
QMKB3aZ8tOnOLO98cL5k/O+ytW/8gvHXSFmxQE044Lbm7+b2WZ+SStVbWngKbsY+
n+J0tNGyq3JGBn9UaW3VVFN/Nuf6WcW19qbXazjMkvVmTQCTE8so0FZXi2vir7Ih
0bhn10Eek2DnGzIJ5bZp4EYrTn6vtGMjOsMqVgpczxfPjAcZ+mwo2bssjlg5r9tg
OGf4gJgen117zJauu2Vupv7tFfqY4i1GTcgb9pGTAOyVP2tMhhd0REyYiXtJ3qvS
kvki0fUTKeI/JfXHNCNKDl7Xts2peYHX+uZrWxP4nHvmypjI9sDFHaIpXGDP7aU4
dLGI8XTUxea4p7mzeXc9w0P3CkFazuaWh2RqVta5g+sshHB3rN2uXkDLXGfmvLQE
IN3c7qHF290twdE26VpGb9t8zu9uW7FXMRicmYjtOa1mnSJh9jF1ImuCeS47nz59
55H1JnWj0h0eUH9Zz4MM6UiujvWyyFCWqVi9yo5fgW0Q2R//k4/Vgdn3WH5YiAEs
R24mNkElSQcC3Gf16p7+El5QoZQ17bUWb3NxpmNDCCTJHtt8jZIeeuvgKZCnFdvD
5Wp9R5gVihEmri638JuCGkjroKS7+50072vIKiryc2vVW9jFCJPXmqsCl4+aOTjT
q38Rrqb/6lrMpCoA6qC8/NDSn2nW0yKl9bWRO4nhDF3CgM0WR/tBufHhdgSfn6MR
+YDJOKjT+NabV1eqbIrGV8nN62rqfAlE+jUN4O/4l90BSC5o5GtlBTD1YDvDfH2h
GM0C+/9jmd7RAvwq2CGT3bCnsCO4am8zp0gDPEc3GTx2PmNFgAdpbLXZEGZkPdDs
/vW4UNgJhhEf5CF6Hco4omfEJO5vZpbXJ1OabqZrcfIg1qnjlBTAjiUFmjMoJQIm
Nkp5pYYZdYk8fdHIuKqG2qiJ2W8PwBpiHb765h53IRVOvU9hOgRrhqLZXR+SmeA/
jMP2GEoqsm+xX0y6VugjVL3K/D7lFrzKI0j9AUvQd3UrjELiwmsEb43r4Bv1ENri
N6kVLnHilJsYUmA4RhsZU0JzKPw824ScPmx6aP6E3TygaQJG2URfiyq1GsocO7wG
eWGN1ALFGQAOU84Lp7h2kjAOFaljUnk22bF+6u/i93Q1sQvOVb5ShEQ1zmj0vZZB
/SwCQcMJsymLMV1QLI0Sz3G77Q0ofJa4cBfmFxKr+8W+k4wi95D73nqRw8N9slH4
/ThuWtcTk7ZTj2A7onL5UdNt/T8vV9eZgMaXU+fFHRCdbAvihpTa+4TQaCejOjTz
7sezvLtTHR0/IdW0XxFQI9yU/fJQWYHYJFZkmRgbyzv4lXWj9R/PtsT7qQFKKnU0
SLk6y6r7MIXGRwWFWwt+IjcNuDmdA10jFfhsPe7mVOHj+lP1/l47c39AiErGVMl2
dIWjjDpJnckiM5pIhO0xX1icqY4eBAF/3qEvYy836nnYm1k4No+ENr3ZzEO0R7Sx
U9LpYN5qA6EUjmQUIDAp1vz4AhoD9imkyLn18UrgSZWNo7FP7A0OEZ0gDr8OVqPD
8W1vTecOrs0cGn+kRxNRHei4reDYgUv4qEynqjwFi+3lMaR+Y+GnxoHafyNw1T/F
AZOSKrP3xPWRu94xu2e8UKXiJ77ipMNMUFv3652sobc7ouVCcwr43+sr53xE1Sei
65ce3rWi9CWFAAd9MQzbcDGiqWdBjLXmCq8LqtZC96afGT9v+V8ZPBS/Dk/Nxw0j
s2/Eo705LrfD082kNVE3BT+G7JUhHAYHhM5QcHshvJRinRl1NeyPfNw+a3ltgeFp
aytDO0erfy5i8/1UfOab02FKFBKVhUqQZB88Q5vc9ly/ODkPWmM5EBdYDDme1ziU
l8LDTEe4YXI6K8lrSua0bGWjhk2jh5dsfkvXWY5Z80PA2xOM6S5Ax0sRD65SNc5b
LTdCKUCKN97h5+x3uax08916ziECPilxnaYi4vd986TW1u5SXn6M7dL0iDWi3tJZ
2G3+6oFkmdTA235rQOpJtcFpCD8rF4Ba5RgDEoNWvf4LUtUTuCnOIguGpRp2uj+O
jegDAxCGYRr3EYaD78DjUu47VJXd6Jg/NwkXcbMsuqjEk+aE7kLZr5ZrwPscs9u8
iUUtIFXoXuPawrWbDj+bzaWNHhMaLZIeFJfo9Fw9LYSlaFdTI31PFK0msBD4nD+c
AIbXYwSc/rxOg+GiwDOPX2nXe/rAUJuJLRu6Q3wRL/uT+O7u0hqUmG/eTsqdxs5e
tKL73f5TjBYNXFVUyUTuzgknDDt+fcX1AiRqk3TmDX7kK8sA9QuSpsPEE/PRL5ex
2VtRABDsZptMB51DjfFxbdGC79p+sz3eKZtEgTUQkJ8x5GQD1sXLBLd+QS0kNHv0
eOlUWji+fYmCO3Io5dBnhrvS+j1djUzsanSndT1AfNnGqC2j6qCCVAUxelWtH2tM
JbLNeVujm2VWGwDpLEgbHxzkPkxWLFHTSpQavEwnhKQOo+C/aQn+8iNxSUHyomud
K+xCBDtLJYBoIeJac4nWZfX0kkQEQigBob4tXnwvnGMx3stqJUG3xugA5S8eWJYx
jqTN/v6lBDpjth720EYncb5TF0zitKFuNVGslZGPgJzHPjfAZrg+uIoFvbP7eTpd
9jcRVVgBuq/c83u+QJYT6aZhJbm7/XyrVP1yDP3R6dJuiSq695kCeEcOGkhzPqk3
dCTUztYS+A4KRCkAiYBgTbAoiUnL9niR03pe6zHQcaih6v2yXUsSXxSpY0LFzwMn
+XpQ0b2bRwsK48OQcSE9K4WC5MFl9myxkRFk6G7ZULnOAZ6tVCZkLic/kS77y1uP
sQb+xYwtmjgl911vW3fPTcRlK/tMGoxCD69sqSqG2zFiWMBi8dGlbsD/2aXapPWT
tC28RxOSx9j5chnMsuhgWGDS0VTzsK9cwu9vhtgOnjhHVdDPbGAxiZkTvhSt0GaD
R7DfvkNeX8ScydBWaxGsSVRySqO7mrNwyHSjK7m6MvBiSm90h8FYC6NUiHMoqThy
LYEdDWMjzFdmEFNdlu1xS/vJaqMLOTFlIfJtM8cdLgSDY0LtLEE9Ps+h2QvIQmAF
M2cojXYkt7R3wvoJsYp6dWFP0uh2olF27YBkeGLawRVXmUPrKY7OVZTr4tVlrnqC
T4q2Ca+GfP3i6eZBkRztVSfyh1CEg+Aj2lz6NdNpBdNZNEl8VX3S17VsCIK212yR
2xD1W/d5M2xOmOMRu558UqpjaYLco73Wq2F3nm+bM0xww/8W6Yl1aDNyh+Q/QHu5
TmfbWsCI/oCS2pQ1zCINGau4C5FYVkmHIkDt1vBB2I/CyoIqc0LoWO5HgaTWE1qP
WBxgOdqrlakXmoJzQ/zWN3xSXVugqKBabkL4RrtfEOu1tl8TKinzmJo/LbmTbq1B
0IB8DiubeQdPZY3EKfqFgb8v1ETcHYeyKuX3LLnXSfNiCw9JF9GG1HXBaeheJ/y1
tyrfcsbHEE3S6NK6XXGhr2hMm+bd1pgFGHD1qx/O6GlbuNMNR+PTe2Oj+a+ktZq9
E7u6lLW4zjKDo/v3mFiPOIesx8Z4yH1q+AX0aW+aJgRnpXCN9ixElZVeMUc500p+
FUj+AjLbBtY9/NwAmMGro2GbjLFy7Xcxwx9IaGAY8eVeSDButuYBcBrlw0dFZB4d
gi68tQkCS097zsR/k3qxRkLoF/B32HdFy73sTrHQGRCUCz7E/K4ljks3pVzpa0NM
IU42qPvsdRMpVY7AF4ENwIKOWqlRInYh6zWkmMxhGaypk+W0TYZM76skcQGTWZg2
VKqLLatkzzTlKuOOyPWg6nbbBvERRbsUStHRMByPIezHYAqoDkuKaHZTEnyYGoS4
txHgkiDFaMjyA6IisTVpbaFsXYKW2F76tAFYDhLo473SlSUv0ID7915vc8IDSqHB
AfVj5dbjBU5e5DrL7UbpySojudQuTQ7qHCdds9CdD/JpOKkBguJVW0jClII9UJ+v
RZoeHkt/blEOfpGverqznSNrdDWL8S0tFDIwXHCnBBqom3vEgH/XP/k/3cGE297g
w6qpNutXs6lypw317Zp6MpJ7MK+K0mLeO2hWbU25HLRePNAofr71zvrl8+XgTYFQ
O2I86YYBCQwwxepOhQp3ue4QZkqiCvN+ih7vbhWF5wyyGXoobdMilPZtzD+yun36
3XbZqI0uCjH6Y8loNOFjB0oUvVoIWhz6VAXkXKLtHKehLDRfy68ZcoeIsDPF9TX0
kXdxMD+EnMmo52INu1O14pgAezUMZLVo+Vtwix41FG55SXKsbxTQYK10SfGXDWq0
gsQa8YF7fBFQvFBosZRWqMqXrApah7dSIdE1BFNz/FstEiz1cc+eui+mM7oJI3JK
wccWxiQYMtuOKfoiy2UEWOAzP4EvF439aTpikvD+TJlzieEXUVkU5L6kJSy673+o
a227UMj+6bEMINKKSwVJS940QP8tN8TSBSs8fhQq3ANyIhVECal8pl53bjQxoNq7
okR7lzuWUTBZlPK/H0mbHZdV8nUiuEiMTeM0BeopUfKwVgM+v9RzVFwnrQRgVVLc
AgE02IxRW+zvi8ftKaw1tpRraPOA87hmb8QhtkuR4JE/2WdfyiOpSRPMtC5WlF/2
dcJgDzn/VjD4p9wgLSTKYYFc9kvTjLF+50RmR5Gq0cTmF5MO3Hh0v0yYMkeff2b/
XM8GauLe5YpDErtmY7VGG+nJHeBaJ2nWFzwjVv/HlGiUIS37jgxQav69ExFq+v2g
YeRapHkB2YYz+4R2WFNNeIf7CEzj/QaV6qA4RfkN6pXgBxl+T7AoFuu+QzMiZpuL
vhursziqQVWi/9k6LQEsgnz1f9QXhy7Ar25sRj6NT1YFVzZVSaXdJqq/aQ5Vy5Zf
+CEMEPJtBSUOZrUG3qGoRp+TSlPAnUlgS4Ragtaf9Uzm9jMp9No3mt+BsVLWDZKb
E9o6eUH5wlIUGNt6mXtlV9/A/knO+xHCrP1cTEbkb0jQbh+ksLpB6Kp2Kkp9PWLX
yK3kZ1nQqbW4i/K92VKO9973FtLHosaoMpbJ5TLagLcOfanbKJX1L5EdDMhKE20O
7gSrP8bJOWPhHGCJ24kLIH2HblorUr6rjSxhB7X/3RfNAHbBsnMl+mWBK/NDoilB
UMAye24p7EM4DHH5tIGkN3pwmEGduTR9EdyUthOL7/yJAP4oEOfRtP9wdWDT8Lg7
DyuZpMeEy//zHEkPnbCgPIPNWHpDx4oiMkRYNTzvem4Jlz4+r0t4tjVGY88yxZMi
T6oVZhzMRr4Ht5m8DPL4ev7I9adEd/3kHwDqzN7XzkoE5jU/nMid5fpEeR2m2PEg
VQqq6Iw472tdsmJ2StK8/PZibpmbH2Pes7e6+NVdGKGOXFWmSF+M6n59jvWYCNP/
pSDHibOLwL7GutMg0IPFO7d7x4SVNf6CvKiCdObp4BflsupoYksH4hn7kUHzfAKH
szNnFi68YF9GXTRKHXaH6TiOXwMy3NxNL+BV2D/egXRYNYmvJUtKJ4WenL0TwoAw
yC0aCj/cr6Em00d8yvIt2cNMUS3I83rHp4Ya514mg62j/AKd6u6fRnq4HkuNYbOh
dEc4g0eJRO/bMmWc32+1DGdnnphTj+GhvxzdLLcKaatPPCF3NP7pEXFt07EF1En4
xwT1AW9jBDli0EI0qOUGtGsb/8SuE97PCiCuCAbQ4PUds6zrqBjSBISK9LRe4RS8
blKo/h8ePPHn53t7gwoo66rFVBPKr0H8RwXKflK6cq0O1af7PZCPqyU5rHFmwZJ5
1vkMrXHseWbht5NTTx8ux98QTwtUQ5qg0YoGQ5hMh5nerB2fFPjji5kj3rue2ru2
HoEz7jlo36HTIoATWbKO4hFcbVTKWCTVSwPlg5Z026xScttMEEvl+IwvDya2pY/3
q1QLWgSVuxiPLKHBORNia9tleHejYmtqj/UBwufe268MCWfV3WSJ7rgWzplDrMs1
eEY+zmdKamSdh3u5c6BbGBfxS8PRQoVs+/9ZgBZEJFQXbt/OhLMnqjN4YB62Sg2N
xSAH+gRyBK2jj+a7DQougSt9pQxT59BRumHfvnpdue+NFUwJH2atT+iTtZ161Isp
ynIVaag/TvxVScIfp13yWwjo8X/djJh/3HKIKnoqEPIjNJNz4WhIKBtuGichN5la
xNxgjkx45ZiX3/eNbByjB2RtxnnjpMk49eQ1loAtS38HciS/+0L2J28S5GfHE1kB
PY/yxdLKzVzGL23zdLUmSrooo0D8mG/HFR50bsEIWmqiQYdiZUUla4iOepE6Ln9q
TYfe3O9HMGH2t+Axca9U0LduCf2p14sLHkubWJIkJ8sjN0akeN9wske3mO7AZYOq
hIXaRgG4PDB7Oh+AjH1E2+PX0EZb5g60CNv/GhBLIswJU40tR32QAourMbtCFCcZ
b4JHI1el316MEGxRUzdRVHCAZqSNuUj5pITS9f/aYBgLRLnpxhrnfn9fTy/ifxz2
pr37CPrDk5c+Z2zrJoIREMqBkDpGx/mPrdPad8opOd1MhztVyF5p6bmf6Q1SiePi
V3gCYcNbGoKf5OGUl9Uqc2zfZUgRffbfgPY7/cayXFDLlEJECJJaZqaucJ4S3XmS
tNtS7O8/FDvuP7G+BNvhGqdgrRqWv1vUvHCVNB30e8SSE4rETjGQ3fCpN/uHQdR+
RgmY6+6S02W9jhxPeZz1Tuq7zcIRs2t4t9pCstpH3Nm1GQ0GvgqXoHDKysStziuB
rQAWLkHxrE6zE01/xT+HHv+5UB/vGHKLf93cNE3sLYJz3/sLL1sssbI9G/5L/+U2
MxcW3pllke6y8JDzFlNV7D5KmitLlOzeeZA5ejktHc7rKYqXhaByWWqlJltdv7jD
tQ6heUTxmXGNiWWhK//74RJET7SUKCBBP/XfFWOifYgB5Q45R7XXnADg0oL4Gz0H
T03OSNBES1b4q75WxnpWsgbOVd4rJGnNssJDQEqJyYdXU5p/3Zp+1jpbjVIYy9tN
r/H8ADi2WLiwBBAN0xDLSaAl9Lqv4ECUUD8ecm3jR1WbCmn4LmeuJa10rrpLuAq/
1LdkOBKclxsBiZDyPTAWY8bbDBECYQiGe40427GEtkT1+kbioDETox4YcrEOqCeg
ywUcTjfvmlyuXgrwrtXHQODMWJjoxUNn71gMl80Rvz4lN6flv5rfplzzzoT80olS
SqtetWiaLJAvc968E2Td6We4SPkjFLnBCoigQkScsNFdjbZ++C2zJVODOZoCHzz6
2t8E3YEZ8S2OEbUCn14X2c94xwtMHxyM51KwSDZtpogkPL/JIc4wsViyIzTRsaXO
ZHYL0IzFMr3jKCq/cANRFQZYgkyfYYr0FmlrEY+2LLlKN5aDmTopeJDDSilttU6T
Rslc+18pw2nisTJoTSFFSULCnsfwiFIvHlGRBHzsnoD3dstg0gj0nk8/RKYnGkTk
8djbEF3Cpg5Q17KFJVquZQvdEoH6jYMjgIjV0m8sbX/3BcjDh8gI23QwlvNo13Yg
tpkzH/Oy2tcK+JMoS4mDMpzlu1v1/nB1qky2mYg1zJSmH4MO6qfCj8WFW7D+x26/
6YHFUsG0FwesLJXTbJ73sm67b3i79vt8kBTATcfF7ImdkdNUMMgUWx2x9g+34O5O
QPUQBqX8CjzouhZyHXCm0cgvT/ZO1AIxENg4RL+d6PqEiRGHrujfpwNJrrFfLZ/D
zkhvigdH0Wt/zf1ta8UxbU3yFVB5u8uASGYfBDWwdaULWJEs1SdqbY/OZ7E/TvIW
LnmApQoDn43/7rhyCxRGZW/9fzUA8uwOVaLV3Q1QlqwbNRRe5aCRa1tG8fdFCZzY
LarrcOLXpK/NbAKqABgmlBDjBTmlFAfBy+bu/Exhyeh/joibaVYwActxq6ND36uu
Scgw77CHwSPgKBnjwvjnqYJ7+AI+LyaQUVvpcbP5JZxGKpCK0iSQsJbWfUGlecWE
UF5ODjVCzebtvhixJQr8S/b+CsR9Xu6KFjQYg9dt35ivkzVrHx1jIQIIBWUCnjEa
DKSiPJKCE4ct7USpfrSZPHFB03Ye81pOuwU6Ajvw6O2dD7G5w5LqHyhK3a6psVMB
O7ghbxf5c3trRo8IyQLHyeienV8SSt/RXOfYCgEucBfAVIr3a/U+3jBgl1+tuiD5
5Ax8X0XOUJxbrFaOJkGkil76gfyuLWUr4F2jRvpeLoWOE9q7xemmkWAjOY6eIiVk
bW5LYKJSbh55aW0hXEeiAMHr8t3uIEiXJBqvLknG2KhzA74BrKZ3pexNrdvY4L0a
mwrbdHtV855j1TZSA4YknAU3hbSMJQ4cIahvqO6kO2ARZ2IE6gg7XfOwe7jV4Hkl
j5Xd1QChYNNtkv0ZxA5gaoc7rpXnBQZrF8zwL5wlWKXSb2X+IVCNN750GAT9tcmB
+GMt22m73YxhluqYtgLaWozXwog4eM1fQm3AKk7nQ2QI+BTugcI6cBYT3J65BLrv
mpcEQn3MRYLUIOW/+5Uf4Ww9ZoR/UD9oEDM3rnjqGI7aUd2p8Rx5om+A2nazRc5a
rmvmc0QGHQR5bXc5bSMvgGkuvkemhIbxUChqqDLF9vrnEx/1fqjx8IHg4W9NGsyo
3IERQhIyzHBjB9yENmDLi4z1FY35FKhJezD41J44twugCgYcNbSZKx6ecja/7iT+
HNXCQxJMkc8uGqCWbGlrFDMlq9/L/yrrsrbrpAZo8eSThDNcAPnp/+mdUdOYehaG
OOx7g1a2w5xey6XcPGdE6pR61dCswfyxyJr4+VftGmOL2cCrsZb9dgDOv8O3w/uT
VPu3GttN/ehWcxaKfbHGpZFouQmZQ1kOAcKWiBZ3GpOBdx9uvbrDjt/6brH/Zuj5
hMuk7Wt+CWA09HFnFVk01n9q98P7HaKIyc5I+vah/eeIVm27pXWk3twH5r+ekR/d
MpiKvo1StL3ljBOtgFe8oTgj5cZXxVBzLf0YYPwYJZEtkyO8xcDP956f/ViKF2dc
2sKTkENR1Y4EOPFMt42LsYAKEWK4n2apntygbWspRK0ikjOiAjvjQdoGRf+mMJgJ
nBrfGQreN/5PecuNSQQotiG1tHZY16S6hrZ6o02udcHD62UBd54x/RQKzfR/GhKE
5t3F4geyGwde4VAiczBAkSX74JZADtHBmEILgvMa4xlUOz9D+0ZgbZ1SNtfoTvNF
eboqtzBUPdM/uXoEWjhi1ETca2DYjXF24MEzi4EgfsGRl6IvHCN7h69DPr9U1azN
9pVmLN+4wi3rNKNIt//sskd+dybYJQVPeW4hb6auwopXn53wCQIfnjcmwrd0Y+TX
j9jVal+V/korwkQ6z8Ax/NgENmTH3tlOn8gg2/Firx9T1k5/g7DLt45UvUr0Ti9q
GdGOSZFKlw05KGE0RXTfXR+HZhUtbyKb6D4mIAjquBGfCphjIQMdaxAFW36/6UzF
aQh0acno6DelXms0/m9sIE5vbEzP6ZMVRs4TFIZjB4A2n3fj+4DTpaMK2CsU76sf
p84GUXRRCYs00+VLz0Ke7FU7beKURHvDYxBD4zpcoEYImuD3xbqm2OUVc0sn2qLk
76dLHiytihzy+ZlcVi8T+8fXnXl6yJtNkBc+Wc5VpSRPw6t18vsg6LMztsY59Ees
cacjdAY/oWVFuT5ILCMA5mMHKpr3zXApX1Tz+T1yJwM66Ahx54oGc6PN+6gpthjk
kGUBDe46Qg9m6QYL/HAtIlQKc7EN9QrwEFi5uBh6lW/suVEsAal0GyBaA5x5bruU
yTJMNJOTWXe7hdckNqx6ciNyOgYO00XEm4c7WdKYTyGESysdMtrULYdXPg7EhnMd
RMrD6rdjHRhNEHbPldZ480xsjmU6aK23+y3zjmAqp7BDkPp5GeWFdMUiLat8k+pU
h1N+t1vdgfz2oA6/MZAVqrsRflC8D8yXVIwYC8POu3sNc3sTdCyJ4BHxch8QfljM
htqCJE+SQbd3VbFXXjKLGKZRLo+wjozMS1urx4PGmILTKaH9mIu1Hzai/401tlpg
+2AOSU8sfqS20k/vAgySAq8Il4Qj11TphuExV5348v+GRTF+7DIoYgftW7JGOzkR
z+6lBfmo3nW+xdMgGmpBBVkavFC6KHy45JFQvTBUnKT8O2pbJlUhBMKJv4VnhsN0
htNQXWqW1o+oTvxx6QOMTdeQ3nWQyr6eyO9f4TVPiAGSRI5QlIg4cAEocQVszCOi
xONqGZkmP+eMgAZ+xeFHDZtFBbtevlWkS65nlj8/2C+DelisRwAKfdpEj0LEkR7T
YKI2Vb5L/rdIv2bORU+DXg2l8JaN2xCfVuB5XyLvDYCDpglPc/70aBjByIFUg9DM
//FKkk7f+22Kc6lNau30PYtXweR3xPCZE9FlWUC0EDh7qtj+phyaxGQ6ws1R9W1E
zwTlzidWfoAJAH0Fir0e6Dngy8l9Zhamq41re0CPfzhO4nRKMjhSdvQwxyJU2qjk
eASO0HVQSAXYkLSDfj+mqfVgtmG+0QISQqONS4r60/RPBFeY4KTPk6YS1cHUmmZB
PT3cwftZOozoH6eXSSY/cKOLRHwKfkLoQ19R3taVNc0qaqPIFHhBdjjgjJ+tZpOL
yPIdmUO1OGW5T0Yq2iyDG3xvW2P9iIiq9qoBr40asqgzD4Ibdm0NmZVVlLDo+Sgc
oNSAS1qf4QtcthWXoXvv791KDXhgCFePPw35Fdnpu4JuxkGS2lKGS0MKHTVWgklY
GyQDJBYzDHQ2WQifKGd0JcOg03uiNO3el7wyOzd6iSZDM45y/lTHPidIEUu2phH5
LzR/lv6A3aNIQAZNXZFcPnGJwDcph2t6ulJF1Ttyx3K9bocfS+LOTsk400CNE4oH
4PFsp6TABz5La5psCV4YvWj53pPu5zyP+b4qq6JqauQhhPtWYinTJWcQmi8RJPPr
6lT8zoXVc9je0iwgUueRYJ9Eb9gJ09gqm2XwKdN/KfzAmZNoDPUH/QPWj6uKL8eh
hlDenO3czL5sqUXpEF+6ioPv8kqiQSnwiGGbgvWIxKxYCZnZPFVVI6mPP07nwAAo
qGyJB+AkxWfwOfNSpu2Z2TRObUGgE3snpVrmyt8imGP+rv0wvRFIKzn9F9qlKEgB
ipfFyJKECOcLDwYPrrPnwu2nqbv6Ji3WZM1G0gF6t3QvP3RxSeXGRIh+pApnqNdW
Qf9GzAYMjA/qNjVixZ90qybYxxNohn1W7Ezhnrsm8QoDmIKWkKcStmx+f28gaSbf
vD7W+exwh1DfV/bmqppXXZ5KMZueFpKRvleKTUuc4l2zeZ3pjKfBsZBayDmcQ7do
h93DNcOoXAeveD/3QcQYm+DeL+EHx8tkQpaj0YpV/zVSCLTZvmVQQle7G2/Qz7EB
u3h4N3hERHjlpyXitL/gHmuHixwqhLubmqz8k6zwqu25wc9ozlyRDQmmPN5pXUMO
G/wH6kDJ+/23qUJ0TXO1mZJL/ZVaQlrBXWZCEWKtT5zOvMabCFTzWrjyseTZlY6B
UBRF0BBw3YtLAgPME0EDbXEU8rsBdgUxGoxFXybPd+Vt+auB4Pr7iuaZma3MoMTI
QeUqR1nkqGcSLx7JyeKBxCWnCEnD7jmTmv0cUGE02wjMLmg80TJ2caE4wVj6k4YZ
tvnNaCoicdSAyKweqPj7zbUBPYF1JxlHyW5GAAfCulxT3M6WXXr44WJKqohzRXFu
HCZMfrNcCbbI1GDiP0yoANwFnVSqqEreZdemzh4Ewkpn1HI36srafPi/XuUyUiIn
vMl2CrzVcrvoq/ZmUHbYc6XixAZdN/NVHAQoAytLZmPx4z1l19FyAWdCO3O3pr6W
N1WmT7kmFBDAQg9ag+3dsuqmmJj4V4yYEAvH0fJDDLocxK0N05eMFjNh5POLd0+U
KDlUhwaLO+s0P4dnU5wkKJb9Fe4oDsCoOZmxqrs15+1wsZb5OL76Pj9zbnx1nYl1
rokZUBohvHdG1DgVU5Acw2sH4/B2ON+LWqHgwhuYy24Idldt3RB2HLRr0xZyVZtc
nJqESi5ucslYfiHa/9W+7bDk9JfVEc3dTJhLQ9bPodERr0IMlifDHhIfyqJTZeYD
8Io91KrY0LDq9Gf9u3ro9eQ5BswlD3GAWFi/t3IdXkofJQuaA9CaafOy0e0/gFn2
/BA5Ck8qF2zN6CydFrmcabx5Q9ANDiE2gbaSiRDIIjd8IqhDtvR1YpN5YenW+LL2
H+bhr+/helnjlS/pR9cA5crjiCo4yr7a8ZI/keb8QWRpM3u4474oTALVpmkDdq1v
4cCNwStuGw/v0a+5aw+h6MKpxatjy+yYxHJVyJ4GfEm507hufNzcSq5TgBYsWRnY
WvnBOf517m9zntV5nqOebpRUFsaRCS6BDJzoNlA6jOLMjgtMP3u/cZ3c3cXzdGTU
zAlI27ny54uy7bRUwZQt1BJkW47rR/s4riol/7VV9ENlYmY+DQ0e3dWYITYTTFOg
Y1aZltCFHIQB6unvDw9JCnhtlRkvkZlBWASbY5nDMMbguoxNJclEgmaivD6xmGBo
DJ4t9RglvoHXO44qCrQ/U16yRxBqeAzK9Ve4Es0HJQIZRUP/9l4K1RkWwaB5cjJS
PIC5UdNmLn8LtMS3MlM937CrFt/0V6hp5Q4noiCjBucfsrs4DaEo2dX3dsQPUaq7
LlR/agfrPmZ9vqhuDxosZOpTMCiFNgmolujMb4evcPBne/CekKOJXBwZPAUNQguS
94mhkHsCSCJZZibjHsc3P8qw7lKSZ+S9NRDFcOaTKbRa43Dq4BR9aWkXJYWKw2AS
Xv/JLv8ZeQxPbCAalxFyqYVrr63bZKzIiqtNkguyu25ism4zxmSScAub7SDaxDNz
gXqODZQbwuYeqBd3Vzj0uIkcaKgPCRMYpDCwEiiDX0E5TSp/ZtT/KsdU7Kz8zW5v
lrN2U4kMzTQgIcgwRPRpwfz+Xz6Ec3655djnzkzqUGc6zOXJsV2FY+zV5lgMsXE7
lw/MMkIoVrTfrE8t6Up+aSSomN5bH+5H0tOR3LTHNVdcKfF3pg20HvXv7gmGFd81
0/GD5g2IVIbXsCXf7Ewni3lQZEUXpORHD8tpiAWQBZlQBfEQ/iqnaKPI8BvLI68H
eWrI5SMxnXUHcHqLJFN8/oRdSEEu8KB+n8sOLYeQhOXjxosfgdiJEU4uhXoztvIH
1dsLSCNJuL/vfGiU1IcneodHH3By8CD6jIqSUYC3xehnYjRZ0dWvyrjafh2O1Eqy
FuFxxwygwaymoplRViMhk0h1IiLuVNRey7dCFWrpU+nC/hgbps66/uU+kHlWCe8i
J7nOj3mkAgK8+m4EO8atFCYRO6c6iZNw6RB/z1gD2gufSczbxxPWLiwoZOweR7XJ
I/sGWGMqS5V0qdFQBREmHPxOZmdQy46jIpfVuHfpuekM4L5DnkLVbGPBUivDCff2
NtucSPhUlIc/SBOfUPUy/0ryrBd9DtgpBSpOzdnEyzVm4fRHv/2/T/ZVzJTMBboS
/4dk21ft9OYX+ZWNaiPCwq7d+/7XkiDNvvsLIvnB3UCoKwy4tIs0fznfP9LVpuU1
Zb6ITj9+etdMpYDXcQuVP1zxCwcjMG60DAmeR2A53JVaMovNqj6YkZiQrdxZYUD3
ohBmWEJbdJlcqVr+vBgspzB53BAhTdo4VdRViyyIuTlgcBkeDBLIJViRjgrDN8mY
yG83IvEQ19GwnlyfZN7v8YipnaL+jw3fYKarIA5nrOMyGHvtWvDrqGI+2bX5duWS
WfILsjxhGMXXN0oTbOiZPOR8e4gLB/rgdPTvaaBfR7CLjMyqDTBrcJzzg/BS/w20
K7/Gw/WKJ6vA/40dnZAGFht62+SiKNbUSUe3ca1D+rIlAclGgWzpMNua/hr9kc3+
Mhh3Sy8L0+R5PWIRfdY//RmZ84Ep43mKeVCrF3zBCwffK8bkJ99L87z6lB5XkVBY
ZrGBbqTMISB2esSTu3SQ43eZKyg87WhgMkvNtKY44OcA9PWhNn2FjAO3Kqet0Lbp
kvD4/Y7CgkPDgF2LOc9Jzfrkq5Ry+sjiHv2hTrDdW4Fj5hf4pC/VIH2OCwRn+CdV
QDGDDl9rAK277he+Jq5WnXNHDcVQFYYn8/5JReRH8WglJ3EWwB/dqCdn9xTJ1tvb
AGyiw9QQgjth7CqGmR/JSJ+XVZFc/kPzYi3to13aoVTbf+H+sbslqeliCChiskAV
zHDE3jLlU22g9I38Vk8HapVqcx2YF3JHyIpcKIo4EpMBrC74YeR6JoZ2a90nyxEu
cXw6Swu7Knsiwv8IDkD5fXQAPtHi4L93Rctw3G83QA+M7TnuooJuC+L7OaaVVJLG
Hqa+dx6zMHlmVLd+GO+qOW7WgTQsSaGgWv/nG0E/JJBbhMqJkaBXbZcnyUcOwqRV
1TQrGnFVkHBWd0xn+uBM5c+zux5ZWmrZoELNSd5AjOAIMXwiNF+0tT9E63bXCKSn
BKgslHQ7ZDkUbWMVWxOlyDKB4/dsJRY5hvk37nPUNPbfoMhcFJxo2hsxvVH8aaDF
wJrCjBbEI86tFeqsXTHC+3bAo57lNdU1XP4ldkNyNXjsk2f4/vnZ9LvDIwy16eUN
yvSqd22T2iYW//gDopUGe36t92/onFvoDadSMCyxQlrcsKqBydBtyJ618bFsegFq
in+9V2TmE8bDVx3Jyw0kIDUkQ7EiYKcYCY4uijQ4n6bYBpUAlYJ4Yy8NlsHrze2+
sxs0f0b8WLIIOeD9S/kN9lHWthMW4ydJH0jTxKqqhZcJcLVLlImco3NDDP2XiOwG
OEBH/3zcFeg+A4blBtmLBGm18xlhNFKCCo06Dgmn0qYwbaNPD8O5LPXN1kgt0laC
bkP4QuMUZ2bxgkrl4XYyMchd8hV6VAdnzlL/zC+d9fU8jljZD2qHNP0zWF4qYjki
5qweve0DLeXiIavWUmbAbLHNEt0YU0Ncgbm3JMRwNZlZj/gEJX2fYmB3jwHg3DIY
gOLJaL29WRsU3dlvCGzXGFZc1lz8Hx55tm2SHOx7ZCLhjnNjqxYKOwaEl0egWfUY
m1hty/NaNyqQECIoRQE7o3xsx3lm2WQzDbsZSz9yOhPVt2gGASjWKO6yQj3nVbik
kn+Box3v6KhpW7hzGkiBRf/eRi4WHUgHMYVq3WOJY9Ckj2e34XJQk8cVr6k7nKM6
G0g/wPjZZWBSFkEVjHeDAq18n+ZjxkpsklqzCN2d73MuIY/7K8QYZFsESpfRaPE9
UxuJuwrMutDay7RlBegmp518OO5uBHYaKFKXzGr1hb2TrVY61tpWhFmkfIWOMLVF
rYicj9GZvXl34figRqP/eEmtegTjv5tnh65S5nGma0tdhbOywLWncrZTlAgXtyuC
uyFFRK+VqwnC+X7nRUN0CjQ4oIzbeiNQc6bOhid/+XgsgqkV3OepmBFuIC6DpTi2
RnNLfGRR31uDONFgVyW6UMv25LgINJMB4i5jYCP5AxK/O6dGIeXdZ3ZVA1/TWEO6
t7+paIB+2ulViJDYEsK4bilhClWnVCaUjY7l2NowNO2nvg7YJFODxf2B4AhDnQ1i
qiajGxS3leZLYh1HVCGHgy1Qqp9oiGstGCJX+NDtUGX4StfrvJ9qBCPbiASugCPU
HOYe47VU1kglTyPPJMvK6IEJDs/lr6F74dkpmn3ql8jg7ZiHooMwGP1At1w2BWQT
R10LsLNSKGI83zWEAzIwXlFPv6NPKy0EGDtpzudHm1oYSC3x6XPPXKSfZNHnBzbt
sCsS05DH2xXU2SLu34Y+LVcfFbFMO+enk1e97A/92NSGx13BGCiytBpUo6Lo58WM
w194UH9uGVIaQC+99TzJUJ6SS9Q0hXVS/yGAWMa9yTsZWv0WmLooQJ656M06jy4W
O4TjrePFEX6Ng0jdysGLuTZ535twNSzBEiv9SgPRCM4KZOypcuydwijXq56S+7dO
AX1xpFabGU4sKeKxzUJH+0YyBJGHgdzvm4YJWUQi9mJU11jSNEfNRxBO096S807I
4Kctw1rNPaZ668HBjkpOMbyPtWqpRtI4GQm0vnur8K7++XDzh+xU3SwCj6JW2afd
EYaiywY+g2YvSHlTrayXAMIG1ZhVUxmufExG9/a7DqFWHjgSlswjz6ckBkUFj1Om
WF7AsBSK50n8heY0rajIWxOYEpvX37GU5ZZyGrg6L2632eFM/4cbZ5OIDSQuZTN9
SyOnZ/NkeOlOmmQs5/u8lbY20qT+lexp4ldxEJcYXMdu2y/suJAk27fDpK85axQD
NneFW630C7ivxEk0pbaOgJ5VFhKtLm0t0wNMSWSnfa5ovEsTxVlvR2WoOMRtcVUe
ueJhX7FikU10xeBMgJySlYllRedixsLR5U7ai87dKH3bF7WUNfz+kMdDYHBZME2g
hYTqlJlZoNzWvnj2WHV0FmbrQ4TU+LdbpQCyTZSlnAOKcyk9i/3wM9nQmfgAgu5s
vIG9Huu+OKgVQ6jyX0KKS8WBrm39sJbFbuRvJqbenDi+XLiQWYJlwV7/z9IjURBt
oK+zukHfsQ26WKL05/jH0Rf6vnvFi7Ztz9JCbr2HfDhe6/vpQLpw6X7ze+i+uATe
RE8JFKDSQtspM6KNBZbLWWi4UTa7upWc9t0wZb5jTXwiIhUiwbdVlwIIB0kBlR6l
tdakX4jccmaYs7mkAgATkhPS+ninqVMG7bm664a+9/vgEF8elfescqRP/SfpCoED
QqV8CoBZ34lm+rhmzy/8WAZHivnU/kQ1D6/pGH9o4dylh0A+CjI5Y1AxKXCGu1z3
upLZEW6Mj8wMtkA6vOYlVArP91hbkz/MJDh6+3Jplrf7qdpsCAINS8uAHEVLTovR
Nw5xKjOA22k670GAnSn7U8w58ujkiZOksxngXJ+cgG8vOR3WkfxFUG6NgQWiWc1p
b7UixouxJs/HNq3GenxTVuMRxUle6jQmWRnuk16SmumytDRVzB0VCMlRXQ0Do2FP
DppnFh0ZyTtExdr9bDCJnNNVIPMse56KUcoYq0NSV6m3ffOXs62jFgLco5qGk7tP
R/3SMGewt6fIcM20wu5ShjZLEIflKEIsAqG/puG2xrmSoNt/mZWAiDwRnXeCPr2W
Yw4xEIMlXERxkKAaWkz8f+0TwOorD3yhns2kgdOQpCITPrdKx1Crt3VqzUk5W10K
A5EjGBqSfYq40QHsAnjkNHkDKD5KRChyHAcv/F6WmCXovntIFGuO37DZLtT6XHxi
XupdOoF+RzabKoD27NxSVSDYNLqnig1FZEVAFAcR39sR/MbnnqKu3uBtRHjRWTG5
xyLGviFXzjk0E3/FYMskGc1HcijJPUvOiFWcH0u1gXOtKWg98RSNB6W+DRmHIZiq
F8dxrNHQtLH0ducuUp4CICeIsqu0VdqYgNEbNpRf0TXTRhavSIBFFzhChwQES+kV
Vdg2/cLzk3XCJqu4s4lGozn/2d+N0FPXN/XzzMvU2P82MsISI3+jQs6Pmp8GHbIJ
h9+HAz9eY/wRVThjDBM+t5h4hE98NgP1qj+FYBuVRZkKM0etqqmVahEQoHwb0KGm
Q0fy1TiH/YrgSIRDxfa8dtU0YSbBBzDI6LZzQ31HxqE8Sm7hljtHjrMjVduV20YH
D74UQ0Dl8lhQG44Dt4e5GX0cDGnU12L1i9dF7cT8f13A8DhSNfDPAffmG5TGEXEi
TKjY5gaSFUVuBIaDWJteqJkAQ3X+al50/Zvy108FrAlDjp753vj8ZL5+gK0eiIdD
u2XPuLnPWgAGZY372AM2kAIpdzM2Y2StJYy5nrJutKSVr9Fz2mvSP03A/osfoDDg
KVk+5WOE2AMho/qqe79I7G69aEFoYw16SUiPxh5XvO49tR/SJldfne8JEePKF6AU
EgHh3hsqOisaf0ncl0XNyoTmh/5jGS/UuJ3/itP9Y33L1hYCOq7E6OSen5wyVSut
F1wD9y/r6m0DMpPNpF9RKwqJ26WcboPfumoX8iBMsB7RStuEXHdZa/N1QdBA1nMo
DTKj8tly8mzat0TEla9kmCTyHioNpZhWIhJU2Nfh3Dlt9C9hdhZACnC9/EZPhgl/
kPMegcpj9+6EMj4vjF8k8FhA2yILVylWwDSQfP+VXfBXzMgRVPrIIxwi6wooPb4S
96ZxWifLDxTkYGS9juQ/41iQw1Nxz6aCYMLwpUFTuxynu0uXv1jGZHdSu372WW/7
YZhJcGwNliz9FRKgjz8ouZ8qqCEbB0K9FaoYv7ovnF2aQgjbsoYmFUpo/8bUCzEH
4j33ZUXOlABpVrSsfHdkc4cWiyEoSFhWXNSq5SRruFvbgqvg8Bl7vDKw0LBxkSDU
vLjcLatc927RxnTesan3TjXTCevszejxc7m7QY12tZ7QA3CmrWmO3dFSrJOgDw2d
R28wdcN30mumlUL/KJsARy6qf37WVH6iUXIQjRV6DfCbKMMJNBxKc/WU/HQIxBVx
Gy3OkJvSAayoc1kXJ+duCRmUlmvwfGFo9ToAgzfRmW8KNxskkZRFlLi/Pb2Qt9qk
w3binBsm06es1byBDYBygTcyqQ/QKlslmxShgg4T4pWqUvV9w9x4VvKuo0dIhtn0
TTfXECfm9M9nBU9VSpLerKegx6wdxyoU7K0y5NZK1AUBuKi1suVWqlmCzpFxgsj1
ipyhZ4plX0XmkIsZLCI0Pqh7LPXAMBb88VZ6SwgccGb4A4CFduRKw0lUDvFYZbXp
zTFZy3AzQ7X/ejFpmwcNtFtTD+H7YFGDlFlJ6UiW7JcNo53M6VhNw04HGmuXyqcp
ZDF/fBW6yPW9DgNYK2neSXAgKsl3+JHnsmyRWUfynbhjGj7vjOzWkLbuLknjAHvp
DnCs4heIGF9RLt3HSkCs64xSzP2x86b6UJE5g6AnidCyI3vQ+ZW7zjIdZTZwwbgt
VoE24iQM9J1M0wykN786s+A9Yb2NFkGwU2ZUq/ch5jN+gQzYU7zsIMaS4PgbJQTI
eE2MkEdl6+2osAtcsSuBw5o0P6+kRV5hlFAgpQx6n5w7Pu/elU1EYgV8cTX71Aw3
T9U9XbBvGoN723Sb1q4degmbWjJoqIqByQ8rY8CzS7XfZwGGvfrVt1U0rMaYbpyN
j6Tey6EkpoTBky1M4oV6YYiAQLMMhoYxeY+Odh6m656vZ+sfG07D6qU2lK6Brf0r
jDmVhdQrtY96W8i0W8HDSEoK9tQP0UU/V2+eKZ9KCukOq72kdYjEhlEJLUGGzrBE
aleWphulAJsTSKjSeVOtfFYF76xrkuO5LpCIIgRv8zLn+2s0XLaw6TOSLEwohtuF
Qwap+0+Rby/Xg2qqYl6PU6eSpTSU4RNUpVkOz++5jbcFPAcjmPDl8oSuJFe++WFa
u7/azvDKuY5QwDWPw28Q+04MRiMVvQC0b42vV6K0S+i9JlicmaEIfCKDi+ainDcj
7kkQcFKoFis1mi48YdDa85kB8hCiWXSvLtTHY98x2oB+6/KRJHjtD9/qY3EaaByF
7aistME3eywD8qQLcVpBoMSi61TOgxgE+cFzZMMEGRV3X+ooMKdzyX8BXxjcKfzb
6IU33dSot2kCGgU8z/xMVV78Irj2k3Ft6eKAnmxktRUAKMwHMYsMOAyyP+RVh/Pn
K68DZInGFjh/qdOYt6iptoQlusbRaXdkTGwTmxyU4glGha1NuWINuCpKWkuKXFao
6wuIutCLSum8u0jrULO4R5FgXD2+rboNxvcbsRuKA8dW0TuLeoTAYZFAhj4iOE+4
wFb3dsGSuLpaGCYDkH1jwmcbxzhXSkAq9LmAZb2SjxMLoNQrL6qg4fy5OdV4JNjs
nbljcfqV7A0Bt5Gl1loYlJkunWoxYIzXmdpfO3o0bkSKht9BTNZONFgA6F6lhegQ
R3+h3jQjXrj6AT6zB9CS8GO1Pdn/lMe61ajTVhN9rpCG+QZNUkPbea2gHbawwmId
fPA67CUsQycNdsQiPnNFvOoLqIlUUXWf1/rkci2TK0ybt6w45QfSwBqp+XQkPatg
6d007z/tSHQ2hDAAFmVQmKFRLAZmZYl5CSHgVoXzBef3S7Hw+EhIwKa3YxlAJYAg
rhRvsqWIEzo2A5rXdxRBK796d+/8Gfj7MvK7njexfE5v9U+3avC4XIEMGDWuim1b
SNlzj4x12yLktl3iP0xHObk4csGsecZ68YkCVupa6/iY9O8lzq2DFt/XoQiqhWil
t34Dph09zWOQmKB1+OVjLUOSEZEMpsPjS47Yd1tJnxNnhrcfc4f6TX14x9ZX95MR
v19Lv6BdwHFXGvj3mta/oRSVne9H5wvqhlnlKGKn9FQ4fRmOnXapy80LrM07C1si
o/BubijkN4fyNXmMdXrnPrRHUTpObJaoZPN4EvV/dG7v3GECFtgbCZl8Q/Ol+u7S
RrE7eda56cOcvKmcOh80CWSc8uVbTzTPx/jdJahFO5o+fqD2ifxoamAlzfEpRgHC
m3I8yyGMNwHS1R+CFTWJySN90TSp85aKKVcBzxUZk+mxYPRa/87a8/osQD3ZyISi
W2Nq68tMW1mEHbJE+yqAesWgkND2WAouL/+fiI60+ZynKGr0y+gW3bgMBpeFEUY8
fwWflfD+gjzQ8tv5r0+AGfwvzgP29V3iYWW5EV+kcQbUplHhWkqPob7uamD5vGKv
yxc35iNK4vPHz0Wi9rRnSrll/7mqJZUW8Ddpv9YG4La7RhgYzcqVZtgJwP50kYgj
eZ7ng4xvnoP16hJTAJK9kQAHaQfwAJI7kwW89SLZ5eXk/O6Zl32kENsGHW50hnjs
VgPAitG+jEhgZdLZldYjUzWEMV3MGMi/l24hoNvxtfTNoGUnhAMi6emIRlqJjKFH
4oJs4jTI1OZeD/fEQ57wRqG334CaMbE3GMpVo1WJgi1Gfd7gQ9TxVsq8p6NXSB8k
6OwQPvOXGoabr16c3ww1ifBf3+NxIwkXb3jsDaPr33S76PCT1bfYXT4CoLtfBq6L
1wOrUOu7J69AfB4La4Th5P1r9x3jsIQpPRXIp9KF66WREr0V+ikjze70czfg15wq
smXAC2G8rpIhER5a68j9AyQhx4L2Gmkau5QGhhx8/deCwq0WM5cXGCdTrOfgaA7E
H6aI65Vi7Ul7D8dj0Ppcc3+TcNrOHZXqPNtaaC/CoQBztMg/+PT6l0vor3ABzbNB
h62tLb8GUIW4tU717DaGtmGC/NF9dK0zmNGqXELdRw9N6CiiwkQ6keFc/YYuuA9R
WN17ZAae6IB5+Rla0LS4UlFpIqmZk5mGH1U84e40YRqoI5x8GkIhSm7EdC4vLiZC
KhQOh4NSS2ZdL4QdRtVdRYaWKb4nRCC/sgrAnTIzGUEtiRPexuoY8u9/uSA6x+ia
2UI4ORVGEgVQrQaP7a4FiqvfC29bTmjVj5aBG4qOwxvMdgJthCvsC9lL7RWiGkDZ
egmRaEpsr2EbJbAbI1mCrzdiO+aVluaOg+rT3LAQ/ggX1/CZiDEhP+afr35wUKk+
ovxMR1ROeMPA7/N/nTvOFeF7JlonStHK/ssrscbWlOBd3eWGjcy58o9VODbGSB7n
ZTfo+FOu9kka67cotimnthKSUOxakht4tyq+hy8kR1W3f+5NbmeVwBytBZiDMx/L
cCRh6wuIEdcnQFYtHPnKnT1ar2h5GROXtJQmcaPUa4uxKPl5gqxLJny2P0vC6QG1
hJMA60CBqU7J+CTHJ2WRK6y2BB1DE5OhT33h5vDKntKebpkBqMvU4XkKm2L3/ICi
burYw4ZU/aZUAkm50SKK8F7erjbRX4f2YvqIyeqX2IP4nbJEqokd6SQwn8WzQaQ6
1ijpnYdVUY/Jpv04ef15VPmI0W34MkWL2+5emMtShUqcdhOOjcqtmZAIykh/a3pE
5HxcyPclhpeCsP+7BpetC4uE0d5iunJ/R2o1m9tLHRx338C2eb1mC0Et3aIzSxyK
2t+WRDBl1HC4LyflIGG3FoI3e6ut1oODC7WhJ2t93HmTHeXDwiQiPaZP+mjF9rgi
psUJPd2maF3hXa3ZFxmhgOxRif/YKuFeoUKKdG8qFPlXsNKES7TpO8rAczjN0zUC
r3TdH6+ITNKLTH0LkAHSySCTQzTqVveTsABHqF9AV/lb8pPXzIDU7w+CC61M5CWz
SzFLfnlCamxT8aF1Rlhx9/9n0AloTGqal49b2G3Pm5M54hvkHArodrOdZdXWHTQ0
THgnbHVqbb70A6tPPCZoCweP3N373jzJqBVN4hGbKmoI65MRhFPTS6UIcoJSIHvh
AIWaH399eNyAeBehgD79Z9GVMyJgMXQRMLHlsC0qhvdI7pcDkth777Lfyt1gGhG5
uC0AEBcVrt4owPAeMwWV9PGi6PpIxpkE3ci7shLuLh2m20j26kT3WR3J/mKJQnf4
C6fSdroHvHhT2b3c3m7AyZXqpwHOsTgMF6CSoWZi6e0tl2iJylTrO3D8eLXMil0h
B4sx+AYFJP9jpVRaYY7364TI1dUlNuLNoK7KBnJaQPNyFK5b9KzbNtYGjZr/Ga/9
qhdewvJypv41r0xkCqriG8HG7KDZwQeNZmADoUddAj9p4IkH9Tbnw54PLS22PP7M
dz6oWqb/EUhYL9Ygj/CRiqTscybN9IFxN8qOSMM9CTIGAx4W34/+shx20T6TAXLr
FCFRL4pbEPjAuneFQhrl/HkBBwDSxJ/DRXRCU8wBFj0PcZXQps+9tRJyE6NbFckm
xM8EdIo+7uRo9o81528Jh92jvRIEQZ+8gpb52usoync0wjnHoNWHMzW7Qe1r9n2W
B7govZjyTaNo2kMgnELpraCW4/CFUA+ic14niWW8K1IxJtyE6gFwcyB3BhIGOan+
WKZJ8DwjQ3bI56AAKcn8woYDny4bfpPJnZbVyCgAcdaXYvefmqtV2IU7+jAlak7Q
9cG8ntfzWfGDsYwcXfde8QlW/YrQaVJf2W0WpUfpYbXvhM9o7yuWuGFn09RcD2YD
unLTVjGisOH1+ItgA30M0SC8KpiUYrQShATViRh9YBDNI9jefI9VBt1hhJOZJgpq
wfxJ7apb2qYvacP0evy7viUlZlITDaa60ApdRE5UO9VfuyRQ6ZU1EqKz1MxIcjW7
OPTmwBYsFyHsUAu89Nh/DnMi8/Z3Pd9Xk5q8fpKNG6TYgU7MlBzGw4snRwCuv4aU
zEem4NqLWZA9R7Kq/2mHTKYRSpp3C1VDJGU0hmxM5o+SjjlOFUPmUY/LI0WkX8Ea
285FD7im1z+Ky+vALCRuHipGzOazMA8ELJtAKtg76dFDNXljsGqB1QlOX0M6jb4C
0HMIX5bhLkkUNnUV4aN6+byCgWdTJOvbHI5zKNdUpqTSWxPtTz/LVfNGtubQylkf
YP8UPERmzRDX+X0MnXWP8O8TSBvYiaOVUw+W2I5UMcJMV6WRjNJlXgjPBQppQvHw
yLx2CfsgwrLOYIMLwvaT7DkIfHNc+WxbPsNWv4a429LFNQSJe/qB9XxklY0LgMtc
mjKheTw4C7Er4TU9FmC6XDFkqvNdIVlpTdSDBy5OGh1Yj4FsHN79lAzkag6Lzujy
NPcqopFL1VIDWaJ4Nr8Yw9Tw9Z/I/d8jtpM1DmrkFAjkjrMyljLyVJMnM70TRhm9
TeJiYgPmO8AF4kPNuBMmUeCOMtKu60HUN2GWLrXNNrUvYX/nOgbQkaThLmuFM17s
AWg7FlyZQh5rxYj5Bg0Wlul+j0w75d5ZdquhTNOindg218V9nTrE2dHGizUeQe1y
1TbGRpgOcTQMVJUEdsOGtOljfPP/laKrZKGjNtiuVozy1yM+OcD8I6Ji+PvkRi4X
XgpaEqNRKOMo7V8/h2XA+tAqqxwfjmJKiyRiJ9Zpf8ciMqK0va5j5X0IhOvp/Qtn
uWgWur5sru3gXMJQfPOmH4zS4qxHLpF5BTb4bGbH4nS8WmoozY4ZTfby3y7GiJwK
BImHiuDL5dGOB1QvvY7DkLHVhdWBzN4x3YsSKKInHN3ee80odpvBNzWAW32Y3VgN
cJ2aNavFYZiTFgW300SUex2cI4/JGXd3oP40YY/IbQV1Grsq0LWQv06DTlDlCXxG
7rHBbfuCWQqPzPr6D3EQiKWMCjwZ9kAK8Vh8uU8YnPLI50Sbea4Zs0jjoDFrKg5+
w9LmY0cWKIioNSlaIGM1twf2tAZrn0M0ewJk4N/e+oqBtnADErRsLvqAaXPUF4gl
DK968XSf3CHb9WDkegMmA+aPEMGKLxoXztWH3gGKeGAiapkhlniUNbXSCtPE+uMF
AlMZcAeOUUvCLevTooKhlnutC/ueePRdp0oNi7s8YbHy3Gc0IwdleSGROBQ8+WKL
b2lwIk5/3VD5is1L4x0ns2eLJ8WMUHYeLROi0OPMIlCySBpzUjLF2cscpPVh9tVV
GsbSUqXKAAZxfP3oKnxKFe6NqylziITOs0G9hcFp8opKYrgWUW+4GK5CR3aGQ75C
w3WyMTPLvu6e3t1cniNiRmmX4QkznhimJmBvZ3i9Z0xGU6retUzZvDOdNdoy+p8K
E7DhdHmDjLkK66vWqQNTAXXdGyD+sVstYs9gPsxNKhYExhpgIdBKjlnfcVIb7s/4
wVfHYRJqRgeG1I1HbZBv6X0ILXNLPlLYgQ/PCPLbdhioe8HlCBg9PszN5X+Doqk9
DE8CeDKP3W0Iask8x45/LXlDHz6XXOnvPGKMk7wve/5nvTFxLSN02r+YWb/6javu
9OXhwv0Uazq6yogLS5RbEfcouDr7gCIMXHurTbupXuEwJR24ZMC6PI6MR2pbV5xY
gl1o7+2yidO5RqzUavzsIWaMq9bARKUV6oMsY8Or8s3G26+X3jdAJ9ogJHfhpwZa
T6mc4P/VHx826v9Ufp8hVedPjP7TZ0B35qm0syym4GQDhjsaf8LucFaMWU9KjTLC
Edc7VQEsmTltCH72bn0zt5N/h4d2zsV2VNgHpPyvbO+LNGVGmNrW4BFgTw/RKhX7
JpueVpzYTG0FXOcyDzEhgdG9WjI1qr47g1dst5WGQR0r6pRsdCFPA02YTQHN+Wah
rmygGU6Q9k5GKJpcPhE/1Xr/dZSoy5+V0HhwLwdUPvslH26qTq82X4q6lJsLcubw
3E3XqX465CiW3QlWBWZNy94JFn93nphAmAujuzXCzgw0Zwp00CEKO3nJfyF6b4Pr
pXPLYDOMnGuW1hfyF21kZagDH9JIIiTgHIab3FcGop8d9mJw5tE4sr5hQsplwpM7
DmqTW+cStwJvlAmoYEZVAC1kuKOHjbR3dRWdc2lwAHb8U1Oa7K7oUp7JqATMfVT/
ry9ZKfM85Sdzx+W3Rg6Lkgl8Jq/PwkbxXCKVOJNqZyY6euw5hXFuJJs672fFOKrA
HozMlpz0W7GkBx9AKI3LzKc6tcHj3/HFHoqK7R9kpHK+8QbMxhn0ImenxT0NMv19
uMXwGkyxi8e5B9LxJ2nv67GWDL5S2LTAEnBfGglQ+Ea5NN/FSBY8QN3KcT3S3D98
7HDbXv3dqvJYw5gfQIijancbIuzQAvQv+B/VJrzXRGXuFyhdNrqMdBI63m/4UiI6
/oC5oOBgeqLzQ88nBGaLNDzq4hplHQLx4gmHsYYnm9aPNorI9utTaNTuQU7OgYob
fNwIKaIt6qiB251CxXvesxY/poj/BuzeTEdljC/vZUPWwpAGdneXzFXOb+kHC2KB
yvXTEJQWSDsrYj8QeTKRA0uL7hxJLj+fj5fJywfFuRrSr5twNNg4mypT3P2oGgUG
9SNBN/M0ak4hnHMwlSyDBKHZTFczYFmPv96gifR0crvnCIh0bS2i5AbjKirRNCWq
tWSP4n7jIF2txv1k8tfetRZ3BQjWKKn3nRqYc9E5+9ZKXMEB8QTGIO7RRQDoBp2D
0/aAjJU83Aa8D6KRrgi6m8cyBcZxRQadojMyZTu7zMaIoY2Lah4Ed1QJpp9tslKT
pHzmY5Wdu7AnS/Xw2tBt5X2kGGBeE9dk0MpX+rJLJh1f9HIVO1KkXS+CvL3x4z9L
0GBRaex1iIO5TzcTp3cSSLLte3mOT9jbePM1jKxSxMUpo0DRjErpdMURxeL8Jvru
SMYy5lNmOvWRgUztcWrZYLt4iQDDEFmupITEAohNBV96elnRSthEETMQkKfUGAat
WnTWbTzIiCkFl/PpTzPfH6LcrJOOkyESZkyqOdHCn4StZqukZhzQqNfLebk2DX1t
tZ2EWA0MNyLtVTFCHGMj2E5eSjd6hYYKpwwQ/5BK1pjFF6h8RWXaWxGRlxYPd8II
/CGdLnRmj4Nus98zbZSmOlnUMElLury715qNPKiihLp5L6maQnxISByPOZe6LBF5
HbePLuaFgIS9wcQRlNJvhc7ClUrJVqx0qoaPJClHyS/bq033bcIu6Od67sZ/oOe9
XRFsbAuD4vCS1vzo/muG1Au0eC/OMX7tVzzWa5uxqolkxJ0IrpKsJxfckhKvXPj9
O1JObFuYkbDQpojJIObHoDN99a+vv+ptNgPNQSbHb+eZ7+vmnkjc3wL2EQiHdmr5
Z4lOGGlspkv1gPU2YjN2gtKayZWbuVFGIbj4nb+48Lt6CMHWhXR7lxzKoK5x9cSb
TP2WO4bZ/bRdZhGcHZgCkIs/2LoiNOSrZcViczlI+AzGrQ5KT0cUXpTWYylYdKMS
SQxRFP9Kf/fXtYU1kFAvqseRweyaGKjibz3g4XdUvQpVBwXAB27rVximkoJQtzF8
g0EiNSc0NcCvP3cRIG6TwOxXOXsXbLu3JFL6BNZWTDkez9UrS7MyDVCUJsPBF0Mc
nQgUN1pG4nYUORvbxjzgBHI9HpD0x91TxoHN/WJXWb4SGy5zD/0c61B2M6YjK1Ob
QS8BSresI/F4+TmnvCOj4GHDryqNTw7OCwV5FHgoyVTRDnUUjav1R3QAResPNjtx
yx7ugZiO1hvEHmFRlMHOOEoplqakphS99t139Yr2vKyIij0OnZYaZTZyotZy2jFX
rZ1HCJ7q35CYUMhQJOHX9P9zGxYmfHc3FDCoaw4FbwfIWMHI7jhg/b/pcY8OLvH8
1gjl4h0+J4B26RlayLU8aSTLCcPk3EK0HB2qmArj4xic5CNuz2uI83Y71c1sexQF
TK49gPt1Hxd1Awn81JG6wErdoe54aSRPj3m/xSr0byke7eapB6ySPAlaWsk2IZsi
m5N89rOIq0kLUfC7cgvzD5YU3y4QImuQO2TN8BDr16t9IiueCjEXKAdQtqUSVMCf
mscn98sQ+cNsVmXYy1wTmmYvEnWCnWw6H+vn53QcMxKx5HdhDg/dDDxTeyWWAgIj
41xgFPXY8oLPDBtBdn+7MQEkfM1z1KID/6yK57qtXkbaU5p2xS3SbuiEzsyL3y/D
4NQ3PmXGdNO7UaBHKk03AvTlM2xkhVUoJoqVoONZJakD6vNaqs6pTWxjEXdQcuDE
P/Ng1bLUnSN06PQx2FfC8jjwzP4vfYpanzAr1Y+AKdpo4Coq8rAOxNvzIZTyW+cr
4l9Z8guArDXQyjyUTKYB80YVAUzNE8jKnbO8gmdmQ95QOmU4Nu1SWA7OFx7oCouV
SnIhW1PO/Sb/pvPSdE5njFyxUsugtPj8ZvdCleNP1J5t21iRFG81xeNTJ41hV9u4
DWJuday/ntXfIJUTAV0T8vlKC6Yc8W6+r4qgx8la3OPf27kKio/DH0v+GbuoSnbx
lbhoRes5WpDvDkdu89rZ3ITQXfebjRA7KlKhIEfm05qXQpbzFRgdF7gxWSSL4l0w
ndp5/tDFQp7A68r79SFpnsqMYeth2XFUI9kns+ZYscpftQArA/xM1bpGpcDYztCJ
TE5VVQ4YVLnFXE1bJRtz9ImkYWbEmDaSoJlEg/dSnpZmtQGu/xJQOgFSOnUxKdtf
J3y1VJ8AnNBbZ8BQeghSDVZb1ovYuOd3Pa2EpPthLi9UpX4h5AkPg9VOF0Jultym
seQrcTEoW8Yzz1jzo8cUf92XE8c7pWCysNn5x7ee+rcOI71+HTn6O2LbbQlj8S9C
gbllJ2YmtSM7OuHSNMcNR6y73ccec4es0JuoYPi8A/FNsdTawPtZV39Z8eW4d6jG
GyBPOyIpeJeTXB8TQvbtnf0GMI8rYtoDU3kt/q0ylXDWxwA1srQPZkKsijGB2mPa
8vo3UgPLkFswb4MR/qri8l34x95wasnSavr4St9r2lQtCFF6lkVHFdgA6FPDjPad
M6Le0e6Q6RqftDL1fAFc5jW4n149tvlM3Flw/USWHsrnvXj6DX1q7wuvga7HGY/F
aLK+pptV8mGShNGOd1pGV5lkftewB2in2SKojlNMiPKJBUl5uYq+4mMYg0u5/q1+
Gvvk51w3Lx9BjaWpM0+kO1hYUHZZrWCdUz+zntn2zsbDHxhuaHpHYc1uF/ruoHW6
cQPRpdxm2qZ/hqzugRIW8cfN5O/EXhdP80hEQL12kxI2sChseVLbex3/99nsRLan
n62Bg0Tgsus/QKMqoEZk/wWyuPuxVCA6gwqDkbRedyv5utTSW8K1qM6ICBQ6OaGk
AQCYk3EDJdzY3rQaY974q6QLIYtfo0jNu2XM5+5V3BMVLuEB5aCViD8y16hvJyX/
6+x4UFKFtUPGSQEMMRsOlCSwCrvJGWTA8aXxhUgoUAar5PwBWzL6+hrbY6f2M3L1
SHtvYT9bMyXsGewWNxPhLpzxe7dBAFpr4zb/csNCP3L4gyPK3fnxjaOmBIKeICKw
di7qx2u9m5aBJbydWDdJOBFsIN4P37HnoYXNxwXnKzw+DP1EJkh0ED1bCErn7kK+
Mb01mOVeyJwdBXA0QjaiaHnxtzMcBE1s6OkuENwAnRjO+paoFaQjLVK3Z9bvOBhe
kofTtmvrhS+mfMFn//dE4VoU8745VJ9FcAPNEIKM11INe1rZzuhm6LNdRjzoq4pr
M4qvAMnF+JT0qUfTuPy4EfP9L1UmsKbogNIqyFuGJgtNVQ19sRAQKYasbPSQu5Zb
y1bgaMC/DYsu1uCRJXUBrXQTNU5srdEZxccz/J5qvt0OTS/yEXfjo2BlqiFOcHS+
aze2bPFmEyjJAFy+VHxv2XrpgKbev7VFqJnbZ+bFahoN0ybdFGbl32yHu3tYuXtb
2P2DNPxr3mTuGSmc8QiOz8nT0ZdnJZWESmUFvzOdVXcOwkUg3IIrOKvhaTYGrGWU
sCQfii0IKM6JcUGisdv7N8BCgwpG1o6wys5Zgx9wnqCGHCeMUgcy92/l2BAmx5sm
GRN1Z6lmLlSIaFw1EdrE4UqfsRNsHYYDlf8L3TKA3zE8axZ0ec79E6/2f6zM9HWi
90klv/ViaolYi+4tmrV6rOD86cDTG0e/nzBU7g44IiPRn78faJmmbL7cdN2ou4mR
hcad9mtow+2IT0nofA2qVT4Vbmip+AW+C2+ouG6OKNhKtNJjEBOw+TUVUlAfq2pG
tRRaDgTzsnoQc6SerMMe8kYDegJ94cZ7TjiHFhsjZQLOgUL0sveGwIjcNZfXEZ4R
MI0ElD9HKxT6D9nhqTo8JJO93J+pQ5N43uW17b+Mk02Q/yc8ENUkJkdHGqhkEZKT
iXCVOIaa8u2A5rWGtkjpFyecmOGmg2GV2OPw2MDetJC5OkbT+ae7McRk3m1I3fPU
MC2JNKu0ukC4UEir4XlJdpgrfTO4Lwam2e/9XiqzdLMMGVdFmHeeZYkP6JAMjIIA
XzJD5IKrd4m4sh0wrtftOm7l5cg+t98w3d8s24BhfkFF7FVmxvBYGQjo78Cp5SHA
BKUSu2lop2COTYX7R+PSuEYpZ8o10migzhBZg9BpcgUaFjrk0G2mXE0NPNx3kOCa
WuE9QBOtMVlpdoLe20MUM/alAEUJ2N8x8exsRR8AUdomu+9U2IVISPomg/Kfbimg
H3QOrcLpsp8Nz4nzuCRhs7mJDY2gsojSb7iStiPD09FPJrgKIAl4uqKNtmazxhFg
+XUWTgTKx1+rn65umYatJAmgXtHsSnM9BIt3jDHufht1J11+dn118U014IKseVLj
rccbB7D9idf7qqNx5K5Zhm2iCyEz3cl+QLA2gmZSAXiFcLiaEli0WXMf7jvdPp8e
waRQo8L/FNUdNq8mU3Y+lN0lKM89m+yLDn+9lEF+H4yWrJNseQ7bEsZDt2hJ0fz5
qQOj4x13WBdXojcPpNRs1dMGFLX6LTlheMcSVq2PKVeYCgAmKOi5CfQEI+O98vo9
G8s0k4SX3kwgJkQnHKnCy9Chk0SuSbNWhkH+jNiqWhB7g/0sT3n3mLurwlVhk4Dr
ExsmzeDRBBBAmTStazB0NepoOQPyWSNQMIQKfAbJb8cCDBNuY4NSzpTh1jdA96sS
vdQKC7SzBXgkOz/p52tic3rUrDfz2wUnKy5mOJSFpfYF3fgezNSwrC0hhqXK74X2
E1yFr1gjf+z5nfAMlc9DFQHCWh9W1MmHsFBNzY1UBf+RQB8uSDHFpV8/d1jyl8Ql
dWqLMU5mUviB+68sAIL3T+deAnx2LhuMG+3BI76JXIpax7xGuaY3FEfzgC54bWR9
ecn/MCuj3rkLByFMSzkEfVJZHD/IiluUEbke8Amsg3AbYytYh7jPMuD4vSZPwdow
1JBaX2dMi8HIZh8aJuvGGYuaQe+ZHEsPe7p05RWDitf3PdUB2/UejLNbdrrjXVRu
Wk2uDktQWy0L+G4xZeSTRHynDINVrEIvmoKLJ2JKvdyyYvk+rW13+s+9k4RgtoxA
meeeOCVkWI5zudx3GkVK9lyoQU6oJpcRQGbRIcmpeuftz+3suT/QMdgrHh/3Xvi0
NwhgjfHY/Ah5sh9btXsIIXMLNXpSFcuiNmbD5tFj6ug/9u2b14yoVsIfPLQdtVt+
DVQFVrzMjGDFb4lqX1R1te7/W5Eq4dXLidyDtmWt70zApbdqP5DDuFSCxutNWYnS
LrT32/h0a6SU8jmiSPDnhsXWz6mp3M0KKg4SyXEzViKlqKhZZPsi3fFlchst05se
nfTiqIf2NGy0RmVvI0xTlGekxgjdEX/ZriB8UPi8VvcwNX2eIN/bC63AXkFJbRFy
pIqz6nSm2IZQkeggpjWSqWo5rK9AFMjO2sQ7d9y2OMHcWaeEiyjEeOUApelNjazG
P8O6aNR42eGV7tk8w38ojKSm553dSXCb5uGP6VaD+xKDHCoK3kpUjrSgsbXA4ww5
TuyUWlAjxQtyXUF2lmAOz5kZxdihSooqexWKjFfOE50fIVDd74sESgcAaITBuFtk
VQQoky1v0/mrohPq6PpF2zekdFH9SLobuKFPPCchVnT6rhP/5QOAETu8lC48w9Lx
B6C3uqR97m9GeDQUO99sbsVbG90MYYUzqX56/mwMOJ47EzEYbXmr/NKn7nc0/dQ+
Vb1lga7R5BUaE71+gEdnkQdtjw52NwsMqa06qQ2z/0rUMbZnXef7fq0ohzqoSLWY
uAnVc9+GGpIMcDEyQrMWC/ah8nLWk8ttzpQlZ8hobZsqCMASKQAkuTZptakDXdV1
RlAl0NDCdhMDWH3HV9sRGpJrYQ7gvKaPMAp2EIXotjnFltGyonXVM/7TlXhWadw3
nIrSWfbPPOLMhJ/wfelB8cao0VETGhTu0F6jshjXqizPvGUhQ2m0B/RUFSPZCIyC
FtO052Mvn5BARpcu9gcBt/n5aGoSLyYfkq9Duh3sdxjZ9XDP0G9Ux1qJpJidD3gg
uCSwyPF1knN+Eu2UeHSeqip59QK0pH88nrVEP53O/5WDhZjY400vgrIRaGyC/Ai+
ws9X41CcyJSjRK1uT7CU75tpwgOnyv1ZujVsdFZQh4MJC2dRTFrZCo1rduGQm+JP
rwxbQnCqrcI37PEj0Q6LsvrQY//fqA7UXXq58scVHe7RDjgCvibcExRFXRHDrjSd
qYMtMAcTHLtlxdnmHCj2Kzx4TIWhBFpDnErOmTG7oO7QtHHJjoBh6MGqg3BQh3rt
o65+//UgpqqCh9uE7RdH2RzdOlhDpGkn8HK5YA8jhVZWj0dWu0QWsFAPGPqgxfoO
Dfz4Sr6j5Ig1Xj2VGpt2D7jXltwqB67j8uPb4ZzWvY/BvafwHo7xRHn8tssw8WDr
4+07SBCEIT2i3kUx75ODWiuA+FA+FS1GkLzNLsDcv9sLpPRogb3wOgCWigHEHZbZ
MQWuPRWrLVBfw79JCSMFd2d3yixEZj1J5CW/N3Gkr/RA5k96UDP73YMFXj4A6HXo
VwKN6b4CprtbHRjYAKJ8/oXYoaYmGdlKY5w5Wb+UfLZLuy1kKBFw70RMzBUJ2VVI
hg9Hks8Mtn/NopI+f8na7FyihXgx9CbY8FBFq1ImQScJ2oVPOSh9oBTPlumdk8d8
FTJUlfHblpeu5isUErlcekcaLurHUqoWS64pw6gfLKJ7IIto4DOApe0+5TSmvmqi
1b5566/pzu8ExdSMRF4YXQAaYq/yRcEssndiaY/vP8Rk+xkfqDt+TqpaB7ClZlPO
GXroADSzyP0PG1ew+kTogZioX4KWKJv0ysojnRqfV/QgzRoTHT3Yms18ys/iF62q
ZIdPtQv/RIVKc8bsmk7gUfb82F59yXVN4q/pdZiyju9X2cA6JwFn+Pg9zeR4mKe/
ir52tD2ZBNzUNo5gHXBkyIW8dJZNnbDVin6z08VL3j0oWmlOs38HMQMKC1PSvqmW
0dt0YEIL+qRlV7+mGzFd5CM9o3ycMMQ/1MxrE444xsJcQRt5PMsiiaweC3NGs6hn
fZzS0YB2UnLCrgxfMTj0Lex3ppRF/PrBv5Oi+ohOzbI99oWWu+STKIKMzo40GsZy
9sjDzZb8Z8vs6D1jk8VPDdqZDdg4soo3bjxD7Y8E9xA94Pite1rFyVl79b3j3Kzd
xBHPFMRgQBz/foWZMGDy5ZLPjJEunRKiSy1ybaqp1hIEpjCiMs3NKARYLZ9FKmIG
zZq0bdG1wIehIeAN7duuv8EJFzM4OOio5+uvYwLqKBpj79c6rUTtbKw3Zg4E2RIR
XOHaggmHW22cL0cPiWxdaUf4NP9WRrf4VghNNlVNRWRX85J9ML3pq9kFWpyP5eSq
ho2t0U7IOxQhhSDaRmRWuTS1zjtMQEco0wSQ+plDj4o1xgWQ7IYQuzkO+AKWwipK
W2InfxYgtHxpLlnOsXyH8U5b57dHWIOPxqJ6luVgHsYeJ+drrXrK8UuVJCVi6A5l
aFkJILxXG+9dUSnNomNNfk3aY/qNKx3OhGubxIZM8ZjdRflF/agrz4O9dAO7gl30
j3gUIY2dKoS+WypjBzP8saGj7RotiGb02Lb0BIm/6s3FcLt6GjtAtSI450+1PuKl
iaGuASjxpt1BEmq6y8jIoaqkg+4xXkVGhOhi0BqIY05Gx/35nCdATWHsYI6uJBc+
bKUJOelPEW7at+LmQXwIW9t7rpqjDEhAUMuk9P9mmE5NjcFy1gkfd+vak4G1GGAv
FzrA32D+pT8LK6VJwkKK+uAvCExj3LzCyp73axGjk1syLHEB222UUQd+Na1eJVlj
fwUYx4LXF111I6L2bCStiGXF3tL2O+7yk87fb5+Ubux5tFKJpwH78K/ZZAnQ4NiA
e5mjE79WFO4ZLrhxrDy0dGiEKcE8sXFc588qNf/gllvE9ANC39E6Rcihy4t7FEeR
xnQJmoF6T+RWoy6cGIOiS9A5SogEDKt95abj9smOj7nFqos9k1xHFqICpoS7K0Dv
bmnN+byzSpN4ybhOAVMzV1J9Aw+r5LlHIEfVOD/veCo1pHL+HGhGC//f+qpEpGRh
YgbQGGSxmCnyVMJ+mR8+GKHEDfjoi0IGE5oAw3G8pVbEUkmY71QE6mbMO6K9GKbQ
XGcM0J9RSGNT4+oHfUxfCZa2i+dAyYY3/Der+XP2LxjOfFrBSJeuZllBzYSFSNnd
k2BaH4118GvRdbjla382L+pWgSitVuDMO8hgX4kVLWFcy9wHxdYFEoyp8G1Tt6lb
FGypFP/pVzLaNiHK1AyBOFJTQLXxnPFsXlGEYqIrtFpGiC25omgCniaZd8zQZx2j
j5s6ny0UjuvO5yR2LXfrk11hxMA0if6W4FJNP2r8/qu/YdHcJacLw8tX2z40hUbf
uXq00PToaUFurTriuVT/2suuXNHhjWWz7aEFXZ8P2uzzaaKpVnpR4BXITHU51/nT
pd7R++CaVQbH3YsoMarclr6wazYFFdSH6w0p0hfPFDACaS81TiGDMANq0BZBmpWa
bkhZpZ3aGIOh+tPiZbfFSy7ouj+LRuKQAZ5lbkrlr22kbBlJFlB+JE1BHoeeRh+w
xKRlUpHohA/oc+tdWDs9vu6+9OoeB6pJQ6RvNvVamlvh3Nw0djJskwzOM8gwA2XO
lfXB8yWarR4r52zZ3v22fr/fyF5Y2PwFpFvmKGM+Nr8+4hkXY5QcylD2NjqhC4zF
Oo0vMGsAdZT3kIldt9/W2df8wCDclXDmxmv68ikNqOzmZHppojeGLiHxuh3EbEtc
WyplOsI/I5w+zxYw2GyOd9kCHnRqxRLfHyRd8EznLzxrH5vTMq42IGRW1HUZG6If
viLcalD3RpXwYiILj90FEgfqR2sLsVstHhpzeSzAnhM6/BAyk26fwRQ80ajIt0t7
FMuwW5nI8bZ3zFWl0/UXdd+ENLVDy3oaSpBjLMC9kXh7ore0b/eGwGoYEXK7cVmr
DNQc20el+JHL2Mv+/O7Mqk2q51hjnfYxbwcs8KoC4KQH12UugS+fYTUTJd9fwW8t
wvUyrp6GtINEdKD8SB2XdEziuV+UbT/ZtVnBveEnfC6zB6EaHo4qipq1yPO+pCKp
19/yxS9/6ryNGWlpGEd2U0mPQ62mQEvOtGo9mjnEFuS+xBCUNRGLSVO9uKtPs418
pWjVpgObgRJMqVV6riCj5Qkpn1+0qPNO6F6PNyqOoMAA/StZqrVH+SBWWIu4k4yy
01jHU5bZT7nqLKQ0G2ukERe6KZzOv7XYaKdO2+i6dIpU1VQ4ZP9J6dQxzBGAePkC
Ywjg9JbzVSaqH5FsV6H4GAQoGBHpcCzSrYFsxRKZIojKvzqb127BDDqgVjoGB85x
7sNggHCp9qjqz41Eao5juPLkR8aIvEhpmmbGQvwfh3l23PNPOk4e6JUPELxI1f5/
uHURl5RRlh0fhO8dEUmBcd9rGPJnTTo1+cUHG8F+Gnbbw7qAqC2aYUVoYaadPRlX
NsJRkE5emQWHVXi9hRdj/3fctQgRBCyNv97OpFmiC1rcwQzCj1f9astyTadZWo/r
LGGp9e51II7pDBurdDsj2nB5pQVdmfd0z0Vl3SZJM1PZihomXHqQR3plgbblM4E8
JfuE+ZwNrX8OZC3pkAvXH/opDdlmYR89mGJ8rRRzLAVtlSCq4wm38aGRhlbduwGa
OrPjCn3Yp9MsfVQs3nYa2pu5T1geNF8/pokp+r3e2P9QMCnyGuX6hDAYWA/8my9e
zTeisyBMn/HRld0P104P7COt6fO509/vdpSbQFw/44VsxuV48OBosVsXBUyzyY7t
vWr28xfpFnXevM9HkLuRpE9D1005qPBN46CBLfG20eqIjKWNbmzfuC3aQJ/XcsOl
NbxQQKtYPpekeY48IduH4Ue/YCSuFqnEdrtPqlAmC5FYE7oOOaxLYbymJ/SLR02I
Y5EeTaGiYyqv8gRz2JM176y1zrWblCswlBbDnwidh+ZZSmPZC8d7/KYKoWJrThS2
HREQApQHv9FNOAhfnHrUz035DULRZ8d0l1QpQSx5CMqBFtQMlk+ykMuiOmDwKrv7
AZRx68S3GdiccUdXpfzLVfR2DO+Gb4sikW5DDPIHvU2dGC38shiqJ+bT0EPPV77O
Qrhlhe6GHnNRStTmeJxzuWqEgTyj+f/luGqDtaIb2jDFo9ezJD1Kk9II+bhB9qpK
92pGhPBaKSlABVnVPOsI1f85Poz2H/CD1hcDqIoVsU8mf2txhkFxDrCKBJBsrNbD
aFE8oJD5kG6NkM458HIjMxOFDV1IEQt8VZuYWOpDvcQHYB0mkwajLe2Nv1lmi6LQ
b66jXiPJeaiWyFle6Uh7KTv6cSxap2SRfHnVshQB1m9TzRJpLXousLRm34G7hW+j
2E2bP8NuIToUOB3FiPP5cwsOfREGtt2sbhWLtwgLupVW4T+Z4LhV0sdYQSChnaU6
nIMIXxtehq1XZcokxOwMuwC+JRPeX5mBcAL6uoMkNkc5VRHvjg7ay/b8f3xf0FXN
nyoy0vN0jSCEufIjAN3PChddsxtK/Pjrl8RmgD8OF2rw3h3uPYqAZ4ZReJDqcQvd
xCmfgGJQ2VvRnOoqBRbAFzXfD8nVwxPrDwxL1m0gVp0+FzolRsF7oWaF0lOIUUYD
NnAFeGabKuHMG8D2vpNPV/3Obb96sCRzp9DGtvQWkqgMuYhA89mANxFNrBwyD9Uj
EbIYoQSx83rPH0k4ZuAt+I5o2XQ4kkaJDqIpujnVYP3ajqYCBWDjJdj4zVEnMH6K
dOhB45d9SJ1PZU7lfk2srqCBXxYzIUIPyRya+Y0mgjPP5gjHtfcDUzxdpYlDfSzI
OZyvHC8M9T37vSEpxjFod8uKhiC36R4Wu63C9SaWJ+kfJrZcdj+cocLX5ONeYJD6
BYA1Qsubd+kdR3Fc4DvSUe5oo8S5o5DNt05DfZWAOHiL+98xw18+59LsNv4W1tNm
2i/PKEzVJHE676DGJFdrT//XxiYJVYgCDSdS/vZO9C11lFSBceCf1ejL5GjJqd9k
z0fbi9y1w8mZ4iN5Bl/5Ec40RDEgjn/sV4SylwA7ezzgpiIvaKjaAtAtnp2HqrVB
jRMh6T4O7o6HKRm8t0GkX/TQGs0oqIUMJaLoQ9gEedZ5E7Oi9TgF6h6/AMU99jY4
tg1MD5bBQCiUYlLoxSpyDeCMLB/tqkuwqTuSuNpVXo+c8+D3TOqpMBrVDEBlEcly
+wk+p2VwwQxXJopzlD+Cn5VlbYUQIbb7VzQQNtMeW/LHC3gaJcD+HeBNPxcO5TSE
y3Y60SVlrEzwW2C3cZehK+jU/KDlB0ymDczHeiTHq1ulHVyZp6GF9J74pEVHBQpS
KAKRFWanAkWyqzT+18QIH5PMJs2YaJzROL6bIJm7MBTWqNH2qn106jhLn5WEj/Sy
cjhiak7Gsc4MLbTlztzEO9dwq4DcUIpHvvqeZyo5YdAciWdTm0+UKhiyMJLH05g1
mvcDo88Do8Q2fg7oe6jne+uSifiC2QiplFI9N+gzuwcO8qv5fHasqK0/SgqtiA15
MHZr+wo5/7vptLviRovdl+WUnDZp+vlT4umRWhfyWoL6Tz/Kl2ANkyIzmRy6kooE
5Fj2pbCq7JhS0ySX/23bBwtVNpKebkfYGlJ3/IDtCrfL3vU5ChLaM3L2Rd2EzU2y
lxPfNRMzDefXPaYcpZvC0Vbwi2ce4IsBkq+IoZxepUR+AV79hLn4KwWget9f8HAT
j1OPrcD25CZhOzQFlyGTV3s3xhpRlcxALA28vHitPLDTbuiNwvGaw1MJj3wcY6dQ
BS1rRpKjShIm71MGU/G5NSuFIuMRpYuLFiYd/cGc70jE3McqZZcFD+5RgX+dFX26
gbt6Paret5t6nPLv+4i04wNC7YzMT4QDFUYzRE05c7sB6/XYAKzLfedNb+ENP7sR
BZ1rs9qcU32PtNFB6EXHPi5i3pqJQ4OrngaI1kV9lathg04PMYGUnnw8IOhT/M47
3r4l8OZHmwFECH6rVO+lQ1BpAza8P9qAXr/+6xk3+2sgmrndpUvZGoOlMYs7CkWr
uqTvaz8HFMjbzm1Pr6JwY/lvg6lHLrfU+4Q5Kj9R3GLpA/iyq4HXo1KIV9icIrM7
+xDA2DnujaLZ2VTfhanOVFTdJAFTDpWW+dpaKXiAlIaBlSxk5v9+D115rMauYmEB
Mzgu+Ubt7TeUPttQ0cN0REdTAsEvUJ4uoIj5OdhBrpmgChdo0cJ5lXS9APj5ieBF
omhLnlClV6DfQ6czSOjzQmqfcWJhn2gShuRM7TPQEdxBgMu78IEz1Q25tHFjUNws
DkogAtK+JGa5JW1e5LS8Tg9bHg5JVWGGHeAOsSlaPK5nPoiSX7K/rRRaiZXV4iaJ
OROoh7FpzcseroTZsHlt/du7TxH9ITZFHl3u4Wg8SDn5ie2v61MXRN4pcqdWxQWJ
HlWWLiE6jFPMHIPujrptJ2v2Mah25a6ch1+HtSu6wfCi4BuyEsD19mMqRc7ZvajQ
Omz01W891/6187ygdT6Of0JC+or7qhpBd3l8a0xSMRbAkbjNxk4ScnMAMGvTMEti
6DFLdZszn3q8sCaSOcOcCThYWjeC15vQcMvhxzanhrYvAx2EIPtmOJRyMQNnV55u
qDjpxoxADToEjf7jFSitj3R9HDihouMQWTaRIfr8R/RuzulC6UiALFM8vHz91MMU
0CxtqJZUuKXipWkF68RbYrnQay+NumsmORxDQQfubT2nqOeOWM2C5VFelORdXD8/
VZCI9iofI6LKmfyM9VkOSG6oNZB16jpM62pMUSqoW3kWotSIZBsOtXKshaMpjOSZ
goO6M7x3K5JPwCESyN2F3MQ9VKTSLA13mpQIrOLYBCYXoymYvf+XApiR3b5EItVy
WEH1bER680KA6Ni3zz9WQ6AVuCamPhoeftjd3gjulh104PELsPoC/gL+ZlASnoWV
l251FiWLHFxWcaL++9g+AcOBJ9nm6zujzaI0ivS+SobivDPA7VV+4R4ZKemff83C
oQNoeJleiOgIr60zN0CTemZT5p4TredvpkQ1sxolVHzUyiBVzug4ZBKEKDAEvtea
QGhJGtUyCvdqPW8h32FzkH2qAt/7QysGlPWslC89PD7/LqaurSd2jsxzX866dBoT
WbuMcCZYMvA/Hbqw5jcq5I2Q5qaYIVMBXa0O+ql7VUIQNrr25rn2glMCIIJE3Va0
uftn+MC122FbTao9lu2EjHzFGTd3w+opsyJVaVABYFWnN+JX5sbJKYPm0ASlFpCi
KMCLa/m8wmhkubw7S6PXIviNw0SCBHDE+rczHZF8pdOWgu47easYkrxsapj3yTlV
Em5YEd79pySh9LukmSZ8ZhLTkjTWKL32MyquyfXUy+3xVExVhtJIR35q/ySFANvn
1uX83x3Mhvk0lsAQSjPOrDllPDpuluKSW9WowVsnQnflotmlCT8duzjouY7LBifi
wdqAbilLx0N2lpXN/dZ3O5Y0OeoEAUwOI9+KO/7VcFU9CaRVLpl9dvAaAsYXpCly
RkaRczsR7WcnQOywDNxVTFfbxHJX0FvP07uzcvmwc4Z2RS0SZhnzu6zf8U8kxPbx
fnvullfU21sudqefsFpUvX3m9cKBPkS9J4cksGAc4wc5nadbavAgMJ0DFfhvqVcn
lr+l+DZx9n9SaF7PovAsdY2XL4WhHKbg44UyfviwDSHeSv/PExrzxWhLViyLsZN8
9lar5AqS5A7/gvdB6hv4b6L4RPp5fvwUTLC0GONFYPep5B/bc0cWQC7CpSKdhUkM
x1giHlY4svVPhyVix6KzIlho8z0T6cHE4lPtiZvImXRDswwsQ9iFkICJomRPW9hD
lBngIMHL7DBDEgxLEs8G+RlgAONMZBdPJpftsB9oA9WnTeY107QLqIKvycL2w3S8
HOWXVOslnWlBlPJVvOV5ZHnx6HbvO6ovVLF6aT/w3E0PLxPBO557+cF8avYeeqMf
uHvJBvX60OxZ5VbDOj9WlBpLtw8Y3Pjb9ySQXH3NfEJn34tOj8g2qjtVnh4pCegz
Fdokr5Tp22sD765SG6tq8pquhWrl1dsWRIJeSxtToGQ52Uxbm1D51FmYIdh0x62R
spPHAbMTfVBhoCalyT2thaIlEQs34Tn/n/oTv06qQSabxGRxcsDglPtMZm8pPrwx
k+QysW1HBD+Tpdcd/a59WvJCX+aACjvExO7JwbZLdu/wE1RpohM/0Yjd7KghtmjN
kkhjRMbWO9iBP0ivkXP1J3BNIuyaTNCME5QUnO2IjR2M16pH/3Kz5QpLo+8599k8
Hvo6niN5wl4zumvh1Tfq0Ra8gppXVptyDJsQmaueKe9fKMpGMfDiuYMsZBrfLlHf
Z7joVV6nOSZDZFpaZTKm8KHE0XXkXZM0rj/G/4cc9KtmcNAGvnV9NO0/kQtfvc4D
mUj/tFY28RhhdcjQwBNhx5s1anEhvrsowR6WbeaYKkIkTFcPWwbK7Obi0jfISYrk
F7/shZivhOAw7QPbpt2O6T5j7b2D2M66r4/4wcnVj5hiPiCtKfGw0pnrMaJ8Wt6y
iGOUPuOnJNKFz+4aK6Lr36agACwlsoHRwDyoQL+u0iY/mRnnu98tL1f43ELIVzqB
x6dK5soufYk9kHQXgMffleE8LPRkDCk2/PqHNMp9iAIJiRtzj0IHGRQyWNaeLXLn
wJccvI+vZA0h71pgy6jMgTmc7Wxh1rerxi9OgKkIkqOCxqKEq1rTtyEm93mAjKJs
7wQZlPDmUGwkbWyNeTtPzPaiVPEIclFEaHxJ8qAeFcRfsMWdtQQxkWyRrqAd+W01
Onlfvfwu0e61VmgbFP/DMwVjU1b5t0cpX/FH+peiFYNPHLD3DdpDuMSFrPKOaFtW
e9DT9S1qXjA99JJajHz7G32EJPf7NcN+2yys85kvkSBmS3X7lOj0P/ZGpM/cNZY5
6u2gTM3FS+TRSztUAPrDJHOT4NP/3nMyJpAFhbboC+ioAD32L+KMfri+VzWX1RKn
ff29nt9sW93nz3uyc5coxOD7+vIWsp8gokcYuHcBAN8z1munk8iIE5qX5ajMFV5y
Qa2QLLVT5wRk/baaXoJgYNhUBIBor0eAim6LEevTAWw6g2FO9uhMvxgsy3dgAqVc
80HEHRhXM5ZTHS9dvHCj90y3cre579k0Xn9X7AOHdCcyvLpYhpC6isWJjvpB+/2q
VEY+CqVjWJQ3CxJPsCih+8Dlgoc8YdFHCL+KN142BSW+h4uvQHUqeekcSQ111xcr
TXPF4p1H/OuG1SU1DQ2CAEX+fvfd6T7Mt47RvIVxDLaUXlX/N5Mzhhp1iYQvs59Q
el05z115yg89/95DA1EruedI3sqTwRxqNSs6YaINhrKWhYCdAP9wOCMEpT4J9KpT
82bC9u0BLvpRaUipRjrc7B0H1Jlr7K23WfNJ4fNCWpdwlvZtttIUjUf0Sr5hm/NR
0lT++6Xk61kUMXF8zHOYDtD6xL27Mje68wZ8MSphoT/thbJXsGt00Kjdxh5wYcmu
xv7aO4YfBvx+i4hDgVfK/f4hhbGLcxNZrTL9gF/nODVeV3/89mx4PF0KYe3/FN5I
pnSwDwMMML4glUtRQdLHsnLm/oHuBaGmo7RguiMEO//YIHM6tIZPzG+7MPfQ4Yg9
9IEOygDsaAQxtkclGOl8k1GNW0M8CIKOK3u0r+jLBpI7P3ov1Z67ZAGQ5yokZfAV
R763iuCf6hJzAaia/L5HFGF6ziMRGmANv+zCgp/HMuSmYCnowJJ9/T+oJvkzkD2K
rVnrc/0Gpb1qrFNJ6Gjp+LdmBMRfzOpl91JnbJNEyDyph+udy3Ut8fPWJaoUYwqU
VWfXSF4urwhCETVMKzJ8E6zzN+TLg4BQaoM+fgD4MGeqkGn9dm5jyKSRkTKvhiG2
q1Lkf6ryRUu8jw/bCM1coX4Ndjlk1/7Je9y/h7Grw4IAighMKHxEJFN/vNYbYG4T
wwYGdwDiqwdLbeLmCVd6IkBsWmud5lW2jiTWfMOf1/BxA5PX9d26VrpKc4jnpkhn
d19RuaQ2RKHfK+4NgL9H7Lw3wKYsYW6cju6nrILX5OqgHDVD4R994Z8dTJ9G0Lhy
Pw4S17UOZf1JnGCmUeHOWVAmzuLIyMMnXa09JMp86+sjbMcoD7ca0KXLVUs23KTk
9Cl9q39L+DX2Rvu0Hq0Gqw6D1EmAusllKvlQQFZBakl/yUjJrktewm/jfBzYyu8j
mtzhgehVbjupzReTUGlRHLk/eVx3DUPdCKHOAzdZ9e5qNyB3NnoIConMm++++LIf
H2JEk94GkHXwmaDMvoqq6PyCDeXQCHtn/10fMrIRqzB9lqrjiSDfaxwdEf6hArD5
lNkK7r8ymJU8JnY4Ni1dQ5pguSY6iZeasW4VWGLEVyvB23+f2sKGz4XspVl0LK6N
UtRJVGNnVN7tII9HfsOYHuYkoraH2nRTLl/lEeiq9fE+5r1wQYQjYBAUqWp6k76I
H4BwI5x9QWcpyf19mKhJGr/8HggdnxBGfSJrm9IeEZ1wZjsPE9xNR5kVbiQA5PW6
0v/pQrm6pkTHF+0XKQiiG/q0SrdahPAO08gjzUl+WVinmL+7VYu+Pfk4ze0QHZCD
H/QLBIidTGZedqHNgrN2pzg/otrj2MmIAsFSNo7rBEV+jELj23FRb292f0f36n60
k/RnNPBRfjPhikZale9iJ75hRib3WVhd25KC3BDrZYOhiKEW87kR59gIfWRUUEMi
vOljE4vnsgyflxXIdwjR7KEmNLEY2fLRABMb0GqgGathUTW2FT50dEcKeS46dZ9s
EtHmylmsWB7cEIlmU3C3hWfEp9S6tQCBu7YEk6H+fjq4d+dOOXsZAQDwr72PlHJ+
OdREbqrzk9SIspgzQP/ot5MGiYmUEeYtaKUd4hjNSI8WanQk/BWdvtEtdlxisb30
3SFDOFaBZLrRrgUGE8wLTIQ+t09iw/HdM8KYMtuxLJDgYBI0wgsnaUeqw68dF2Ko
DHVMkKdKHsul8/I9trNSeaolco7GlboHMLmUtP3/LBZc1aMlm2P20MlD1GtcLvp5
Uaf6R9kkCCiN2q6AwlUlxqnqs5lWQRHbmeDrxBVLzNPYpz+68LWjjX8XyJAZXaOk
TCAljbCmDb73+uATcI4TdOm0DXhJtAya9awLbqh42Ydb/O0gHkTRoz61c0THtxhU
GYLaiIw90m2IFDblYrPuIweG3NUR4sBK3FAMrQLHk0VZBiEJY5z2lE+W7zP6PLSF
SlYZ0HQ8qfzoZ/wET06K7xOGTYvUrVQEbS9QVLUkpHbT6qsQ3Ez5MyT/G/AinQE7
qbzIIMmUnU7poN64NPnS3p1ul3uWbCAo4lvQvKK89RJEGtmk2dNQO1sb88pCJYCi
vRQ+ZNdFpVGNRb94o8FS0oWjrErwirJZZJ6anXQirQNbCI74Hie9phFQaCPFbB6r
souPQo5IcnB/eLv5x1rJhFBfcFV6e1gaRzPsLsGkZMYU6psJvLfPyxK2G90BNSAa
uluHT2WcwyGVhiP5+dWibglXas4JRIRAukpWOFiUNwXfsK8f9FDZ5HHUTiRyLC57
+cvwkFxH/wwjMr6V/nZV6jZ6PP7hmrVitelgWpeesDQnJGX7i5a16UV33JixfyrH
CJKKZjPmTbkh0xemATRnifbqeTkGgE87HkckYVMofIRQ547WXvA1iC0R6RmaJfRA
ictcvDSrGDawqOkHBqK7hElxjNeP/tbvVVLSFQHms6d9l3YVqI82Db8fSSNuPyQA
3wFjNO7SBuA8x3H7yciOZ9+aBmrlUy6bJyyedqe5M2/Pzzd7aymWAcQdmjKj1P0I
NbDPzYpRgTCP/25FVqLu9Uc5LbedfdV4/BWbzcMddrqpumNWHMfoxrJUtBz+uDnl
WnZN0DvuGOKj4tJMrp73FRKtM+Z4/oPyNU+h+Ho02K9KWcmVElAexuq4pzQnYEgC
isMFno050/9IbDw29SWESw3OZ0W4EfCCCqmwITkdLd/uMOBnMToeNpBSvh338XbE
9hCnb1WMmK3ke0WMER8yM+PuRqN8jCNUZ1kCNhDO/DvZbkNMAx47ZT29t3N7ffIR
Pwfp3QwExJs7l6CkId1G6Z+z5VY6oRIBxDvcBCsvrxGYHlhcBGyw0vv6EgzEWhC4
1BwqLh9SFUeIa/6V3tWhaZJr5VE2RzxoU/iQLFzzC43mQfGkaHPxDqtGIj+O8STu
aW4dXe/w44Zh5PO/2MKiGX/UJa7Q05zm9oTgUaQFsCyfXvFdnWISmERp6scOFt+j
dQlg90yPu8jv0atmVjH/94UBR3GWnpmezt8EzrhA2+9e5Bvn6jYQ1IOKDwcSpoOq
ZFcRDFkTJG8UwyKgoY81uq4N1ahuBg4d4Ia1EmuRV/POaMDFtzrMhjUDAaUe2Nni
6F/gRRvxteKBqytictrHYgrf8l/RItYIosx7QsbBFf04MFT408sbrDNH9ROrXOOC
mftBCas54n+PfgMC/cwESmfuR+z705MLeVpaIhht+473Ehfl91rkkt0JbWql90+r
KE+N8OsUBNKGhKzSfQYvI/0COj0wJegKFbG9aH1K7GqXqhZzQVx6mw9Te2Su4YB4
POPU3zA8PM1Hqr4QQxTWJ2KhHuAdCl7+6EDscJwgHVcyNtjUwZdEVQ0a6CRVTWKy
EwDt1oh3sJ0+3NVLo9bGX2fC5lzsa4H8d8qWZPvmmy7ZS8/pb0tYAGZQ3zzoUrJ7
hs9OngvZ/0l0Oi3htjD6BnhuRUE6ViqnqDKv/36aEQOV0XDmOF4rgil0yPtJQ1zW
yGKw6Yp2c9XZHmppwl/f+OcceuEcGm/yFwCO9A3NczogveC7Ly/N9ILQaK9V0RCw
uTuGqomNbADB8+Xdr32DXEudct+W5LnRVK3ZcBAuX8Z2MFYCg8YmSBojBQVgE56e
fc4NOQ+N1NJbzEBc9QPJxTBX6aecN9xE/a8QnV7f4tPEO11qGz7S7b9k36d3cUfm
TayYNUHgUU9A/a4C0S6Jj1u1YBXr/nIog1qo4NJ6kuQk2nDpnojb2+iWP+VqvK5V
s1wMlOphloEY9pWEsdNpLM9s1Y/EFqa6QroIGk+v5LMzKHep+0j/1d5Otei+IIvS
zuMd+cl5h0Go2MBJoH+b3lWd1M5AnBibV91ogku7ezTPgc0WhCyA8sVKqVL8NMl2
HuTMGJ9SJjyypnLEQPQIIFmKdEXoOALQ0c2fZY0/fFdSsGBjv0J18PaD9qwvX9Iq
/TLplgpuZHMzT63NrepxevLBbk9OJmbRNUB8exmbfeCtAXfKYjyv3799oquDhFAT
vkOr70V//Unf1Fw6NmQhVjaALrA3OKpuPlJVcYxoPSlRpLIi1jyCOti1huFwWnh5
3JrSEu39+WDm02pt8bcGOvqOEgQ5XxgDWWEhVWNmNmtaYaqWd5kd7OqkJKHFVzLP
XLs9dWiEjGBM2znHZDWpam6jsWmEst9vu3tqnSz+weazYmst49mdRyf+DAasXcpD
I6UkKxP56KLxGpIABChYaqeNEJ6zsqwdbNI9XCQU/qFdlB7ua9l2MH2ggtfq1pvs
+gfLmgX5Voo4OJG/Z/PfcpvG4pKbR5dOPzNEJD9vFd2bpbDQXQ0Yr/s7V8feSE/j
5VImCdpEmqODkshrzYLaKVmCAHIdL7ewQhNJak3BG51faALDz2aLasaW8xN3Mo0Q
ZOc802LE0eK2Fp6YYOSs6ALaAkj7VBbUR1dqkf5/8yQgvlin9PHWBmJR8SQezn50
CuMQblSfhOAXv+oDzT/AmQO1yXOdKBSo5DNjisALid/MZSNTfjHfHEuDfXQBNrGh
BruX2jr7VdqpJ1jfSSY5DxTfFNo/pOPe/4Bm8a/MW8F5TiVkYOo8E2HcRiugmlQi
BYnq0L/OiFw3qmvmwYRpX00Mn234fP64ceklgYw9XKMYoHsZJgK/cjEM+mv334Hd
PONBUMKgHEfBrM7JdjEZHoKYD4NHuYGXPlCavYF0ySc2HFLEZaTMiuMDMNHlpf0w
cK6tUtZ8lL5WKdPeOe45w2m2KusGzcg1IbkECLLc6Gz+ScE5aiet1VoPjVmWDfsg
mEHZY5ePeZo20AJfx+i6ETfRnrnvYsJhcg/ijwShy1fTexIAYjPiWuIBuMiLNgvh
tZobcjaAFFFvISaR/6AOypa795v4FOELZUnCDXeJp/cdbqRYrz70BJNdlXHUG64L
h8N1zCvcEyKv927hzzOG8tyUYgzMrkQhIw612r7k3qcYh96uKAUzof75K6pzQ+tf
Wh6Qs5Qd/YeE/O60MHRQOxBflUOuVbqZs7jChhbgoqk8Q65kfCi7oaqWxNy37cVK
SYahQCtnb1PysonaWKvILfyVAmLCZYMz91JnG8oL7eJ2hHWZUr0P7uhXzwjL0b4p
Q0K62Zc4RFqOZRm4i27CMQ6tb2FvRBC6EW6W/uk3Fz6WyHxrG6uTLhfpyHYTu+A8
opXh11uwlWhqnJ9DCMOfurDGSpF00VUrkOQz5eHC9ZRmxn1G75Bgzzld+SVTK66M
7Oc/uHaH6aI3OhbynkoIOZx5n3rR5BDob/uRCOCEo9tHKs7SvrH0CurT6AGDc/mM
Cc0E48S8czytCK0WGgU19Gz3wu/h0l7qharRC2JYLILoMLuszyGtxTYxPq6Gg4HZ
4fFOtXFEATTkFc83VRIOBdope/ucwJCDCigdUCQyKlC0CarnPyrGnvuB/T7AWUo/
VFcOhBDgpCg+H2g5QL+MZxJ9n3uOD3plGVuGlU+EPRfU6a/Q/M1ab8kEgjC0VgXI
tFetN35aAQ8Nhv0lHqeb3n5RDUueFtmq3KNg8GcCOm/xbthj88BArdgGwTnW9OdA
sYJ8nCk5IpvNB46OS+LxLEI60dOQnykpn2sw1A6OtakxaF9j4R0YJZ+w4Varszp2
8OxLepCC26XoUWMMeivoorxWRfEPX5QMLMCOLrqatCkRuORQXzUH6LpbR0jTGUze
sGPi1HdNcrtcHT6sYBA2R1MpOuF3cOox69Z26NumM1c4iNpEIPEQ1UwATQ0pNe7D
y8Oph0RXKAj9D37dbeKFks4U+6xBijwjTv08u1nFxw2vGdpb6NymjfESLAKxd7Vu
iSy7+tJCqIFOwnHQRWf1JR9+sH5DS5g0ZzoiT5vYzIJCRJjaK3TYK6qcX7xBZNmr
YlT3qdc9mvC2qs4h0HWDosK/ZvZd3IbrAm9/bIe7utoOPatVz7R+mTUKJbFxJnDx
xMfQLGLEMTGjG3Rqs6Alj/RxHYlr9Tf94/6M0htZFljEJoGseqZt/x2zNMrOF/M3
6tZDHI6BpTOoFEv5w4+lZUXaOuY/wTlbRsMDiLyhzH4K8HFD6iSwNfy6bC4BAnuW
InDJHVmJqR6HqzqYul1LrQ6e93Oc/uMLqeojkYQZEfyQhxdXNvrrMzO/IyeZRYUu
gRyXLqrydQIKC0VER/XPCSBmFNPrt8DqkRSq7fsAEnxjOhEXXGoiBQPQX45dU+7r
cYHV3VRfaOSfqbCxyDN+PaZuw8wEHSdNSyjRBqDpxx2YQqbTT7MAKDkfBC/IVzSj
D6VTS1w6LVNX2IRtYIVX2D4SfgdHpvzs54AS/TMttKe+CUT8LnRbEqLljyA5vFfC
2qLLwRUUeTtG/cNzOmdpUHkudlDWEVTaCT3Ubjql69u1LXTgrM/SrcdiWy3XFU3K
y7sQlbqoSKURlIuWVByVvrrvqQASVezXKX2pAdJiSfsYaM3GUPDDpCsJbnCeR8bZ
DUbJTuOBm/DDj996HI2BiGp+C40jJP2O9ENlq4FAFIk+gneccbS8acTJ1X4tYJkh
GQp3Ll23OElAoatp7Ll2JRpBLdN2sOdQpODMpPmHPNqiruYlChqJLLS+xa4z8wTg
uH4rGAqFVt3smzNBIoyTaaWcsadijtRtwAvj/3OVAXvtWc4LHxWCH+hijcyGRgTD
l6xONHNjiu+gwjJmarysjJIU2Ji8VVHeAcdUdZ/YM5BAAuxav4sOsm60S64P8Vjq
UC4B7pZJhvcar+q5kCt/3rQu0+bhRZqOQj4INz1hnTwPrtqNHnSRici6Srd2Td69
+zZWUWAxYIL5DdPpNskUmwfV7wXjmKduTiEvcg3Rdk5c8PJgpJoBwZf9VXORHWed
3iqprhpgviTRZtJ9D6bO4yrpuFf8czW5p0ecAjasYXGShHZDYRTSrojUsDJWLrlv
Q80c2DOC1C0eWlLNCvqFacy4Nr/AOucz1kkjphIfr2MUI/7r2RahIIbUzRoglXU/
I8okgh7UOqjiptdKYnz4DIfs8qyqN2Iuvvu68R7oevUE8bpSxXvcWeuRjtxoHcks
gAe5vP5hj34ywn753UHdjImzBaHK1K7pzwiKHmiDmYTIuU83IqkDYYLzE+e2Xzrs
3GppY56KlHYsaRM28k0OfBdJSl1Lj2ODv1ynxqwUn8njh1gTf00m8c6qbW7Zdy+h
eBxUkfk7w4dAbQch1ieSeH4rfnTI51Jb+4JGc9iZ3OQi3OU62aX8YaTT4MefDIIp
CYayFKY41VVVU/ATuYbVL9uP4XNNQzGcb0+lAiIgIB0rzMRN37n1YTAiq0T/xBKL
`protect END_PROTECTED
