`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FSKlsT8UHcJ9CdTMP3HZncfYlJf4JO03MxUv8dJyQq2DHwXl0iJI++2ITtCkABi6
PL6uxf5qjQM+n74Lqqc2EOHCPqgVTNlSpumAG9aDrain52/mIaJd2k3b+vX5Xfnx
fSeG4t5uIObBFhRllw5wqECwZJiEUYxYr8XCDVVSY+WBwu0Y2gDlHiYx+7k5sXv7
T+f3mwXxkYg0qx/wtuWwZz9sRNOVo0Sel/G8tgvDmiQnJiryfhqYMk8DGvOO/4Oj
3UEBHyOEdaDAzcp5X4IywRs6+KOM8cfLimo+wikRrxm+gPrDxm+shzNm1fBXylDY
xaf2a9UxyxpepSqItkBWhserWl2aGXOUXWsMbx0I4OM57fLoIMEskymi4JojE+TH
45qcNXQ+GT4vOmGzPjIPrCenmzPknSppHC3eFcC9tUoMCStcmtrMxm3U54h+fZr8
Ic1OX/l/LWOd1e0d/WGrQLjsqd0A8QDmnOIQIP3uglDj70HZJlJeNklAqCA3TL1e
U0cwpaKuCpmpoc99ebER9JIj4ngGTcvRr0XEo/p9FnD5ewQVb8iI0TwOW/JLIbYJ
a5pHEplZSkCe5TfCLpM/uMLpz3a+zPccUCsBIQg+TcspDeklrCeGEjEjvxs6MOaq
D/bYaI2DZBSSj+VefuISUCVuBx2woedkEYk6yhGhNEZNQebzLq0n1jEdIhxGLj10
xx/zCKnQ2ukzRZZm+u0ELs6TT1dFTK0GrcAMKYMC952YtuA0pFm2+eQXMZJr566x
u2p1LMKaYk0doBpPUilBaK3Yab0RFoZBdn02RFxKGncPn+UBVb6cFx5w1KG2IWLJ
N6gUkgWiPqPleSgtECkQRIjkPsay7GLM+Y+TGNSDG5D1qOIH7V8fTD+DREB8kT1N
npY3JvRTX3yLYvW+wDEFpvg0YDh0j+bGkfCWapQvhj7xX2N4uIsVOkcXZ2sgV0EX
HTPM0TouHxm5tmlBD2R4hBOjwwUw2NDjE+El54tqV4lJK/GGFtJ0ie9dnt3L4JH/
dbOFgEESD5+9ydupKDs0icqqwPf2cp78dnMLWFF4UQ1LZy5dvmWH0ngmgmEvyNkO
wiPMKdhCTtfgn/yQIL46o1agkGmn34KisSjEYwqZvsRZl3ds88Erb3Pw3GqqZ9uw
1XFJYzZNAbex2WnbFYGnX71EzoM1fwADBPZKIH2IziIG4pwb7SW4MfL+632S5uvh
BQXGJ2w3yl6b4ghr8vR5aHjpGElOR6Qz3xQ1GAY+qmGeYDtz6ZpoYct29PHQJmn+
bEZgQ38c34koe9meSvSycSyv/4ZXGf8c4WDBy4sRCy8jYwMHftAex5K8a5lPo0Ro
Z3v0/aPN5/ig15+1tf/XI0jH4mtd2awehPxeQlfsmyhrsflEPhKFtKP19FvtVBxi
UEkB9+XAkqYIN1AyRrWJ19Ha7KthdHMpxulE7iPpLcsY69X33EZLD7dNWaEwHhmH
BI9qaVi9LaDued62diZoaYnfT/wMc/5Xf/WaqxXKPdZamfDeMfjpm7PC7BVNA51L
vZf+NFMs0SLjBLO6mjal02I9PWsGpOi2PxRWqsWOQKhundd2ZKfdw7z35nh+fAQz
sJyTN3hpCbNaZgWZrdmIbSx7jQvnMNCfD5THpcItv8Opq9qDwlXYT1Y44T5z9EnQ
zZy++sFLUlvSpjPgKstUAfqvfYIClhmrZ4140O3UrqKTFFJkDL+2N8H+uw+AoEPy
G29X8/QizsDJqQbY47kfY0eqpvcaTQnJ+b+Y+XqXy3nKockKvxfAidHMS98rCh79
UzUrYuQZk3+0jjQ80M4CRG434uQD40/PBH8j2xind1fllS2Gf07Sh8Br2VQPCI+3
v6ew8XE8LENHKm09TO4w57RetB9k2bRxUACqq8y/sxiVrvrVnK/ekSWwEHeK9Cht
uTp4HlzLLZ9DzpkYNv4M5/o9sfovpr1kz+M0EVk+tGvEWkZoj28A6qQIEbbQjOog
z05nVGL9g37PIzWwybr0csLrlBrKh1hy8E9cvFq7NjpghOvndLwdNul99yEs+DN7
69T5iapQcycvzA6wCxR382Zm9OJ9zG0kicLhi73YWnqt0psY31p6r+ZxbmR/8Q8l
wGE5WvOvM7F0MknrKSz2T9Ompr3hMKt7nPuJHlfEhWPP1e0kU44iNlpEif1hX1dz
5UZsM+yOOYH94qln/Hw1Il9UNKEMt/9JSji80WnppJ24p5MkwKjnpeqEmOkN3wZv
u79Y/5JnBSTufUq1plBVnoNCugCmzAvY+c0wf7m/0BBJsNvEQlHd5fAoRfLx1pcF
/HotR56KjplRUGlXzcT8vvNugmbka2805R5tX6y2YRGG3Pa864RB/OSk0oqCVJEd
15hEooc3WcmCfxT/vZ5LL0IVPJXsTXFonJ8Xf9scVG5xTdOW9511enxMmlR4zAxL
NM6oxBxNT4144sGUWw/mmjs8hhihynxrt64SA4tm+iHO7ohXbjYHL/2oy47xTVyL
k2Ni7U5irYZLw+sJHbKSSnuMNwkyQidI9lN/qHvBc4pD/YfMo/eYpivR8NXxVnQd
tKt2NIQSq/mWtGmniecuPQYLTC7vYc+L5mYavYVkzRoZcuBUN79kmXjUZ2z7arYw
gG8Jbe9uCfIZA6XzViCvpaSJgpHR1ts8JiVkS4UGxo+qmKXBdZ0Q4wus48PBTuCO
C8NIZsag4wRwIkONsH7SBsRFpLBXwT3u9ZkQdcKOhd5u8I2eKssFI09kOcr2QEtx
7fx5dRD+2NjzlxIKNcvutht40YoGC17qesJEpCBgoG5yI1c4PPGTkvjY4iNHsvyj
tjik72/Z3Le4MPuJvWTOXxc3I/jD8Yoh/qGHVQ2iudPXpqgl7ELo+ZNjxTFGA4j5
xs3UmkVWxjAcIi9Num3hSlAFUhsrQp8D6IJw8mUcf8bE+BLNOOQGXFrevmYGs/6/
0Lbqi4eJzTGmhPDtZhKM7l1wAIIc8X5cgMytY0/D654zE15Nn+enRMriYPVgdPyW
ZcDypdJo0AJZpFjXt8P2lGGZuOUqvPCUSdo3rOkSs+BaJS0w4djzgzMhlzwyzmSY
iyD2uNn9vYMI8lTl51ar8YOjR6HG5Wt3hqCoPUFCAdxauAKBlKheg+XxG7p1j38L
xelks7oRW0bzfJG4T8xFM0NRQO0J42iFE3hpLUtP25l+ViP3q9ZhB4OXlD5bqTTC
/0UsoruwuCIC217VjmCEDTgs6Dn3N6r8UkEFN+wNeAD+YxFx6fspJVbf8/kc6HsR
ViIgUlj7W5b2S59uDkbusovMtxg4Ivw4HWB5WeDdkgx4oHMKrp81tTO7VSPqL/Ap
h7KxeyuBYEQXEqy1wy3TrSxMEDRpr55LPgpZbGv5EIoPrYtOJGoQR7HWWMOlSJ72
6YfAe/sD5SBqx6moheTLrAVgSMPhMD1KEm0sMclZ2JyR+YNM603B5bvDoXF//NwM
HHTc8kItkiG0OLmDy6t6loR3WHppnaZMFzNQ6YGnHk8GPJMt4E4pUGg09HCqPi4m
PBcuD+aDxq5TQ8SZUjun1vfUo2DLVmrmtlqLHQUrgD5OcQHZeQp+r45HfJTlfBwH
iC8BNHWfJuy7jxCM+9WFUarCbT8lmv9krQtT+8HtAzuzwqkbnAIWzBwSm3YlC80g
8kL0RtzcRJoo+wnqJYZQlvVw9gCn73FJoJdBoja2W4R1CdSFphU71cB9JZWLYOSK
0uNIdotzahP1vkBkzlcHIUF/xsmqhr3eJ4h83W0a6j5e5HjccQbF/W9MFXUvQKqV
QIih9YKzLKBup/958ozYOKdjGc/Kt5Bd8iPAi5Ot5GpBpPsTIWu4BuvkedN8IifC
0lbZaJm+eCTHSTfKeEAj+equYx2bFBPTCF3WivM8D86c33yd265Bn704OHerHR/k
FBXc7Bf/tWgzE0i+0SBeu0E3dbCfbiUDdaMsZB08tc2ak/ei5Cq0XBrQpG8uPMRA
rUrVlsa80H1eTV0OdrDjOBYx3BZ/3ubJzbmYRPmrAltcgYu06dWTQv7JRQvHza7x
tPmFMj/a4DE3REHttb1vN38/EQ69fjU4vLhOPiksomWqKbM62CvHn4cSdKkpiYQk
2HuVqa7dLXd9+3bcadsIUvDOf3IsHmpJV5toZdFVCEBBII4N4uMvGfOCgcFKmQEg
f3b01iLq3Oh6CPxszDkLNAqP0s2uh73nZi4UdQJRE8+fPxF5bMUxIFRKgTPA89ep
YzKhc8wvEgbVLIV68S/7rads/5nDawrM+YpXNMFMLx7mTMOpsIqLMXUB5UGWiDSc
w4KDZj7tuXp56vikLU1OQUFBZ1YgEKfeWo/s9OKRTzwc37o26JKXXkLXFViIZUiG
te/mE8fe1AR05dVeuJkXdxWAnnClTTePcDmuEpfFBN81xT2w2lJwW8d+17mdii7P
uMkj4qAiciKupW77bI+1Z9hD8BzbJvWTARXLMNWIR1jvt01YW5VqcwGC6EUQ3KwC
nOGwuUTSdwVuy8ElMFj4o2qaIg+nWFsrgElgkqoiHLIughKL+pRkVsx/VJwFy823
vp7QiTKyackRPOo4l4X+Xx1I+yMPB1b1ZTEo5p+EQn605N9PlD77CX6c/ke3x+JN
ueCndwbLhz4Ox8lr+9EcxvmqA68o9QsEoyFWRqa2tG+WVlE1Aw0hy7AI6+1Haw13
xKTZ5djGrtkfEc58LMbAW0M6xGJ+JVymhVGGQjMjNwWUJy6JbfaCZWHqkfaKFDmX
V/IA3/b3aOoLhURS+NewGySJS6bwmxq5Czl1pKgfncr8TqZy4LGVw/pxonJDLmoE
PHsfJlfYSCO+DVxP5oJcNEvmDJIZTJX7c8H+eH/j7XMSP1P7xGgv2rjHEioUs24j
HbDOhm0c4jd23JB/XfL/zZ8atkxtm1NmjlgJNSvN8hTOuaHWqO1aqc0yBe4E54Xc
r+u1af6r6W6pVCMZGPB1pI/9+csbirt45Qi5vCTk5UrbtpcjWMQqCRag1YQj6QM9
A7o8daqG2ld9zB7JIaKC3c/qnITRJI9fCbPwPMieGcSB5US//kzeFb2KZTQVH0k9
RCobjPmDTTJj1PoVln3/jJ5/Qqr0mT1tX8ZPJpOQV5HJIR1zyPj/SrFTrzPxLWQP
N+UtM8Sio1fB/0XMUMNRTsfkTEBvAVg6SRFV9falUz4E/ogzFNpiHMTnF3IRO9fc
Tw9ZzoLMyo1mGPjBZCm8Xofstg8Fmb5e6Ri7goGAX61lpgP+ekCeATlPsyxutXUM
KKoe0PjP1i98znyktFyyj64+RK5RMXGKQgdtQ+Xc504xCt7LBceduMMBK/kVrHHa
GeGXAH3u/jov89r6Yo5EUEsToF7WqSR4FA1b+IC1YefxhlIuqNeUW8aOGxAYUTeP
VzVmQ0bBkBguMKKKCJe74WDfx3C6EpiHUdaw00W/Shj/AK/Psz2PiIp9Cozfpbwy
mgAWbfDIGmaVJQnyDgJ7aXP2X8n7izaGdWa4jjy7QULm5XxvT5aS1T9fgLMDJ0a4
tUoxWbZHyrPWVGY2ubHbMV1xuckzEzPFDgz9mVF4OBNW5nwLpNG13P4/rEDLoSsV
/3QZKwcK49IYWsbxdOXqnUGRslObs+fgHg7N3kJNCBz7gqeIQmYtM95+X0iG1tzT
MYsiz2zQPd5Oxols680KKoQXATM/w6D1PP2NnMaBo38PT0ZLPpcFidYVJ9WNSFfI
8pEtTMPF/6AVNTcFzAcbv1LX98QemHSsfHwczjs4WEkLpkw2+IyCzzFhssMk4PnG
sZCptMXfTIEgveQP1cJPKwWIhso1o7Gsg50/1+5EPIzYd84FM/Ipw1JHuKElo5rf
8OaVBfKwBq93eYI4MKjnft3cC46N7XDZ9pOVYWE1mFSWfzkHfb8kP9E8qVOZ9EKz
jXIVZr3UajnjrDdSgRK//mNNS7uvjA0xaIKUTcVqHZGhz00J61I7LOjSISMtYL5u
Eaad7FoI6knT9Jxf+2nPvKKyyTN48779ZIxqia56FzIVLExiInCyU3KaA3tdscQr
GMEE60ZBBuRPUkPRV8Vh57iNBLnEkjEyb7tnqCDoKKJ7rk4MrMUZOgVxJPC8D1G1
4nR+KpzucY70IOPOO0Fy8OjqaePeo9HBqS1RTWM4Yv9lOtctzqdW0t+XaP+CYb/T
TESLRlXcTusqfMzP4MUrcfHCCZ4foq3XV/QJNny/P/nxx9E3BSmSt14tdO/MJvLm
2m4Sfdpao4HtHXBSOcvnvb5Qy3hGVtb40b13ZE/AP2Uf3RyzniWeAxKumGjb/GOO
oq2F1VBvYANnAgejSyYAdafhwrrNlCJobscJonCNzh/T5VF0l5AYMfoCRY37bknn
05wtZV+1h2LlpsHB6LofurzMr5PKqE18EG1OxcF2wpOOgFMzP75a/Q8hSW4uKES4
mdBTodgu8hRPtnvMwlcJ5WYWOMeVqt2Hp+pPC7BQmRSlaNgTo1pDqvWWd6Btbnji
0kbIDTrj6O7V8464CV7be711s+EVdOwJTJ19BaQdR9R38E9K8cTQrfiZg5IkoSAY
3gqztZDAiPne38JMiFF4m1ItLTKraR6b2eOr/md2rkevFA7YM3u99lkdgM4ry0MN
TDuGczIE8tFeevCZzfERxWmmHrq0VSMdKESnkDX+geWw23ShTETaIMLX8HrSvGEY
eoAypK07myVLspnBwuqmB0iO3dBmLlnpSMsjxyhAnWNQD1stVQMB2BVKwyVlwbEH
HfDewnTcd8PDfrV4ZsraWXbssmPqhkrsjEnldDEIS+p8OX2sNPT/Pzrxr8mYe12u
6NNIkyJMpPhzw5Hi3zhpB1nyKwjSb2LgMxGtF67Zo26sqeVqH3jJ0pgu1cc4f81S
PPbFVWFBUYsbHUDhOWiy5Y/+yIMhIDNU8BADaWTVPVQ0vgRqPLxQar184ZJKtgjR
3MzYslnX5sFcPs05DM+4fVEgcFEsqA2Ymu/zCbN09FUo5Yz6QPNJpMKcG5/TYdv4
738o3uCkE4Fx8zF25/Bcgrqqxf5nUmdxXrWK6OZDc9qghCaXp7u6C+KnMMLYKTFW
VvxZs3FTQ6mzzJmykowwPa3950i7FsARuycuGIns4DC9JL6403+RCDrOAgoegskD
h/k4fjMajFW5cQo/13gpNLfzQsX6Zu1zmM6AF070zPHo7uoebYbYfkjGSc2/DtOL
/izzLhmYAMB9cbp+CCVmAUrPdZB5m9JOTieDsj0pU+8KBMslIuieoCNz7/10Y+Dy
Yy5c9QOeKNANz9ZzmYlSCr99WdfGMNfJGJ/263oqYpsuAIrBv5iznVK4umVG+Yfb
ls8RuRagiecoRELbQ9gM+rabA36lc91rWgbagsXv4tLSLsDqoFCCnZWr6yvTaKkM
/x5d78RQZWLDvciHNd7m7vt6OT1ExXcQ4F9u08iFkUAs5w5jYjHrfohr5jgrMpWm
UDx5Gf2GQerZwuT6S4xDa/n64RvuqiD8pwAvA/HWKR28tY03nuZnSZKQnd4ReL2r
2n4qBvCO4j+4xbvjngv1IqoewLBeODmFQMHb0G1HTCjuV+RBghoD10qrY5yzd1st
QNkaa3/9PRIK3QGchlmXsP4RPCtx4mxxyvAZMcvnk3VLi1vaNc0Mr8bi/3IXguRZ
e/8P5ccJma3jtqOhl2R1t9oAZXZwBZpNrkG3GkyAtfitkfI8TZLX7SiiDnziiujU
QRySOAX5ixe3HsVdy6RUaOGBBFM5MG63NeV63El54GCQT5Yp6gt85Xqdr7YXFS9q
dIcthUueHcYH02VchJY9kEVfZLrXx4McaxOb5F/gqYPGA35iNnGzTaOM1MM1fbcc
elVi+eUSP9Pe/ZRCxmVSR02HaAgKnQhfsUrDOJIR7YFFHnMunMsFI5szt+NZv/ms
MNgiDHKiLeygivDrcFE5EdaUK0yqJm+ODAdgEVZMEADoYbILIPKA1gSQC9ZwXZtk
R750Knh9WJ9zdi/MYT3emsNBAS6V+HGa3yAO4sYzfMZqW3anKXhDqf0K65titI5Y
72CT9xjZV6pfHfgBF7yh6tARxlLIi+Z3v1DFQGymPcPiDRYN6oUiGGrD7RftrZw9
96Wl2gMfh+l4XYxdXe7Vqn39CFfSYxzGCzVPXJN7JuuwZeUdIV5WflBtEVim7UTf
kQ+6fY5WTVneqm6f+y7nnLE+y0adttssTc0xjSDQXmtBpXk8d6d0prn3O0KuzLVr
/CuqmBZCJ5Nvzt6CgYGs8YuH96aEUMqWkNc26CwICPKUeSXlSdl3dmSMR6djnZkH
nDWqzod8NE5nkadtsYFQRczXrOS33NjlFyi2SyFWgE5hPGxylGX8pXcvkVJmc3nK
/Pj18LJCg0UkkMJCSjb47suoc1zGc4c3AM4jeuYPRjw1PkQvELLviT12MsXpEbKL
bz1OoaR9oRuldxsyYsEUnfH4v73ISlltaemSZOpV8sK2XwnmTJOd3nXCQd55uIRv
tFoF3EMftMRx56y7Kb853U4AKHjnucmrtcgHmRItoOfdaigFhZuhmcoySznONZZR
0fbAFHsPcjjvngGCKvyewXF3VZJchv71g9GvO2ClAM/yWL1aul1nmNCT+g942GMx
gzVJWKk4Y7I7k2qL100zByvD/tlVj58RiUXdjqsq1tWDHeoPngnYw1SqUsJvJlec
L2eS/xw2FQcI4acY+u1J5Bh+B06ZnBO4/17b9elW7xQzChQvYsgnSm05da2ykScO
zAZ3aGw5FBzSDfK2sQnGkbdMpgl3Xh0eDt54au3w2+nGmkF2zumkaYmqaL9Ebr1N
CSi4dOkilx3zxFnI0TKmT5J5Yw1S9lXJCYQV/yyFVT/0YzM/9NQTHvzMPjt5Cf/C
bFI2FShf8hhMVTUREp7Af1EM/Zs63KpKJadD6DmwtGj5ErS7xTQaLarTLySDbPkA
1KSKHEE+5fCfLrYD2fXLhwgqY5TWAc0g/ewAdY7tZQw81CwiLYf4uTDwVOM+4O/t
5fIi6H4XiOOK/M3B9oxgnn4vOtNq0udPxYjXrKLGsn7L4kGeaG+jaXqsyQpx3qsc
eimr/pKdL4xe1UOpWkuskJvVHdlhG73TfpzuvyGNifCxLSDBvPpKHlTsAatMuprD
sh5jP2iUnXTkpOg/+jo30por8XagzPuKajYvNAmksTZWa7649Fbc/J/i0vPSYLS9
/WBGphcrwGT/xYnOXc7QvnrQMafMN2GKOv+gak36vb5IZv0m91IMSUUJL/TVm5Zn
KdCUJn8CmXjBELa2YiPeX8bqx2MXeHnWNS1/c2wuCLCqI/QOBrqza0FIY14uNTNz
XQQEqKbgPE7gXM48xoUX2/O5VhgucwsA0uz9LJ1AnVonYi31PO1mtmTaX7JsUNYj
Mq23Ap62wfxmaRq3FZQWh36yOnt2qOzOzYlSgtcWetDILcHX8H+jYWk9EWtFOw0k
otwMW3m3hqBXkccSqpENTppYIf0LSfiufv6iK8oy/gVe+D1iYqaSF0XYRFCdQZT9
3OZ27+2QX0DYdeuDmZ0Sf4B2vAX2iK8GAJaoV/Me812oSl4NjQjksPR9xWzeNfkK
ibk40+Hfb6D+cII3JAQiH57hntyhcguTfFvbarEaEpoOH0l1mvCMcJi8eAhtNcc8
vXXgD1HlNaGe5+B7/AMi0JeE6yvhVqQNZvuUK74DUgaBRpTPIZsb0gEvPROZJwxU
+rUxlU/bsXHtbLZHZFDrxoAaBHrgk0vlB3CNZJyDz9GBIfKEfRPzGNG/efYEfbyf
UT3P7jrCa0otvtouvbsxk6/u5qVjSYVx5elq4kN9VmC1agikfFb1L9nnsVU3cDYi
JxDXkf2iQmUSHO3uPMJ0AU39Gd56ipPXraqZOqpoCCmFNe11ZoOkDZ587mfnIlP1
Z0Y3IyTU/yo1W6KG0i9Mf5piBWwHBg7ZOZaPwE1/wllH2xzQ48Y2RfBjM3ehrhJV
+nIlt9b0gM5y3S+ELDJRF5+RHVGWZ8nTIa5yoJt70iIq8VH4m2pNk/3GusIx/6Ho
uWDRn90loHzYCLYR5Rd10ZhPygcbXndiKXY4OYUYhrnumpfegcCsDHCWqiN9TU2t
fw8sUBT59oIGB00jfJm0d0EoXppI8wuJGyXufj3OYyON6AeREDt2NXKdjCKIo8iE
aPu3Pj5Mgyr8JaXvH14FvhXl+P7AXMJiIZtI7EbDixaVti49aKZJ5uE2Xn66s8vj
Wg1UL2x6JjdDF6M02qOys+Mzsdh0/mt6b1EExsMFGek6FwXCuPZpQMIePYalGaPM
T4/w6YqylT4Gx7gn5QtdWKySX6Et+jErUyvJ4nhIooh25BOZiRa89b2Iwgxo8wwH
JRvWDhPFqf+xoPuepJWqDeE5hQhxKVy2NinHuEEObUisfEw2AtINKsNqv/kGqQQw
hli0LuGwUVk2h1lAcvelsuBFMYteL0ZAsgrVT+FLCTimW0R8t1u3b0VTqO2hZ4KM
eZ6hHjV5gQVtzFVeOdklm87Xu2G4bOImnfEd/ubgoDu8LFmK0MksCTZis9bBVqUX
scEcBmJ2VSbN73oCAPYc0RwktjxF2nZbwr9FGDZ7/+uX+MdKeYGGuYtXxoISufx2
KeZ09XAPcdKDTasNxrY3/Wa4mWyAJ3CHoHWijHYOFsY7h0PNpAe8Cl4/xk22n1ac
zBb29/UiglCICbXKMa/HucQCxyN5jygGBx136RcJd+ZTS3ivunMOjPTRz7JbPPnj
f3dZ/JlkY4PUAdp/vps6ZedXAqC1ECfeBpvXHQ/VOTJfWoKl9yRRMoj2jU4QvmLP
Eo0W2bED6PbTrOmlkMM5nroE+OGFOTCnpvtyk6ojJ2As78DzhN8wlOGMp3Wth4TS
XkdlBaaCUNmqD9PVoGtY5hNybNT6LQ5zgayqtrdliwpVmCDBoywNQukvAdPdn4HE
r22S+bw7cAYFNjwWPQEaNyihYV29vLgSBuOKvAwKXp2Z6hYUwMUHoel1bBqmNa8k
41DdO6nlDsxMyWB+QkdtVlvF6yi6/7SJuBw6GkNQNEUVd6WoVNfu7ax7tcDukmiG
NX80n+TGSimpCq7GSZlrUwYb41QsntMzZYD+H2mzvApDZrKyKdpsvIuWiwoJn5eP
smqL1omUI9lmRYsnNl3FGavBWg0WuMFNOfBPTq5LQiDwih+OfU1/PAQuATbmcNcF
JyBzJa3MiNrgUInWZehZrb+8+hV2/tDZ7mJaoPi9D+qyK6WDK9Sc+Xq8k218XXO3
7gPQkzyRjDdaj8O0IZnCVLwPjYNwXFYTL5xY546ygfU5i3YzHTF0sXAqQi3evYiy
frjIulwJsciFqxeKbZAH799jA13WROaQTccomyjXzkSeiVLx5G0x/tivaIOGCWp8
R7XO9wMDanI51icr8arP2KEcxvUiqtMaEfOSCbg8TijtVqKyb4ZKdiT8LDG9wsVP
KmX396C4ha/tkeqNWlhqoadKdH9s2pQ1ARczX50t1uy139DLHTaPK8jCFEcTPIsn
XdfWtlWiUtvYhQwBAGkJT67yeCDL1WOdlDDUrk1l1UxySfdG0amYNq5BirYTb5VA
GISchlu/cljNiCzVu0yaNNPJtiZqLMU0rR7fUrebHNsTyXfDfNuLH8VAjMtuR+L1
mLVYz7kQJ7I4X6zHhgGaeQoDqQJ8ig96EAzLfvZrr6jytQEU4IEJhvaYNorG+07S
EWFzKFWJlZqV9Htd+GHCDrrKCGCEXgbaryD+4fpRTVg7XMjeRt7fjJsDfTdQVSQl
wAxhv20BXZKDNT4D+dyecthJ9dKCx0/zq31mdHGmCg2Qh8qAbJzlujWBuN64wZgH
laYJXtXsuh1OkR4dU3W44Xxq/U4T0K4vJ19ffds60s9jQbgl8F/QgtZ0McVPIkNw
FhE3Cohwv44c4NTb7thgFo0sl7QU0NwHyvAMCOUC3mYlSxxbzmjIm0rywDkyG2QN
ZKrn0Vnyl14cBG3HMZpEQrEa+rZG5We4drXA87tttNysQ804fNpikKtpV+d+W2aS
mYy+g4lfSZAHDdlcJa2iyKMqmJatypNlGNXaLIwKiQ0kX98/vqqnTzrw4L65rX2R
kdxDQFP+xkjh+SIdGwIkkHbdJYbzprs/SOztiBTBWnzXHBB3qxHDdkqfV4QL2mvI
TQqwebqWbbPkD+teB2XZtZm0Ictc/yNoAn/pdyLBQOw6SxfZTTnb88B+6kpFyV9q
mWygQm+EZZTba/WtU73abjmbQhsxQTVX/56XSFcZYSqir1eEv+eFDnWPU8O2Y7qB
vjcK+YjZZouijumq2qvnFTy4NVH/hMpAp6dbaTOlPkHBUdbwspxXeqDIrgHqLgQy
ZmTM08r6srw62KpFGNhOyOGj5AsQOmV3K/mdKotMUyViLjiyE0QUknLDSGv0hiHB
sr9VMo26d3ObEILkmBxOJ9Ll9/C/3VyA21KjzeOB66mD+hPRx26WNsX7NRoICNSb
NAaTIX2sdOFIyr9hA1XAGY1hbY1+9/+9EPcLlpGu3NPJ0XGq2/keggOwcYxEqw/y
HeuUslKcP7UqQQTNslqg2oS5j3x+zPSI0fy5SYWqh7hQ7oPyUgDjgAS0bR4pAEA5
yTeM4py74OWq2A5Tfk6Jkq3OeTzOrVzWQdTlbSgboNHdZ0OVcWQkz2WylGxWdfh5
22wUaPE5CvY9khyQyZfj//MWbHCN+OuvPA8+IR4PbMAfQsWftetGENTcaeX7sef+
NgZTZ6+1EWQJvjyfOEi5IdLKPDQ2hQPNoEgW2gSLKRRdFJtKOAwOq3AtGVTtSwzP
4HPB1gVR4Lo4Z0ejaHtbBtm8LY0NoRzdCCX7FGAuZzwvzCKBh25Kf4MTPW+WT8Cr
bl/JbRFZQDJ1On4OxoRr79gaRqLwVqPmPiWtP2M199PueM0Quy+THXmvFV/McUyi
krYCh7Ftn6rycBh7FqwK9OBlx1CBhbfU25RAmxc/oSOzCkipxUl/LZkE1f18iYt7
eMSGHC24N70sltfau505hCKvQQYDQftlV+VIBwIbNnKisE80I2zqARjRGNcxUG3e
mlaI/D/4TnhzP7uo9DhRPjHVwxgLGmn/VsARpXzXAqraFlH/VqsKdplIpKOx1jgU
1l/o2+FGue76aMdtBg35wwqY5rPya049dY4k8HUFFUwbpYqCYz84VtbXYD/kw8we
FoEVSQ8WvJDiUTrmB1/EdRwnf06eP0Ky9f8k/nbzY5qCx9fYsgngSV3kpUXSqZ8s
N7FAiJ/sjOeIRFNwWHMKWkmazYRmvIzn6KMIQG2Z6ebMrTXL3nsIh3BD8PvTfcPr
PoQt0rWQFgnlVm4xyrie35cdplEHffrWypBzuiqyFpIyxSeEuLm87naGW3eXTcIu
nNnsPGcG4fHkFQJp2ZeMB3BxePB/hs5OWGFhxnxdKC+cEfKum3XXsIlVCQ1GZvy1
qwI24aIr8FjDKO6iUZrTNf47t9yd6+bhkzfQ2EteAyODn4XzitDc/fcmmjecral1
+cuRXHNfvqrrGgNn7G4s8lc/zo2KT2NMXxR9+unGdFmlk68nRs7Z7mBU6pHmC1Jw
YxKgKjCTESYBiBREdoT4lI/oo8AOj0Tcp4v6Y/JNoAR+RMd6lQBxhZdueiCyFeIb
lOBCU8gKd4MKusVBtjDfZAwbVtOYMUwBwDwIdULH59a4fsIPGa+7LNBfxlbhZkhJ
FnnggZlN8hufTtZSwglION7NLpi5vdDzCHmxbFv/M80Ejc5uL7Z3pvIEFSXjD6Wu
ZM3t9u5CMd/9yLyf2EUiIOgst4GenAvwSL8vR1ZppVwdv54Vmcah0X72eDMEmYAM
4TIGeVFExgSXfG4dCxCz7mtEUZDS6UoDQfxv9A72BGpQuZhqVnHTWW7tMRzjV0yH
Owmt4R2qqD3BBm5pMZAVv8vO2LJ52WaWtBgBpowEhgpoagTi7zf+4yW951Li8B68
PaCARstt4BvnT+tM5ORYupPZSpoZ7D02rhZ4E3VGxTLS4c5UElFBoCJVIBq09g2R
cJj/sUWxNGOVG09XJuZXT0w0UwRmmBM/aUw6O2dHSOyTQH4LfiIKoxId2WKHe8UT
CinTrgmfag5XLNkaXY3MjixV0BEiOt67ZabPG2alHrM0o2tMZq4vAaTKariA/w0u
0HEp14a11osWMzi1/EyIQb6BixuvLvOfGqepC9sHovvAoFdVBj34zAKIBl6Jp6oE
PLGY2cQv8Ey0T5kW/npaXVzUQej8G1gB/5CqnTwo3Alnsxp61nm+thysjzzDoIOl
MRHQYsxoskxYa6i4HpKg1QNMnjImVUaJwBkIUIGZugh0MyFdh9xE+nwZtZ0JE92S
bKz8Jl2ezJLYgADlCO7S3P0vN1JVrUFGg9n1jlRUg+j7ghusd953n8w3NK4ae7tm
+PW6HKmL5DYzr+VChZ3gmOAWc3dNb1Gjnp3Sl3eGnNL69OpGAUoFq3S2uu9iEZZe
Io4K3Q3hm90Twmqh6C4AO2tTlc9C0WOVDIkXaZ65RUfxvPpoN0rI8RRwiYpkYU/i
DVRZCYbY+eGFFrQSTXZ1+3x56DXvwzaue/vmwydQTys2mEy4RpioaTTjlBQHfnIu
A4jX8m01X/woWlVjCYvpnKDYIrnU9+/ym/GGTh3B4Q0U1ImGeXMGMvw2ycblya5x
kz7fwY19YicRrpnSWOJ9beJetYUAYGm+e278dGnjnNLL5M4nKk/sN9gbwRfxOYvu
mFaidRR8X6+iWBsXDrP7fF05yJYal9QhNjs3TMKXhB+vuk4jEDbVemZEVncsTdHK
ntxWKwOy0Ak72uU7jh69VJzceejHv4oUnbwRmwT4kCstJn7p6XMYAwrwQL4nPdoy
Tka+hKl5AN4su/Z+z2iGmJMi93udJrzYVzw2itaTbdnqxO7YHypYc/LoFessX1tg
Dge/qY/UiK5EPfdAy+4mVN5wE2Cklt00vAIQU5hEzwjBblDOCf5N0Ui++r24E7D8
g4k76bWWrcOX/EnGbdnatBv0NgdgsrNaB/5Gs4YkyRYUVjpp7Qz7txJ/M1kP/Xwa
7UKmw8rGkpacl4GmTpKxkvlnSU2pjDNxQ/nlauQOc7hGo5AAXLzdPDWyx8+6IvRT
TKgrFiXa61JPe90PYH7wQnNPFliv4rp1JKdlvssO7m+eqbCClt5skLA4Bffr8lV0
quTdXmVPGgh2IOPmqgwe1feqgpT0es1i1ndIIOuUViPWG6o1IfQjZJQekKyhd1ye
FZFLhDZ1ryICgx3uFnVLS0zrI2JIZjtooG897UP7ZuO/bwBZ4XCPHOsR2hO6LxxI
y5cZf1S8Gr2rPmErBe/yAqUVgXGAbKUdsPgXHVQDcMFDWb8NoAhXkLJU2z9s1X2D
wGsbNi7nVAc7/NuAOrZknEtbQjVJeY1dN12qm3z0l70cL5QUvrQI2eeRxt9s/k6Y
o6AJNl0JKHl+Br/Mn0fLjqrg9VwJsJypSnlo0ilAh259Tc/xuTwMoTy00588lHlk
T3/w2LHeaP+S4WCaiySQkTl2llGHu8ueUht6NKh79EthY63E+F37PLBB9gYv6+G/
N7pHeLlkFLBlzchs0zR7YnE1U9ChQips7keu6OB29Bfe+hd62NmojEqqec5MF5gL
7F8FMaysloKBCuF9qy4rCRtiJZgrSTyg6JD5pLc2zSC73q/1t3eUoESE7QO8Aqqf
k7nv162Ahv4NqCfrC5hWD1d/WhL2XSIrAA4izIo2LxxYPGK3vyNSzdf47kWPB9Xa
4zx+HtxMyZW41HFj0lDrjDfm9XHZ5e+CmKdr8UJc8KHNCiW+HZxdiJzUWz8blJ0X
RiTcYRO/ePaJpa7ji+jeP72ingKiZEU3BbBdfwcw6WABxII1830aqT+dcZyksDA3
mWZ5YGK3noqSbqBfXfXGPVZEkhZx5BlpQqI+uCY+BThd/faYvJuFI9inV5qmMpgM
ebGMeJMZiZXJb/7Da91pWOgmC6HxVoHqn3ATXGOwArSogAEKi7lELEorZRFHahSX
gxjIcITbYUdus9pn9+eeRG8k1Nz2NmAL2kHJoYMeAeOzvyq2qFajLMbRY5dERYV4
Kxc/i6sk6bJ6fAiRLfLd1KAFHwUXBv/Yc+fH8U2HLl7H6CKIUABxPWROzGApQZqZ
yrTnR+Tef29JkWfl14hxL4tn9/c33iNEkk8eeDxP5oeqSILBHNoWr3w0ndGH9f69
8NqleYIoDWrueNprBJy0XQMy4N7z9UXgMmfhabunnO65RhMYtU4Wc6cq80rDGhFr
l37hQ5mkeNDS6JrND0rZ1W5xbKBFZxcRgr11m0d6nEhit09RqGe2QQvkCBjHuX7k
4UITs/Xh1CEWhuiVoj4+AdxM026MxwyxKrvWjQa9O/EYbgOUyCojlwWAvag8dCPQ
qx+pYdHP4UZdxoTSrrSyYRou3JwmRTPjIS/v0CVSxbYrsGUc9neBeznwP5NFMRlR
HvBxs0QZdTweJfiFtQl+tO3UucRJ8X5LiQ6NXKwfp/BBxbmT0YRH2tq2yoTEKyLU
+6uEDGsSq9WSIiji4K63e3N5/JSdxL/Nd3h3Jbtn5sESQSKInkuqtHOn/LBPUHLf
hcbxyy3QFfH0lihXbC7iYv/RsK5U0mLzA2cEIA//2Kt48zlZTctisATUSFjRnEDi
hdJ6ADC4Jj+lEizhfyufYbvh/Pl9Mo6H0dECh1SPdduvUs87Z4JAENhLiixip+4k
7+dmr7SXxSUQvchIGCdC+YqNUPanbMTRJJxRLRJzJ00Xn2FP8kK26Quk0d00tVUQ
JJalTHMF2JiYYd5ofK/5rCQfzkfgRNmN4IMeahjTiZY0V+PG91lmJEYiLrJvwBo5
r/d52PcZ4GHKztNQ5/CC58zWUJtPSlPh47FT5Ik7R4c3XGpoROleSGhJWmYpw3GW
hcWsihsnEzlzFfU62S6NA/FK4BYIcGJunIpap9yhG3fx9vqGg9JI29lleXMEGDVg
cS3bDXIiLsmaYUqLXRe8edZk8470wVmVG3MMVvUnZbA+Kgz/AZzfmKxrPu8RecNH
Fc5t3QZTpmu1iEC2bA4uzLbV2wAUb9Kxk6OZ3L3Ai57rHj5uvJsmsl9kYiJtsxWd
okm2ChVWuD0eie7bikXylEEJEijJdI21XD0m20NnJHuEtf/Wu931uiWANyNDD828
tbTfvwak/XTp9qoGdRcnChuBIR4q+r1zf/KGLZlK0p5fDXwH8Qm3+bj0TYzAp/8v
KMxZ+EkUacRo1FGZbKC5TmjahXrtbddsbiA1qEPJ7loGPQ/QNcXGcYP4EssJNNUn
N5v43ovUoPCnnPuWNESpZv44iC+AwmE54Jp46p3Q5pazJqqEBWzyjfVQjOtaZZxg
1YzJtkIyiR4HdwM+qIxhqZ4Tq06gClIoFUhtk7tpuYQSXyCSQPTzp/XJdeMRisKr
ZCQJlDCWzap5ZURDht535xVE60sFmNUlVAjEGkusb4TY2DgB7S+R3Iv4zUa8eQFA
mqvhLe4P3pRNaX7TNvF/i8qMsn6cki41+x5h+xLCni1qOIdUI/hYj2ljjK806AS3
QtE7D56n0CKAauXpE1ISPlT8NfIdr70xTUZahqbjfnr4HlouWFTwmpH4ByZUXHD0
0bPutgGSUxZgxRjllglpdpC0StuQnz+H6wRSkAqzyDo9NQo8f8w6YeTs1nVrE/vC
mGOHsDCbwkEwgmkLGgAzyThGmAwjX+T4tLyqMRGF0BBvZB6EXnsLgm4PI/Fswekk
to/kcYwlR3GbL6Iu5uNdJt/1DIEqcaR75eHz+Jj3FILqlgQxUoqqI4VheVs9xq4k
UBewYlBv37HMmhrssIGZk74n4UYM9xZ63rH+bf8rWq3S24LmafWrMGoMQ7/Pc6jc
Kcd97bVYptr1CKATckdkO1AnC97gAI5VDBvX1hNJxnBz3Q3GHF7YKk5hkz5yrQ6Y
xoJ5PEvi8sT7fexo+4wDBeTbbarMXw+GFQr2k44iC4sDinZ+CxjSqhT4EkX669mQ
hVEghmuqfX1/8MkXWWS+mnvlJekDCg49aCYae6465N04M+Kmp1E9hjt8jjiwTBi1
CJvDOiDfuqHRLCMx/RhChHeEu1eECh2syM/enH5RAKxgGmwhztpU8YDDzsl6sHZ8
rIyQqx3QSuDA1njf9Sz7H9B7VIZiXEZI4MZUwqn1M+ENH4GuUKqENOQ1uDGRvR6n
lOvU+9rRW6GBN//AjeKefoLPkYtClfthTSzHlyHy6kHgBSrFulI3fB1L2rXU+Pwv
gNC+UBiF1qkGDqJqIT2OI74DWqRRIQzld1l5eZ8Uz7sXXwPtL4teFsMs7xeGJ9TA
VyZMkmZeOUMTCnrkQ0G9VSc6CUf/AXwp4bODi6aD5A05dMRT5UeJ0h4b3TaPcTk0
cxf9bjtZZC9nGc2UYfk0Kw7FXLir6ymtu4z3a1zPq2k/2zFq4qUdv0RPbUPc7Ouk
lMf+htTZqRe89j7grFp/3r0r6W2ZdmjN2EdWSPYlUTxR128k5YdZCiIIxKKzKUfI
A7mtnYJsDvK2MvLQVrDrnYafy4sfUYx/lwudHkmKcaaSqiMViVPwMQudx9omiXBt
aXFOSmLtHmCFtRD0FzAZlSh3WHu2VxS37SPo5+PlaA+VQ2Ws7k9Pe09ZmQskYRlB
GhjdPWTuqcF6hsIYutSwuyMqI9b3TD3KvpT8G7yGqo62uQGXMxQ9ix2CxdoewdYH
U8fpAb7ImQamuYgoKnw0UyfcgyveCCGbpQOjvWXglL9wFUTO2FQ7PaxKsbUWUOSg
+mWfU47SorzEEZO0p1MHuXmxH1JcfwKoutB13FoLeRWqHXGJaOYQbh4l+il22A5D
ziAZ8CfGnDYpt5erWfAiG0u80jrFHOePnR9QKWyWDcP4z9OksdCC3xrTdomLRWF2
IIEPHG6AZcVnyllEFUCfUB9PPtkR9PXWBpHqx9cAO+5q5Ho+UAJGrt/QLjYK5mEG
DUBWx3Shs/y2dCUWQypjwNIE3n1eiWdx5EEFnSBIv0FKt5pp9J0bpqYSnjpff9fK
Q9+kd3ZdfBGeHdZDyszsbaB4DWKCPga4JqaaxHiya0dsd3EDHd/kH3qRia5D6vDA
exexNJ6RgUl8sInotQW07sgCY816a7iGwZe42JWcEDxoHb3/ibBtAau6SpZHQggi
em0vH7DnEVBOb12wtj2bLssvp6Xd/JYBK1fBJR+WfAr+apPVjz4el2Dz1Xhxrv6o
7wszxw+WqCt8BpWgRw3M8IjmfVSCsXYM1kGeyFZRi57bFH0UwI+JINcJ4+uh014c
LKSW73IN3nxGwl8NrJM3B1w3d/a7jBWTZMkwAS6txgxn295krag4JxdAGbQyGy5T
UIt8OtmdiL5xitmbEKfR+k1GXeY26vdXdqX+0GoirjeK/Qi8gnoWCjCA4j6Fbx73
kXDNLhfJJCIj3FaXb2sxxibnrjORZDHPLujrx7GRiLjWo3B7sYXoMoiydeSyTQJW
4sNkdpRGCN9E4uWM3inkIzTgWUJ/xcKkYFBP2AawaGzzNCDQ9qFDRY+1kW/BzwSj
+acUkXR8YS2T+7ii7EgVfxtFhAKNxRMwA0RTGGb4fyKAf1+ieH7UNs4J4F0gC/+X
lclCknXkAE2RI6QVx6M3p6i7tPVIdEInTfV4+LWnRocYrl9758RC/JZa3JQoJPgS
XP81inC7UvM4N0tZvgo6up5EAfJ3e3oZ5XujwUzIB66GXXqPt7ix7yQKtoyZQ8XE
yWavcplOAi2PEEeMwN7NGW+/jzmyRde4FD8DNx9HLV6Gajxjfc65RcA2P5K4h4Im
L4XFnwjnAkBJMhaMv+FDVQOG95FNL/+3EnqzkDd2NzMyp5pyHyPAaV7O2sOFbWio
+xRayyYAEdQsJhTI8YXZXu5BD15YBX745+rc8h1fg0ctxAU55eXmC9owxlUrLxlY
d7OtYmprKQaaV+45Nyy0tdN49cZeIx7dgPLwCN+nd1tg4WqCJ3esT/jODqNfb+od
VyAn+3vSAkhrukO2/waMKWGr0FUVVOXTkHhBl6FbPZ1J9N1qJugtux03Hd5qsvb+
479ICjhY/TGXLkROIIXHWTpIMXdUwW/P3ZDpTp5G31qbY5n98/jtFHygjAFdedgY
dcP7HMZnUWh524QXKMtQkLvQVXrHyo4UlOXxV32/NHdyeCODQ0vAtSwaJ6uDGi8w
A0tgy5HxkczTpnz3bfxPBsrQkkF6o8x0CWRlZqXEjnzp8+NnTUB4NM1QRDam06b0
V0mFepB6GdY17HCvyjMTEXbPZmrlHgASXsvHH1iWh3dSwP/ZL/TCp1svyVsfSLPo
DguTnyUyezRzVPVJDxNZPkG5Y6BO8xOfs5C9ep78pw0DxX3HYV89Yi9fh6z2Y6xP
kMBihGnZg9e0jI8PbHYzlz2qOgXgqh9yEUgXe+G9rTIkHH/1O11IOf7sRpYVMTYD
qQixRwaNu9baqVRf26OJT7iSYQLElPdNJ1JS0uGzWP6BD+l02zJYeNi+ywdO3tc+
bmWx/YOUeTNcrdS/xUXtt5HnsjIokN8PNpg7iGijfZBEjvx4EEoROwPq+KyHOS96
yP5pXu31MPZi4iKsUjZZ1nKakQnCSrUBYWjTK1Gi6qB/HvwIDbtctbXGIgdeTQkU
ph2Rulv78xm2/mowDX/UeltXt4Ns2aT3b1yhgCgVZ39Qdd2dXX5PCm7qUphytOIm
RFf7pvkETWHDEhRCz8bvQ1pUcGKA6zviRKOG/c+Sxr0xMapDGp86/BxGTreJHf2L
p6/X1Z/NAbZAug+LG1Py40FLtFWCCSuR1m2US/0oI/zaOotdRvUJjn7l2iYO4KJV
qnOHAiTo2QZlMgdLCjKTs6hmq16M30D3cAazgw4e7K0k3WrbSSVI556dXlIbIQNT
snLPD94TJrNTHjEtMwRg5H+Qn6cL5snnKQo9dVcnxR/eAdDW99ZL+NahiMTzVasn
8g4RFqPrQQVEeAHu1wERpADlp/9B7Es+Cg/lGtAURPARwsPlJfMOPlYTmV9vjQAb
0C61aB3mjKZIF14Z/XsKxdTgLDdkvLmw/TTU2V0K5ATHHIB+5GRfAW8As3/ibUhF
c3xyaNlYf9u1/ZvDQNLKbwMtdbCYp8HNwSkilNMFMMfAIeMAqMMtDAhqbBHtNSw8
NWPa/df5VlTW7bDsy8il/5gaQlvpnN9C7vb0VasrG0GUjumtJ9E/XzgXkBJbJNMe
wBK7M6gEtM+AJpHzD42IikPyzxBhGkrXGVOYpaECTWj3Euxs5xG3nbjbYZVrV6vz
O/WVMLXaFVpY0S1M3AuTpb9xJrEkhxRzCTvhmMtxsalCHXeNb7WLcxuouET5wFJe
p22sf8NpzTX1od5mFL9hya86hRSJArgqOMiw4Pmz8SOb8iP6e/EWP3WSzuVK90lP
vZUWxembHlyg0ydRigwVTjI1FpQ4KLyWnuMCb+i/1Un9SpX7RVeMdMf/Mi5ZRPzu
MC8tOKrKOnjuT87+5JXin0qCoQPf1Nlk8NIKkx6C/qf81bb5ozS/CYKh6U975u1g
zV5W9x5ML6IaOCOPq7UdqVDi1E8AWZmtkplleV0TF66/necb3zZrGnl5YX3Hl6gZ
LVRv20GdkqcHRcrRVZgPuzrDAX7oXX1m6oOsYepN0ttrpXEynst3T7fJDd4EKLNP
mNpn/J3qtEr9K1JKJwcAfNh8s2xYa+HFvO/WoICxxkMh4Aw9P9V2mFEsBQqu1BVC
jrwMYPUyVr0WSyLQXOda+AMkXYLIFn1w9h4AS58ZVOEXwN83s43ErX7X0vAmt8Qt
IO3MzBiPu/6Wi766VdZ4UIVwpS3u8ARdzKERhxK05sGq3MDHNHZrcxdebN2n8/nG
vXMsk6doOvLYtWUfyuIczHKc3SB69dVHSTHV6ja59UnD8ZhiaGUDyuKz81Ja0vOK
u7H6Ye4ykxlCUcktdI4fV8q0PbY+vTWFO1ptk/C2F9ZaqXUgn3snLV4gc6b87Vn8
fU636VtzWaPxfZHfPiwjJjLe1oqE/eaqCOMoBysMIS/L5LorKU61jauCHG46ChRZ
lG5V/mD2xSRgU9qfmJMaD+fO1RuaoxCLPOYqnBqBDacxCrXuNRVkTYctNkfUC5oE
7ZD4mWAS4sDwd1w/wo/RPPMVDmVJJHrgWaLBvxwGwxBBfcyyxtKioHvQ0mtfKELa
L9qXN30munz+XfJN4+1W5kOezNieBR6xLQVvK7WkhvozCsaQ/KJ9RqOe7GBwCWyQ
O+Rp1RoshSm8wMAak4HFyGg3Vc2CoUSStESk/5AXN22rAgFZ7tJi7pTxFK2ma/01
AklbQ38vKylqNJW/4HBYAzNAY4tT8uIuS6WGFYFaIAVTq5rqJz9XnzCZylzxB4P+
cAOxdncYVn0F0qo9zXpo8PGV15QwO2klVt5cCZuT6aZyFZMdcZ5D5IOG3sAQKOZp
4iDxaKIGkZ3Pg0hhKcB5MhCx8jnsDGHHkygv3b/NIlzI+o8jzAlKJJvcuhRn5BNF
XU0NsjP9vozjZ23Ldg4iwnVLg2kS2bRSGO7mFEvwnvdsMqUf3oWrLcDFsqJESp4m
AYRFWnSaSpvux153fSfsJbBHDEOlwErpb0vI9mY94O6P9r2GNVb61upO2klCI3Rh
ypmFkeC9HuLacEur0vlWxNDD1wrfFyiwT/Cu0R/MbnhLAZJQblzDcPWAIIkFY60r
OI7ghHHHtRvVZB/yszUg2DBr5DfsWJhEBBs2qyzPhZHWefOf9jEBYwA5qbZTsK2V
ovjcZYj0PLh/7uvjLpOtAQ8IiChKwNiWga8habWk/Mn/NlVgAsQiKNlzq39+1141
ve29aWqGnrN+VyXbwErpmRot9tqjrVcHl2s58lFaQoMPu/I2hFs7x1sQvWlSgjqb
dj/L5ZHTIfWvmW/ESWFuDmKf+T7tHGsShqHR7FZqyPQqgLsLm0OnZV97H5QDMEdf
/9/5vKj3GCFnEm24XFFH/XW6FVUEhDpebq+G5BYqZayClQYJT7oW4kN3tkaiVL22
v7O3ximDCZGh8xCLh3jitgsKCPyf37l2fFKspBss1WRW1KUqGppPMq/0O35P2NJp
Cddg4O3vOTYX2RFWpsyfQZyuM6onTDNjKNrkU58mHqXSRy1AFtIMcyIxw/kfVOOd
mQ3QgFoWCU3t2xzeSvVCJJ9j3NM/IxnpTjXoFCKM+5GSX0Ew0Pr0ZPpiMqH1UuEO
nCZowLVo+6aoSqqRA5qYWVBIUfYsq/2Dc9NWBQ2MkVKY1TC6W+q/5XhTvRNs6H1w
idGk+0Qlrw9fTKYjnO9qDnE+m/hDzBtKIqm7lLh+awc3yrxC8WEsvcOU4gMCUOLt
eW7LkrupFslGXTRn3aioozph6ItpE87qqR1PeKfw8mmwgwbIt9RRJJ9F5wMpik3d
C3rg95enWnznEUA9KoDP+7d3i7FDGeN/68C9SKReaiWk1VOFyIVHv5s1RzS8Dyom
tH9lVBHCLxpCJOXaGdNoH98qzm/iFXiYWLd6OxcSk5vUW45x4MfEEJT4k07LcpSk
/SZs4o5G6d2Z2AWTpybSjrAZulTcAbsDAU9ouWiByO4mICQ1dMsN/xbzoc5SPox2
Z1VZSsKm+QrYLgT7UCzQYFyRu0K7RYDtT9mfDiIDMt1/OoLPLcxcfcibH2yEGsus
4B+Q+C6TPi299QZMtMB9c/pJ17scdZIaOvH0TfXGpt5B4p+lt9w7t0sEQYHXhSsm
dqTHl1Sifz74qdlQGJBT6Ox4bA6kfHr0G/lPKiZcPllCWmc0IFCH+JK3/Riv9A+z
CfOhdVuglXmJwFb9FBM2brZ23Ax78AtPW24kcv4VGopL8DREHrntOMfEzxicVsLu
L08LCzymQ4dvSgvjYb1s0rm4ityWelUML2UOjzNDEbuUlWwOJOYoNVXVz6fkiUyk
e4LHV12dnTQxjKYlIwOWPMeJx7/clY4O6CIxqVuoPp0rDncnMA7AC+TWtXsx/TxE
TmmLQXXVeuI7oYN4T59KgElqqUnlrr3RjiLLIE+LwbZ1qsoJ0WPZ8R3ogbcVaWHV
ij21Gw6YwAT8jIARMOvozFugAXcDbcclkL128cjYOiMGW7hvqYwsaXizRHjVJzHs
eDGsaoi3UAiPRcIxqSqrWukFp7P0RDipDnpIMxJtltOYuPUmV/VT9yhoEkJm7Dhj
28kLn6EibXYeNWjHnv/6uIK2dKk2sXfJ3nIYFZdnLO5C8T/uEEwCrdFb9y9om5mm
WkfSjt6cHprmIgXUZdjIEAC2XW54S91Cj1A9hGUp9DqwVYaEki7snBrNbMMvijAg
GTop2VHmsuR3E2uHL+IrmB/eoJNozppBY4x9KapbOcKZYbMxs9LSPY912k1e6bFq
qSYs9/qAieJaKzd7MNUWsgKRLaB83QkBLGmoHM4TyYU7TEGeYTjEDD11TljaNtPF
MJ1uSWn8ugpLBOyBAUYZ0NnhA24u9r4A+mb4YoaXwHSkg/5+6/+8etEMnumSLXV6
NJXK+94nqW9jPZLEUQAEFDi09oA3VNPUA3KHuAUbPPnOPXiFvZ1++Jk4WoCvPFDX
PNABg1I3HIZ3smJErW9JXLS91RAOoqYhW+4kqWnc4DdBQg1wZ5U/ijtSxvvYwHhC
EEgM1cggoPndJSV9C8K9YleezNwLuSOvcZxEjrEHJbEc235Aa2cjjyAasttn+g9v
8s9KAe4bhxfL47MIYi7lMxgUtfEcEfYG8pbIM+eHHPYXKf0Mc+kNHuskANttrzds
4+7lyXsHtNhoOfRtlp0CK5IM9dyS6tvu+3tGPmjR3oB6IrqQ88VKN9EDEapk0gSE
Eja8ES8F3mXbD1npE/QaItfgAPhWkVbXp+ueUNS68m6i2z3x50DJ7b/Wi2ECWB5M
G85D69/KigU/M92SGNS1VhiUjuLTNgjI3BCF3XDNND6h6Dhsvb+IlVm6KisBligO
Gvp+eJUcGAQ5LGZZNwq2lpoqQhwsgnBVd84Hg6CLufzijVUf80K/z+b3+kBaqsoZ
Ba6xU/2u+rsWgqpTt5WdtNDdXRiwBKx4CA7mRB2RJdmOoXbPoU+fkHlf+Q+6nb6J
3+Q4gbvVJUlge0OR889exTBxC3RYLuC7mvquT6zhiZIKTdZp8WWRgEyXOhqEp1LS
VZ4cgmojqakBnzfgBZslui9ek2sAAIaK02gAiKueHVTZNacTQxcKr9jxHAidftPu
nHjCNJ02frZsWZvLZyr3ebstwMtjC70jq/0CKFtYSd0BB2eiT/qwiCvoMx/t7rsS
Cb7D2bCXI6gdnRsF1irUO8KVqjozzPCwCpPe76cN0dqTWZYtX/XE8SC8mYJw3czR
op/X8GdDDZ4S6rNEFu7dcT2na1qfb956q+hvZsat4mTm+a3ZQSWz/7VaKLCq/n1p
ohDF/N7JboW23qKf9/i4nQ8T0Jffk33DaNu9jtOjSLUgKPFSyxI67TWURvIiMHKG
muK0Ay1IuwPDLKNRuNwoB7H2Kq9GSJT//jBdO/5PFoTcSjmdpaM9/3mPfEnGKboz
jqKKu+JPt2IJHOzsECWXwQQnAXGhXdGFFzi7c6QbbIkmOI4UH9dGsruxiVhWL2yW
ZDL7MPLbNLmeZH2WkGBvTbvxaGx6P1qUV5KhLqUENV0DBDmxTnf2mvmHmoPc8QEN
LzPGoZqjGN9Phe5sbVdwtw818g1t+iR9d0OfInwRJeWVgiGSnAq0NJL6LVLjEdzv
Dz8y/7QdXBRcrZt/+GoBTI3P1r1ZqzluYvVvwAvk6E4uAyE4P80w1TEiWFQ6WJiT
6gdpTRBf3Zjv6uXfJQ/57Dyqq5CBpEUa4USfmxQPq34wDgyLZxxI/joc+4wmj4D8
jCuk9U7TJhieg6oevakE93jR0oXl3dCgVrbpfnXAE0R+t8OH6AaaHEa9PFb5HKIp
7exk48Ka1PdePSswH4aAppORa8awg/SbuikIXgUFQ/w2HkIr9FITfQ+CsjwgVfgZ
U1Styf0Lg/yK4nfIKr/ED1OxyoCYjLwsaL0D1SXzCiWYmtclmeBs4dxUp6bI5gRM
nLFluFbklv/dOyzI7iKWy6bs2Sf1oN8kQjN+lKO6dNLdhh6a0UyWU5Hf8J7Nf+k/
wb5e5kZynIlpjsl/BvySS1QSYJwBdW2uXPM0ykA1xmdKZi19OWUBML+kpiP1t6w7
AhJLIYa2/1sZudbhymHGlXvIoIc1J9xWq7uIRvAk+KGevnEOlV/bkNrX1V/oWspu
NwcX/WBeKs3k98/dyeEdVN9zdxT2DXKSJR/Qzvk6NJnZRJPjKcJ3eCNXT+RPkows
PnoZkbbG/ocuOOy3dhor1ZSmVpG8JKVcpzWe9oLeX7Uuc39tMYXdz7EL1bbA/NcH
zTAKr7+EEsE+JbHSJmgEIDjeRyYx1pSNbjPUW5/MZYOkWZGjyfphQlhpizimxwPy
s7V4N9FD44gCs2kt7kXhveHD28yCOz7CM9YslbyDqWoNnRSyfoqSB03iPTJr9j5Y
KcggVaSysvy0ycThHh3CpKKzSrvZMyeKux+sMSCD/QLeu26ZoNCJpTEPRkxZtF6t
gd1g7ZDtvFD4wUMiZfZ5u9N9w4GYkRmGL8p1hikYnn5p/e00HU3ZcSDoX3tXhdqL
5fAkF+SQQLFs3t62jHGR8mRDcP37Xs93bkpNVfqpakRmfjXYAfftHrudLtNvTZJY
TJAxXpJvimHXVu//6JP+DcAI0yiHPCOsug9MqEziAG/OHg1zVTBDiNMFXD07Z2Bo
n2AThakJFR25VTbCO7eLV3kGNQcWr5rGPDdSTTSTnF5n8tHCkAoxI5S7armosC9D
CUFLphqMX4LY8QxrwHwUIJlE/dCQiAR/GvkOEP1GrbOEJViWU0R2X/ZOUBwjoa7R
YzGQTs6XtJs+Lbhn9xEQ8xXF190zknLC5Mii4/1vNLaK2Ip+PrWDdTx0GMzqVnoT
ms2LO+emp5l0AKn+tmUj37ROKMtSWujpEavO0MO+ha4+Tygz9b/lUqrzZKICqIgY
ZzV+mS77tHaGqxjjcJeUCFvKqqWAnUP+H3ufVofv8C1JwMmiXUQMHLcKhE1rnQ+g
FpeykW67aabnLfLNDxXGMNqOsLYmtBIqZgpZMGM8A9BsRzuIqbCFYGXFi7m3p97W
Owev+IFWsADTZ4Xrcf78Ec1TxkJDQRGUuV41c0i68E+wv+N8cJtunVY4BhIjswnE
CaqXKb7GZe6RDlz8i5e/dKKK91qCN2c8F63fJ+uH3z1KUmA/OXo8Zf7mGEaSzenB
cKj3aUp4+EeSnXi+bOPI6lv/m4P3FjspCzfkj7rltrB0rkd3M4cRC5++0t1ObOyl
BDu2eJhG3zV4E424+E7UXRY7OrSt3FaAp459e84ozu3MDshzUxQsnQf1AF41OUMO
UEbGn8Z7kBoJhhPXeY16Cha2rYjgesheHvDdApprf13z08igrGFituFrJEz421lo
weaHugOrVvbinpcID9o62K8kMNb1xa7GkmKFXUhHNfXBJP8oZzcPGzs0gkpLWfjD
FF7tRbBxITIFghL7nsx0CEmehJAwzevCpWS5Mhq78gijOZSpieIjyiOIGBZLCLaU
bdO19NEoGAsY+/v4scfMtcXm1IIFpRfYVRhtQC88X0QDG2YNcHBnRFI30mnzOhRC
hDbR1W6R0ttyVDJ8Qus7igIEHdeejavJoklzMvTqTHLy7vrxvLNJrAvvZEVr+JzG
fa8beK7P7e/ba85885nxRCgHtf4sbYoooOcw7F7VGOFcvklJoyqbNXXTUv6ukGiB
bc10U4XNlLzAj7SiwhX//oe99hjCE1iFExyrYGKuyHsjTJqufeHvHALIHIEKbFHn
6xjK8O4G1RtWNc/qdPVrnP+n9oqL/6fNmQpQv1xSE6eMOqhGWpnhRoxfU2ZjKoxD
BvFB3hJ06GQ3lpc94aLs/OEEdOxuVw7Nyr0W/ku2PqirYOfFexUmEd7bNOEKBXUi
oYjeSgXq25lep8WI4CzXwRx4kDMcYSmPVLA9OsTA9TpyudW7MYmmQOYG1mawKb8B
zg0zML7p0ferJ8KbI11/QX94mHds20tdT1rgLXaOXUai/Ire6oq4OS7hHneYUgcF
wPDicyQaZKPAMIK7+VDB9OugAAj8bjuHKipT+HFF2Uxp+rUIDeODY2vxKFC0NZoX
zXunHJNEdBoUOyJUUFjOXzIrBx2RLKTO//o9fH9H8JhRpWTYCTkIUaCZ1DnPUspv
gNniWjofX3w/uJcG+dHcMuG8Zpmhm8vPfOsJNaWtX3M31lpEmJeGrksQthNp3n5Y
BKDLeh1TeZrLOYdOiZL+sfCM7gEJ23fbDQBT/hjK52fyh3EGDUsOxcv88Ju66lxd
ZJt6bSL0b62u/2jhieptavyld6ugkZdDJxsNNH0S6JYXYf+WOG7pbNBHEX4VvV5P
yFwYJY37dXRZrkkdx6bjWH3If5gjgxVosVfUOvt21AIJ7Pb/xwiIQdK/OBHxaPW7
4gNMK/KlCYmLxOFJXX3SH1PHIHinlE+LoY+J3SK11cFqEv3mHEG3bQeahr0Cx5U/
7/x2E7DYVBsJHGnQ+nmJ+0FKIDeyaQFKJPej3Rq+NVza+oReleW85nOquMqpwFYz
BL4HoyuDEJ9VlYAx+s47IqF18BuySUdHTYKpqbScZckmkOtWrcpV1UUZXTWtw5ar
F0zstfBZ9BBup22HwjLlnrO3TrwozBCwyqNtGbzex1d+TRA4dn8UeI0lw212YKrA
E6vjxF+1JSailQpX8tCWXYdI0vALXBq3rEe1G2A3iVJLkpEIsebwkxWMCkDIIm6l
apAyEPPnqYDku49DWjzrBnmvBuwOQ6GwQO7Ca/KeF9dJ898bJiNAZLOaOqU0jMZe
Lks9Y2RmY6sZ+72Dsa8s5B4lCs0oLJ3ucBuVo3hEjJtZGGecmqiXV1ONfKSQ1X6f
gig/BgYXKIow6aSJP7d6AW5LJYaEPqQaVCBbypzeAp4mLjQvkN2PGzC7e9AML5kq
PQ8psJ/qDvHxFGw3Mulrda5oZ8MwZZk3whPeNW0eBUoRljguY2tWhh+9S1sV7eSk
jH84uDFhBRz/hQi6mewo9cNP+H5yZG+YyO66ZBCe+6/gf2xCEcW+Clo3gxgQ82eU
I6Yu8qjuUonCNvB7LNi7zFowbGdSUxGwf9VOQmCzjan4a3eFJUm0ZEGiXehk2mZY
GG+3fadpd/mZ/znPAQk/nLqLjkVOhQ1olVaNjd1je5SJsMOblPQor0Aj+6jo2wpB
IzoRoqa43Aj6Em0pmIjLoo1iNp4ZzEXPTNyB5gesHd70PjkmnpZsX1V4z2lEZpcH
qYErq3bWaCCX8iTKk3TjOnCVBhHozJ+cS5/rIUG4r3F2E5XLCAq44GU0cLRwe2ev
ttAcWCq4JdUgaUobHwC0qZn2N1s9a//HuBbzuyfssaUGkzAchsJ+meDDO4HSUPaF
OZCojqoNZyn5DDPoSqxNUXBb6uaueZizcToAGq9fxhZAW173cAOf89xkayEDz+JV
QHTd7SzwCPmVks9tlRK78oUSlEBAsSKvkHOgi4YlrK8HAZEAyF+m+ZcvB0yVGN/+
N+lG646QLb+NkLgYrAdS971/lRueksOtS6Nj0J7yiju2oHlWCn9ssfCpkvEb6pb+
65sY0P+D0N993rOhp1PHz5Slt9p/bjSTpqLdv6aYdQpHLv7+b3Qz1tY0FsqP4JmC
bAN5wCstzc7q5jFGlmnljEvQupHuqW0WMlPY4abRbzMSLecYwvkl6nBW6bkIFhWz
K+6VB4OAyEotDAZfh5QlVGNSEM/rU8wTNbKooAvxL86CfsaxatwKzsVNL7BC3LsC
TONJbVJxcl06lSt/FN0Pq75hiH+qsOdgRwEvo24v9UxTxHecgzeFwdKgHFKtgrLz
zwQAzyANlvIG/JKvBq6lMLfGvgXChM/pH8rivH+3nAXpPaP90w9fKGXFyEoU79b0
90af/pNNEf2KjhSKKxYrKWu4DEl7OS2NpT7fnQ8AFO7hSloFHSer83fhZowVRbKu
SGPxrxbAMmzgWqLMjU6IXl5nbEv5y2vIW7cn9rKC0q0oorwxh5FniOzIhf9f5U+O
vR68fba3bl7iWpvt1L+Pal8qgzrp3ZsJbnTMTPXxNMaeMWK6EznOKRi4/A1NpBGj
dkCXT5bKdDXyDg1h4fYBfwGpYmIOIfLF4dZ1syTr8oOil8gGae9qLcExFP2QTAvl
TZlmsQJKSZnHVHxCkXVFMVDWyCrlItTIznmuuKoH1+VTI3Z4VoiiVfwi+hBWc2p/
w32K7BKKBsIFTPSs8hxVZRPw1qyM8ZJ5ZHFVbVfiniPXXbYqX/uu4sbHru3bbQNW
NLPsD0aSficYMO6QkzNrRIEX6MIOPIqgrMeJnIYJxp/+sS6OZoi1LniU2a8xJuTR
FHnADjfkzWxJQv1sWPC+DvxrPDkGprzxoD5IUXgKQMI/XqzO8ZJGWnfTkqROFjUc
nR67Yv8bBv3nadkb8FT2TBrr6Z1lj7BR/DH3Nu2iqQJfNZSGRr+IwsPu4im2cZ0M
5BpKBRzFbJrv1ZvxIZCjQmu5Khqt4rDhUYRa0MdjzThlfTvZZfIHIsfj/933FqPY
koRwOrsOEy2T1xe+JFhseV82c1C5ebLqxgd3npXydZvapE2flR6ydSajPlyvECgR
9JkyCWSopLgoTmvV6+WzhoRAhyAqLNZdzXcScm+6kQ5BNWIV83PAKY+7HW1vElty
b3qDKKP0PfcErD0aaUUOur1clAGoOA1gWdxJS8gx6suNAZ/MhuvOvSQM112r4feI
Gn9YMIVE5QdLqSdnac/eV6spcYXPLzYjDz+Fh60VFdB5nO6OX+kSMsUCa4tv6bFA
TcRT360RWK+7EB7YpH5+el09QW6Q42r3P7qUZVKWzOOPhPkNla8BL0snDr2pArXx
EzbKgX0LTqySoX16e8NTrDMUDvwLQKUrZw/k5OQUUorsdAuM3PKFf3H4KgTnYRHn
O7gTomxN7Yjdmm/xuu5CbW5XJrR1yg+OdqLTH/fgFte1zWe4RfQQIvZxWaar0/6J
RZ3W6v/BoPXmOuodSoXwMLlmE3DsLjdY0+1XFO7QuuMvhhR7KoBL2UIXkkIJkwYS
WtS5C4P9JF9sC2i2YBnNfiFCvEQOC0KMPugziJslEbXUXZUgpUnwLIIJPmk7TaZh
5pi3e9kGVbTZ9LiMo2kZ2/Ywz7eEuvC58Do8bivhq9lr8hFOvWnzE0eV9EHFO3PO
P9HL35+Ej8sH0Q6vlRDllMfsl0F1wRP9YUcyNU8CEiCTmW0hLAJuq/bv64A/SULx
oqm0LEU+a6DRLmJhcmPLmxUPJCbrjWivo+tXAXR6ATEjA56d96/u3azOF/qGWC1L
itVG2buv4axiVzOmnaQxcCulRxTs5LYzaAIvdTKpVGgnc61vAacYlAuYEUECQSpJ
Yd/PZwUUQW8yn7muWd5jD4BarG29siSJmln7qHT8gu/R+Fa/XZ8odqjdrNd2i5pW
jy2eyvUC8g5ERxb5uC2bQ6bvAiUsGu3MTOf/rbgjFfDdMUus4OCz04Hi7t2NDAnZ
161E2jnKAx76XhpdJEjdPXB2YvnFfgN+5aKrYPBRj8EMxlZtFzMHRvP5FFrDprKF
Zvn91+EDbcKE1j/lN3Z/GdXypExuTPHVHqc+F3kwzcdCtfhOe1oF1X6EZTWC1fa5
TID6L+wjxsUMFkOQs13ZfH4KwzGnXnZL4bPxpf8bKeHYFzu1aM/qebuXUdT6QMxn
qwHnm7cWp8lXwnLPDJTQr6Xmb4UQjdd8C80/Vtha4pmLomkT6GR2LETCNHzvFm1e
kDK7wznsNxBD/EJoRWgZ5qo88nyGrhlr2N6UOxCYROZiHE1H1vmSysSOiXaNmhXQ
R7oxE0sZBhtyEfD7SyIgzKZ4eUybYtwYvYc6cKh31BlOqA/Q7XZF8BO587h4V0Fw
bqSJ8toRRDYswrFbfeYQ4jqJCOPLSoUF9SA984FdwXfgt6r8EeKcTPxnqLBOU92J
sKm3qaJILslU86P7t5dh0TGlFbN5ghCuqqaMbBJfCWjD7Z0azDBzXguBp7gNC7BP
7kQYDoC04A3PBjoU8zNOo9+PeOccy+hizWhhayit6sQnmSxY/mXr2+uaNhjMx9Jk
mNq0Ta9mb5n/CRSHw/p+OHqR0sDoqmn3PZAwlvwN0FLzWvpg37sTF13lcxc1Deba
qiPDTEbZjpET4TEwLJA5RZbbKh9XXBMvmy2ZLY6Cvw5kojn5TbA88lhWVrfhA3wz
4I9y11S7h+3cdaTLZw2ATdX2wAvjfa6nBU16IeneK/Kc9O/J/DcyxC9LZtgnrWEC
t0P2V8+5G72CY6qKK7wHBuRj29hiAub2hLQ4bLp47BBkHsoT4hU/zSzcTh+wAxjZ
guxw2IkwScl8xZ4NktrHEp2XZyF8YlwUZ3ZeoJNDp+YNB8U0+2vgM2aAzTavcZj9
9ULcorFNtER7Iv+KmYHyL1Ufc96zjHGQGMeOJU7Vf6QjFmPmAKSZC5KzT91JJ/np
tz2RAI45H7ob8ZwDiyoxktQyuawhJ0o4IU2HQ+t67Gx+kdBWu6lh8t85I0aaWzXl
jhGVci2/DMFNGe7Stu+maKdUA7l/0nSlnV6QcokyXtVPkvRXFppPsO7uerxRRTDY
aLBIrtRMj5HDKCXmGpaM2gW6Oi1EEg/nVpIMLOtffEu9/9+IzJXab+xM/QTiwwWq
8OlulX+CQFHFFV+pZakru7q7jG70Ix9yDn77ykmegHZHmL/t1TRnytMtnmOr5R6S
+xHya85ii+9nsx2HGFCPmT+DNsNLq4W3oPX1PLZYObulFarHue/E+sYB8Sx6YgbE
MfoWjQI40BWkNV5JDukrWyXggW5x5FSxMP3UVqUeq15nC1ETOl1QsRhPhtwFvYVm
cGDDlTRpHjJ6wSfwhVVLdfC4eKf08sRapkfkZGLJ+pcZopTd3i8t5ip2KCRoFtwN
kYUKEBccybajuScG0zB6ZEw8rIA7szmIb0EbaTPLxIT84EHEKVUCkVE0bSx8/ime
CbnXYeE/W+3xD1YcjjQboMejhm81l14oUFW6AyzxnmcaVXCEXZV322Iv2ytTxD3K
7NVW+Cd+iAmu0Lta1HQL1hC2Az/Qp3wEUHhcfqfjmveTdWW6I89x+bXam5YUuw4E
dO5h9AxAXqIzAe0CUrCY9hADITJnWNqp/3lqXBPqqdDve1oeaQ9N+ipDaP7xUZat
SvsJf/999xxS9EMJS95Wtm04XJ3GzaVXH8foAzaibnYYVwLrf0ZZXRcUYEyLeAoC
vOlHEQUiSHKiJ4rDMy6cthJ9Y2wpHwxC9RUU3YeLoVJ3cbn2vQYZ/eLQyRX162Mi
6FiAnrUU6VlGX8AxTDDtY4p0+CHPgy0QR7Q40q6F0F7oW2uXr8qDzSAdSJEGTPYf
W+aU3en9oe5ydMFoo898T8fRj8G7uQFOFMG1hNePLipjh40L9AJEHURb1XChs1T/
i4XOFrNKoxnK1f0mgnWwCEP6jgf4lqPCxiNwCqKxtxwX301Xyki6JeU24xyneRKx
ncKQHDh6Snh26b0TNntsjMS3FKNjv/NddBb9ZXaPiSt813VA8NHdJrp3RfWdtXsl
In1UZaGXVpd8QZi25kmsZ9mRNhQf5KNe4X86hOam2tOAsCukYVaqlkjnd6Bph1ZS
FTR9uXG/JdaSaVtZW5gFpIquAcigz1pD4Vxh9fgJUVb8gbK11MBol020+JIMhDiL
vhLJI8Z79VCsyPfzqDtANGpm+vpOBgtCKpxoWG8hPaoeVe9F36GKRd9xAg0Y8/09
0eExHuVN2gU5ytmPNrz1kHkK/002zHPbt27F3fGZJ0kvnMmpuJL7swvXCgpBrh+q
9EZOr22gLlIBexPLzr2QlkB9XCmrQTvHKMH83MML8B/69bLW7RgXnFl09pJnA9LS
RbyCxrb8rixLhtQjuyoPSoobrRQHgbRZ7V0cTsTqqsvC2yrZ6Cv73U0+/tmffP0R
4JdffF5O8lILVQufCtLGWzxOw6tsHwf91iMdZ4D/5PnQ/fn4g999EC26KJnB2x0r
U9m1jZsEV4gKl4kPzbQucqSvOEO8i1N0PlZrQuiAndJEQ8PzuuMK0dOpG0G0rViv
J2Wg7qFOi5PUZHi/OWvCBVewzoUO8QUcF8iY9o7zw2YokeRXDYNquimuqS/fjw6M
uj8a9ytebOZXqykOePpCB5rp5EGhDSyFMzygo666s4V2+eQqvnM4WgG0vRxi+OgV
n2x3x/P0iCXKyXnxUpH8G7PFKiSETKkPY0MK+Y4rhoxIM52+IAVMlmB7nvTMqpH5
l8jpdY6v4d1HvV0UT3ecbQhiKBfGUHyt1v6SIXMnf5OpiE2kHIKZxFEWjTt+1Sj0
VYALYkW01Zce872ho30XV5zckxHCWx7t0MQtt4l9qQsipwIEh1nTuwpJ02MzmmgQ
eHwJ1b6ZNnFjjVUgPhXFkyg69tmvTTGQMLcKfMGxKhj/ELvUWqqb6uqx8pEMA9ea
47Dgw/HvXSe6kd8uLScFcE/j3y8A5dwi3fo6QzklYFbOHmuqmpNZ4N4vC37JudtI
VQJ9OWjNjI/cmdRo0O8hSfV659mup03g5sH9oStejz3N1rF9KTqqYgCxUougg3g7
wfGLE1eYu27jCxsx1JBSaj9O4GVb4VdOHsfx+oTIlXGhXknvn5V3+V7Km/UyUygk
Pvg/ccsqv1F4xcL8GaVr346PDwM5hBj90u9vqe0f9zhALYx1mSSXcjV7SFJ9x7UM
aed9r/9M1RlCGVcQhstlgTUSDJLk+C7lEaPfCbp35dcnKFgFWgFT6VhaNcvlVFdj
HMRJzgcLnwJXqlX8Ko77QTl+S2mqbTRUahJwxbq8axwtP6lbfJ8reznlkgxL5QNo
txHkm/jl4gfC1fcZu+1I/Zmn8s+pfYES6SR+XJHEU1XLisTZcOiDMv0IYg0puXmb
uS+1rbU96V77oJVx2Mqqakv98eYJuP8+4OcRTz18vKF0osb/cUcc1QjQL4fLV6mu
291aqcWLaVmE3R537RCrUx6A4IfHx0ECKMiQPQLkeFnbGaPMZ+hiOJz+JOe6s47B
qHNK2M02NLFmyseYJa6e/pcCEgAE09b/ZMyRSeVHuqRNGEVlBLr26j5qDxibSPCH
3tDyE7bmfczbqh8OJxm2DGCjS7iGWuZiQVsxjT/aUIiwCDgHvYjHWXXApvzXRCah
KRwLxxBRCdkx6zu1z4aLpN04kOQ3K5FhoIo6tqyx/PFwWU19cydLgMTEoDWLMRuU
9BxW4oEPRD9n2b5P/GNR+iSsR+k4uXtV5bhkZpPl9EKGs516SToIiOo6x3r4+mDW
CDLrhZ6ZHEJoaUvVOFFiK7qZmygCjTQ8C+cx8L+n1JnThNIn00cWGQAess9/4rKT
yPY2+IqTyt4nkLOhwEH7T6tGLhzbNbYMkpasB0kAKdj1Kw9D8IXpoxTdB0nWzjje
SP3+BNzL0h38H3Tp92mH8LNNKLIxu4fFLl3F5Nq2VIMyxnt6Br9zHRrwrAn9LzI6
oparhC5Z//dMTshYG/OyH4EQ/6h8tyNjAnq9JJ1NHmDMzNEzOS5sblmZ8L0j8tGh
tcw+eM9zbv+/cXQ30jBDvtxn5Td/glJxzeczfAg3Nrd8qqLxzhvZ02/F94iJKD8P
C3jh21jnuYZyF4gHLU3UPjrzpuOl/VJRJPVl5yziPij982NVvtuBXyZCspyls3hH
rTEpNzepTmPMAeZ8oc2acbYQ+J6wpiLbW/2G0shIS2meANGXUCVURj1+TOpaG4IP
AcRDIAEyIfWSjVuIbuvE7oh4WfKkCcAWEN2BjIItqh1ZJ0oEcx6CivbIhSc/ee2O
KGy2qV2CK+qx1bprEGtp3ZDqrKrPjinm3T3twVXUB3TEq054tha3f8IkXJGjDD0k
Z6ekXFkKTGEgPUZmR9pGmCTdiWxFL44lvczFlp6hBkhLGSjRZ05+/Ilb6itKPINX
cyGGBX+HepSHnXDFtqLSIGOow01hBsNKS9BGEghBoM/YD84G5JLGHp8F+11YbBwe
1n78W+bUskw6VifUj7M1JQUbYYkY9w7b/5tj0ujiTTznEjQ31YfhtKA2RMnIqR4N
grWIc2bAn2v7ct/R2I2b8E+e6ARwq2u/R98uAwFiyKzqHlFNQMdJt3evwk7aYcIi
3yEJyzokfVQIEukRSjywXQTTzMwIXSSN439xFSfb0ayeQhkYMc9UMUaQpH1WMPB9
9NR2BI1yBYko7Xw5v08+9AJLA8a9lAlasV3HHxaPGDdn/z7rfmuIUKkmOPklMDF8
YtqB0K+0uluLsCn7Qb3Y6xGtWwwSeI225BtWM6o0zYh4s5rTEQckehoCpB5k87Al
OU1gf54iJmD20vcsBvSPrn6JisKiDeqUzfU/QWfNBe3JiZ9Vuexuq6j8pjD6YVHP
jSq5LV907BsEn+CDn1LmNPwXgrGZMHWqwzlb/TFE/IwrKWT1NVEJ/MEUyMVe784m
gKAujjHYaXFjetOFA7AM01NRBD+x+lSzUf4Wy7Y1mC1AA5htZWbC6bYNrcV+A73I
/e8xIOXGFmVs56Y7GxDuddFe4STmDPQ4PH1QBnYcBFNmprX7aa0WdZuxLVKIkD5r
1HmTOAKmwxhJ6ticRXEyrd4VKW0qcGnZSv000syYNTyFRupabEd6NJLUvvLvZiHt
Wt6qLirIcRIs51MNEeNpU1VeFfQ+tL/mJPmjodjdoKDAbBraNnaxyR+YXwZ0yFy7
PAf4yL0twQ/uSYRSU5rSE2QoUhFVKRecr1WXBnX3kRQkKCldW7igx4DaHdU0REfl
OGucB2ZGs6nymsDjvrS4C2anjHhXkHAcylfLjOgnPTv/YnYTyaCE45k10KRBxhSF
kyJucBjkcYaxBl8IGPuPHXkj1S5kcIjdS9FjiYHDl/dsKPvpOMXLZ7+Kyvu7XLaT
pQVjVNobKeYWd3A/ce18Y+It1TenivziCaGY0ygMC9ipc1gSh6rXyCY8SYIQtqHb
+yjpOjyxclf5IZV0qJshhiA61slVhY3ak9cHeoHIDUZIo6qUJg/z5w+FvQYUXWIr
BIGaR1+uKlFaLBtlFtLgEulVX2N6uJ0w6GNOhOBFR9p4V8S7i5s5lv8Qq5auWA2t
buFuTsW4AGeGjFJYSoZOpMlB4usGuJ0+n0oikJHCwFpXHmwVADr8kINpY1IK/rR+
I6KwNs1SkrjK/hEQjUfib9O3TjuLZj+cwSU0R8RuiHsBMKkTDzIBPIE55KoIhZYB
EgDAhqvhTnTqiUVxNdTKgGaEfXXFMNncew6wVkfyxxSuhidJAjRX1y2NG8tXPcyD
G8ifLiua23rxkHVFR6cq/JMj7CU9UQPnBaKLCOfZFuuGHH5F4N3rInTvTNAtG0lx
RgZ6Gz1M1XK/yvp41vCRXToj0azhXhOIwJ5/rHAuUK2rGR/A34CaG0VgUYXoR/J8
BkmQgoOKGjMBFku+gPE+bw+oIDgy7j1CVtKnnh5630UYe5xtFXYUR8pEaqdK5Ads
fftZdwwW0DcAZyLYwS2dzCKkxPPidfAUaZ9Fvw19TCaf7KuDNjqJrVnhlW3UwdLm
KrVwli/+N0LD9gDdExr8BVgixXN1+PdmoGmmtmTA9W0qGjVVlbRZJ2pciFlkblLP
pB8CvFs1m4KiMKFvl7wCyLioFQULTG1qSfa1sq6RIp5jdgNigmvqxox+ROyE0CQA
cmzMG6mTBa9sELHzjWsQSgutAErswB+JhtqL44h7eqhnjleCc8PI76fZ6JLjH3qy
Vru8euZ+94DHRjeixv7QBYaOaud/bmCgTZG2N3OrQDFBU3+4HygoBDf15YiZGJsb
YRul5Zqg+xVPXIyodJjSOyYf+j95z7fqbfawOstiKFBWsg0JaYm4OAWnTymZ2ohX
0eUr7U3O8Q3NOWeVXaw6AJCR1c/wbz3KilGX6A18OdnPbmVPPptr6bxXoDUcEY8Y
O6MgjzZ4QpYTCd7AUhzTPDdyw2n1Q19GNZ4i9Nk4IB+1wZCSHNPPLFx/4FyG0nxW
EHoAjDgpxE4AKTs86mlCR/GtXyZNTbwpTAGcyw8RfOm9CjURoIiYB1+7cRm/7ChF
ldJ1gsUxumjfbGaJ9DSHvIBW99xVUHIReOLdwD2qigTk51ZTKyE6fj7pmsIgpKkB
Ky8GgRefaTTjoUNEOi/oLWUMr72dIS6r/j3RF9BFJ2H6arNKG+465xw98dd8ktzx
/IcWtE2JHVWk8z1Qbc//tWYD7xO0Upa55uAV2mpP/Kcp2/vJS9F1KYQs2DKRIIwq
Q4T2KtOsAnchvkCSjQD89thyVSKwmzcj/8T4Nvn5/c3ubJHn5aishsk5YqOfubqV
FBAwRizig6ZWds2A/EMoEKOI00XjwR9SThRgajCLqSSeubMX8wwSSJMfDEHXmP1k
Gn6boIxcAMhdWVMHbKPfSPdT80KYi72M5a+7veOy0vB0p5bfjgVPSgukwKwM1+tT
C6hIF//arrUn5wxxKHECYj9JeCGWAqsbfy65IgqM1tDKy8rv7uHqI66F8gUHmCzR
CS/VBS7B6FtAQJYL/l0/GqKyww1Z4STjMkGOQVsuDTsElrFK1JyBE+wchwBfMYJL
Qx7zNRrR6wzBgf1Bk9nkoDn4Mr1xp+Z/7rk9ofR+g7UcWdlQnzhPUHDWISk6NLfr
HiUWGXU6XcWlqvQMt9h0cB4z2Qt5wPndYG2e8+DatCoeZwsMJdBtvTGMpWRg59ye
bV4nXhh0uNv2qAfa9SQa1dc1ZAd6Z4i3ARrrrUyIpisduYz2Mmk+oFMhlg2hbpmS
dCV2iUOXcW9Yg4IiM/gZF+XR6xvPK5eyFWHfT7Ir9JhhS+HNCvbjlggeWIpH6fa7
Hk1hqWypmJGgayJmGELSnBS8Y+xwHW7bxWfJ6aLU5jHY1nuxeEOj2PomiRSoo/t/
uzL91Y042+fdYYpu+6fjTJkXYm4qOXI8KBUYGTJDxLumEdwANlr8nYmuOA5Jf+T6
EHS8DWcxMqPfRmXCCwELG06xLnxqG6e6EeN3ZCnolV0DvGWzio/I7wgO1pieCLAF
HeDTA1iP0i/z62OwZC1Ay/BLky+O0BS7M15z2ciDfEHdCpQDL0BTBFYx9tH/ZqiY
ptPtDnNOuyWa6HpU9bjODl8K6YhVjCa1tYownbmIGGH3TzHGzW+OV3qmAwE/Hpuq
1fhKfp0dPf9a+ugjifR1vPJod4S+DLhjkBY70LRfWlXJOXmdxw94l3yJ0277JDH2
tTL0P/aHzQPG33YQnhKDg/R+bjFrySCu3Se3eawbLiC5E0xWt8pdi5Xi0cyZ355H
pIXrfy1odys8+YDeRSs22v9IK80etGGAuC8UJP4a8G8Fd63a3MbyXxQaQbjSFU3S
RfS/lSG7b+U70omqfgkjrDt8HTk+Qa00or2UYFMrEzP9tzmQrDMrUzyX5pwmpskU
k8A4KPdKq6AdGoPGKxPrQrushQ88vtDzwA38y3Np5bRdfhpDx/3dFjfyWjtWAei1
FuglIawPeccGgAxtYdwmBZd9l016ZAM2kQVgLq/Jds6T01N9lZ0hKGWn1I0xq7t9
nWagMqcRl8qv3c7mbq8J+fyw7lQ1UkR3u/PPeUyIp//gmz9COlw6blSGRUFvVmc6
elSZmM20T1soyrjVZGfxPz2fJtTb00ccHxhJEfQJrSa55PO0X/WF22w7YnUZfMwG
dsSBiVtnNXzpU281gWvPfcUUFTdLLptjcoSxLe1YrQRqYA/Mgb2oJE2SQSmvTWGg
4/e4T5/RwcPlGlXGKHFxEUYIfBQ1diNjCNr3SSDzJNqGyn0URBGDDQK2XMqUEkDu
KMw4+tMmdDuENWi//i4MzKIsKCNWWLqu3wTRLl/m1oX0W/hTKaeo7SX9DNkUqEOT
69Ni1JvobtYeFqCr4yeKhhtspUS5mnQkKHcxk8U1w8Wmdou7HGwoeXz2bd0XUOC3
uNwS7J1s5BA2fdLz4Qh7c1ukCqc1fQEBJHzex/CHKwxB+KeQ6aDxmt9Yxk/he7F1
+wtMON5RKBrotoSqJIWH6ny7udfhWQEkGZK4iV/q13d9Tw1wfkEcVpR6B1QmdGMQ
uT4qXNF59kzFMW+nrIZTfIWkbbzB7Mc8qQb8ksq8BjNze1BdvMUYUElQcmNoqIBk
4bT3XOH5gEKZewX81iEh5XGUKiWZDb0mYM8S4LTkqib0jXah/48vp7miNUp3YQQ5
nKVIHxJi6ZQxc/hAaWBf3jYt6GVW5+tjwqvpELfrxAogm3ldvDd94c5ClL7rPZpb
IzKt7BDZss3FXwiKXrjRpd+JLBnsnPKcm3dgrWzrpcDPEB2mMuNMb2jrbXiCj/BD
laGyvK37NrhiQOwMjpT4trlBKF3izsRiqMHXdx0rHjsSGn/NgtdmH/DKnCei7h+f
yg7GP3lEFjs11RixOAv3CGTLd6V0PhkMvE2Pm67h5au2FNepIpH5miMX16xisB9X
g39HijX/l/ZFTJvLeZrmCpdBMDJskCYizwBwNQGy4+0xGXjEvaYzoFLk+bqdZhHY
S50LLfjb0oSROLKwKEQU58N+mMCA8YZdnpdeHH+tXwjpCcTbza1DjctxXyfAtG8j
f4R7Ev+QWda5ASvmbTu7nHHJgJxiJCMUWzR4kt0sHR0RJilYJvfhJpMFI23GWwpu
tC5bV2LOyS1nroXw8EAPtiQM8PcLYufH6Pv52cja2qRWexUhKRi+iTwxeccarpOS
4AyMnBN4eSFWg/R+bDdhk+2Q7AQjKVmZNyCPlZL33bogvrEsvYT/QT0V8KOPXatI
/HJotYeOFITO/cidjB1gzgZ1SH1bDmPT9HVfNd0XmFnnA2ErOnnfx1TpzcEOFIH9
0cOgXJOF/7HYy0u3+7Qpo8Kpd6gcEgE3dp7DKhz53VOD7oSdXjNgLrLj6ZDRddML
jdWIB0yQ/BO3j8O138Q4eB20NDCPQ49BBkgQ8RLWj9hldsPeWdfGBf+HPTYqYil1
4Kfbco4DNAjVB8GaymCHa65AQOEiPeBpwdt9Y8VsATwRbxM0DJrhKsR/l26zZH8j
x9b5zTQ0Z+Ms/yBoRTp5Z4E+sih1CPkg6zV05dCnDQepjMJL+Ig/finXRU/uc78r
qCq3n0IROYFEaavjv50atnCQXpAWCUwWzVWn8QvXHhK9i6WYFGsOcv4SpyvKxi9m
crPB+UL1GWI0Hug/tTjWPR6GmCwIqBZp91it991wJrsvtHASNajUN8utF+LrQXDX
4jD7gtGS73vHXINKs+MPW6fmyH2KJJPXrc8lGExn9Ezay7CKlU7YBLF+HAUn3s4w
4/zyRJSavAKCOe+2s/2s8YSqAjYqD55O+6vySAS68nF4n93nxsyqNZWcrSVHj8pm
WZsZjS34xS57JRqRbyoPUozosGVyhkdr7kGITdJcLc8cDjFvzl/7D8/xL65breMC
5CW2rfj4ilzOEYD9mX/36akUCb4Zi/rrMfoEkTtfTwt3mskLWAGLkXraCYWuBdoO
0fr5wxrg4cfxwVGKNaZwn10mC9TflHFGdLUPBJuaD80rXir1VGFTztX8CwDub+uN
9TKWpgDcHaL9kNxJtLfsBpN7mZfvLkQpelP0GO5RFGhSlxz+91qunpnxkcPkLe9o
lFQSdLYfg8ynXblJxnR2pPTyEc1Ic1SNd+gZcAcz79AHgj7e6AAHfOV5Bm4uIaxu
XWZTrUywCbxzPPqBb7Kg22sDc1RfDm3QAx26ku8bEx4eYudUfie/6LVAB/YO0kRA
U9pJrhaVWRNbWU8zGtGssGGumr/+zUEI0cmMLlNZEiPUYS8HLLR/Blh0ScXh4zRh
567nQTnjAZYuCi5ifpR2P035GQcJ2eUM4zVrvx1nhOjwM5SmNCD92E0WKdiQq7iJ
AIYoW62d1ETy20MqiRDwMdZrCX1ntXu2AsxrcLGlpAbT2YmIuSygciXGPWj1P2Tj
88vPOAy/LZqHx+vSfQdhCO2itIn+LCl0vAZ5iw3Ve8bXDwJt0XcyiCDE6CjZv+XJ
SarHF6lu/iGQmyzr0VdrbUs3PIcA0aKGmCUBB2sxu03zv/p/05xWqTBytqblY0Nb
C1DstdvvgVhqeniK+5vl5eXRgzIrjXyoylrYR30Oi8iVs6C0jwTTSVmSOY+ecYFY
riY4J0jJosLg1QCokMMEDdBg3gPJY7YhzRUhXc/Wf7yrruEcpbMIlp7hUd2FS1A6
MrratfG31ndOZjhwmvISGrHQRDFFM1krrPhpXW+ZBZ+rjwB+0sQj+JOedF9Wgsry
y+K4hsxtSpqh0em51JN7oWghspN6d+u6jPaQ4GzNZezuG5J+KFSjQi8QyykwVO1y
GnWXZRiJOOnxGSeuFoMzzzWU9fjD3CGGa+1UPnTD4LIuY/oBoFwNM0mm8T4JFvXt
VrqpcGQrN6j/gANXU9ngtyKpJZoiqZo291a7vnjzFjjsGAHJBQ9pAwebjH7ph40j
V/TJE87VB/8+sXUSX2G1GdBb5QFMFGi4m8Kf6KhJXO8SgxPxVNFZxfx6I+8nviz3
vj9AuElBtDB4s95CJnsri8aetTw3L4YQmtQ46XliNyQ8csnwPpgzZgY2SgjYArLQ
4Gr2PSmfbOOAPebDRpmVCUQNSIjBYvNs4NQXUbmBEwFnwungY88U18UPar24Vwss
6Za+G5VGVsbXdWW0WDwplgbCWD5+65ht+IkxNR2mBDY/CP4D7KE8x9o8uS4RhgX8
1ilp6+ez8HuAol2ygDXbRt5AWlSuZz/vxfRnrQG8Zwd/cW6kdfEIeVCKtdCz5pNL
Cww6s5TP3ytDR7vq6aCSsc6A7KYwjFpJaOOVDqGtmpbGb5ax1FIB77pSnCUdMnV2
N847hPJysRqZ1MXAtCSFd06xLC35u4RpUIzf8L7HXGS9rNufwg+Yb7EAQsjtGuTS
53cAq78qTLITlyc0EqM8PsXn0G9jImFPLSVnO2HwiMyKELySlqD2avG6rkSAmGh9
I6CVtAxG8BYnHc4SW9wC8zT2TNFnDRNuSetmAyvDHyOHVnQe0MOLwbnZVaDfZKJ9
b9AkuaghV61PXbCMwdhlK7KA1JoMKvl5ug9TDKjcOg3aIW81r2n+fjCzJ8gIzfo1
gQ07cKjOLSDVpJXXUlrjZbbS1NT/mMiupYvD9UeN3Sd6PtJkIyzbEzP9BnwOA+bT
Qu0MZLKg1ZCeGwreSANGtOxwPv+koUCUi9b19BJtIE2yBMw8paIJMQssoQXYBSvA
WfNJfK5UrjKWUV0WxrS0XHE+f2vDSQK2vH841NymWq+NBGkfCf0mNfZHfwi8Vacp
64n2LB5HuCmOSX+UTMWwZGOSOXPCjU9spBdpc4c0pLgrdCv0gFVHDxXKnkEkNTD4
YB45qeCm0QiIm7stug5J8cmeAgVhpPv6yuJ1BOyjDgb5ZeDAbHNDuEMcPv1DbzqD
iLEVZDF/1rK5DGvjZy5tyLHnrA17mIXejmDRJwXmjv74RfhnKuLanYi2/VR67Wwl
2mWXGcbYw1GJUIVu6b52g6QVN7lC0MBQSVGUqMj2BtsiMkiOuUx7PUU7f4tb+VOJ
5zVWrDjU9/Ek476eaAfj6jEBRJASksN1HZ31YY6TEQ8XnmP3OOUnD+YdVJRtMOjv
gnS5ljlqhmHu0FnnGBmITwv0uTJMtSoNUiuIUSGXKVW0Nu1E2QL1twmSm0QplaOD
HuAb1VOpI7YjlX/ugTauw/9NpmA3Nj3oK1t0wr+WAjLf50FfVenzji7SPYZsAOcU
tUVwtEcwS0yTDjbhB6hq+2RVwsunZ6t1PB4E4SVEhqOQbNLxbGwIYyvCrSqFWy4y
1Wdvh2gduPFxSE4fZUhENZ0lAM73Q2J/Be0nPJMT7d+xC9uEW8QYDblFIzjIW1aD
IpztDbI9j1Tk486t+v0JDUKA3eb597lu6svgCL7wMCsHpiSdTQqV+7izyXAax43F
EQd365mjfqHxVLAj+bs3oX06ouME+SlF9ycRNb37a/EsG+El0329jZNHHGZ7dSKE
IKMid+CIAOxOdmZIAflvmJvpH0TBnd5AO+4YlazRk4YTHnX40igours1PfOD7Xl3
WcXjwa+Syie/CqrOdEu6GxiykyPZeYOXzIxL1vHE4Y6PQPbx6/x2FRNWNk2H1oNA
jT8E30Ph1zf4t1ZTdeNCsRqKl6/TcprF5OMwv4rBnWoSR+UupPFl65XyqDsXf7Pt
ms6BE9NCM8i/CUoIHn9InRXKDKR7KDsin/AA7aZF4KHl0NPg6fRxatLPbE27ma3o
j75hjbPbyxdS/7ewhX85G6aiIxeZH28ZTMFvjbz8bsa6iiUl10rfpdlwJ6Beufqk
7O/nBb7wtywSQDy1HwKoHrE3HJB/UYxXcM/efy7hZfehc7qpPkTE6mR7cqvwNT6E
BEpqNIoiLDikEwZHLTRF/Xf6TtQXryARrqBQWg+xHMpQQPMVNZTF3U9/MRhwaj8i
SpsF8hgMLvNWlPpfMNgKCi5DM4rnwhEgPpQwFolUbqr8CovY4PWsdejCJA85I9de
ANRSVu4JKlj1ln42fUVAWTD0S9fg4Ngz4r9ikOzc4A9UZPbGjnW/WHx9Rw2DYPPX
oIyC6asouLpPA+KaJAkhpzbv4rS21jxRpmHg9asFFojgITp5A2Y5YLMH4t9nyF7H
c3qiy4KPm74o3SCu88hRrz05JOqTCARKj7K8L2UXQyam2TQNwxyfzK++ZdeeZeLT
h93KgPqksVIJj1jbEiy8lPwFbtEEAzyL4RQ+8jY00FOG5dp7eM/7Zwmb5OD0aDh5
qFk34VZtSfjBxm2Favn3mnW1a7Vf061YBh3ANzl3V3JoHmp6p936KmwfEJcSH7ld
GEqc9JCMTiTX4cSRCnRBJzBEjKAluWXUjLHGTRuAYcxkm05OZ+6PNFymEKhUeOee
oxQ22SB+w6id4VcJOuGU5I609RlVPWEAwU5mq9aSAKT3T8S6P25n/jLXwsjKtCD9
QcBdanbJ+KY+7RLY/pyeOOv+oqX5rnUy1owJ1HvW89LYz00hDwLuGwuTIXk+evF+
0+CM+/i0T2053WrWqcveN4cd+orMlWvGmITo2EIxY+WfRZB7wpZioYqRCpBudz6D
xzfYkX2uyzxbQXwm5moJGn/okbLx93XDUehqMJ97zhc469emMRroCBBmjOTg9Rjl
A22LhhaPgiEAVOsNGMO2kKqei9RbTNUBZftNuGYuWAUG7jIoZMtQamq9Yzejbc5D
JqNTdRnGXafrWlyvw69xANlW++dAf8OqKBxPtkF9LPTu7LbqCTw/kc859pPdr1tz
PvGh88Y3OMiq6S4/Tjf5Quvwy0srDZv+ax+e3vcch6Hb10jNxJFWsZmaWDl5vNo7
IJSdDpgVM3y+yCAzQz4iX3sntWDl8ZNhuOMOMlctB0LuUE8LfBbrQexxaj7ixZ3C
7scHuB8SVJytlRJYrXgbZJWIQ29a+JO/2Icrx9XBXP4wEQSeBqKHz0FaB26PT2vq
XMHbU9VRF4uRInh80qaSQCKH3aOVrS/MO4P0VnFjsPH0mlEe7p9XL3WWLZeW4ohe
4fBhEShXA05eXyVF/rkYNtL7l8oYy0ooVL1/UUQrQf3G1mbaB1Prlci0RPTLFaSc
xJDepnKvY3lB81DHaEX2clB/QF+YZNRiyyJ55tozVBs2P4LFQe/3VlvUOr47HmDw
LbPgA63IwawVIx7gjN/FYFW+fgWkaKTNiuBTBL9d2XkM9FFowDOolNMXkW70fPNG
BAl3ypzrt6Q8ln0n3vP/YZGflCa3SgViphYalHfaQy1X5VR6zteCmwDfbYbH5DJd
Mgy1KbX5osW0QTQ2iuUyMxkhIv2JwIdsSZc0KuzMZ2sf7C/TP6icY0AcySOx9vRy
MBAqSfoCl2wX2hfNIe445PBR7z1dy5o55AOGp1NKBee/NzUdAv6pW3aT9lRv/Rou
XnwgLTu+CNraLN7QfympS8seJJep0xV8mbISbknVAYrwuRciMSrlvGVdAeCbL0ra
AnCnGw2J9CS9+xCyg7BTsaqUN3Ep7jU18q7rSP1VruPmOHnwGeCqn6gVD+uvpBAb
mfR3hnpmm6fgndBXetkb+Ayr8am+oN9N+ociS62rvq2sbAsXFXSmrAwYqQjPI11V
2Ao2BlSUi6jKVOhSeJWzP49Pv9wa9o9dFahnoKRRSDXmPcmPkUjWdRJM175AOM9C
B1/vj1pSvWnPak2DZOdKqe0fYIzEuWfhiXNdlTw24QKKeAG6GeD/33a0+rmp67qA
LjDBrAjmdB+z1oy4qIuFVpLcZQ+MjVt5fFleVNCVQSeZV4r/Gvg7Mp7ipHZrxORl
L4l9gC5ZB9ct8LI+MUPbxITfNDM+rhdXKGLonN/pMQduL6W3cPiPNBVR9NEUdE86
rhQ4YwIS5Ok0owKeaOODmonSMq2QfaXEypE2VUiCeFfucIQdKgDvJ7dXTlSeijW2
i9ardBIr77qkxhF3De0RfMFYvXqAXCbt00n2S5qp08xzSZNis+nfT5yF0zEBxEYT
TafmT30CWWh55XooOsZa3rDm8T7BUl3EZceGG6AA4s88SeIwsfmMdQ827yWFGHW1
fApaeFcxckfgFDzUK3jxSviugZZG+AJjKjFRUvlzDPYLzL49vhHH7yjSIYQWpCWH
DKXfPdFn4fJ5Zp0m/Yvkt4YKuJmvZ0yzO9mBaZHi2Cw1cdOzDgmZPZq5mV+5MmFo
7yeHZU2C7oLPhY4tah3M7fC3zW6ya/u4rPm0iS9ZCoHvLmrqR0UcX8dzkBfSCvCq
CSUJ36n7ffWbfucATLPgOufHsBQiMXG6o0VTJGGaFhxYCpU/VDgwt2P8PrY/SyRC
Y43ztfdh0AThBEQs0HZmq/u996EAYNgdsEx+7Lg5BQAAWRLANwS8IhT87Tze9wJB
7MLEpz9B+F19FFW8p1YBMAi5R7zXax60IWt1E0kfb0qZzubtUk9uQf9ThINhG+mr
kH1OBAUwVsK1A96bXIc2scXzY/aSUrQ8b7U2vaWYgZP3aKzcq0tCsadiaK5ngMG2
MvQ2wz1tIMx7XFmhKOTRmXKJXZ2KHnsYu8ngWhb/IRTEJ3+5JiZXp5sApCVS2N1U
fe3eMu05VVhk/jMbxw4kAmFFInpj0WNpf9XWalCjvkcjIQDqahbvLK8XdsvNo+9P
aRxQlqwA6HS+ewqOIWzF7xmf3zzL4fEMPbKX+4He6Rb8ozqlWkypxkzqjFiwKRlG
vfYh9v8PK7W85rL6CrIQaCaytjPf1rD6D5bRu2+w2JEzmZsYC/bwasPEXHCfZKkq
y24FG/7UNdOnq1tOYKy8Qrigx6XnHiIFNV63jMFjKwkqGJHohSyZp8bXd+hBaNCR
kXLMgdM4C1iBKM/XIpj9SIQNCgs18ql9JzZLLLU7MC2HpZSy5QJ73uskwWAKjwqe
WXKb0Givc1emKzPmnrsNce6cUpKMHtIHVSMZyBgebNnEkCaxxd2CZQV0KNydyZQy
2UndeS0lQt2Niz0f+pbLNsDhN9jwk6n644L8T0hUoFd29sBBui9OdV1hWICNKVrU
g+c5PwZEi40P39moYpjDlLQu4wZ05yaP/r17Uxs/6G4tUxp1fegHXcnZUPx8Fy/6
AojaP2zjnf122imJVj5ddGPhVJM/y74/p6ZOekIxm5CMtMvnsaXMF1fARtl58F19
jTCqxYHjqH54RKnAE0zQiRkoYFADyiuYktVRs8tcTNj5X2rPV9fBDHblWnvk2be/
jJGKI/O/KRnQq6q0W/t5oiAO/qYeiGpEhwHpzEUcgpusx/t+Twq2NLJhPaW1U3ey
2oPIwQvngMAKoogPQbwM3704QeGiGSgEqPpWm0btC0/u29XZY13sF3i3/Kl39qgX
8xx+Nh/CXhFiObIf9W9PbnuOm3d6v4ElADIB3ik97/FxL+aXsNU8iMeAgBB0k2U8
Ig/EZ/8cm4lkNs31LKZ5HKDV0J7H2OFqanBV2zWUCnZGQ6RJvPOT+aD9NxgIwg1A
uipsCwoWK3A3J4SkwUN6bnjt9H4th1211oqDnEo2fYXcNsH7nBsCXcbBEbI7uNdn
0FbXUm94KVKl5cqsIhcy2HUtDZK0cYGm1cGRR1NDjbJ7wGumjxJ6uXboimM9VIv0
4zqIpSNzAAZFX5bfcFEpXi5tR8hVYOf+RIsIlqWoEkmKPqZoV0SkHRT2Mk3+nwVd
lXPECHq7zySIXen0mzkvEYjeZC5hGasKasOdFq/7lshme45rgWpk/6oODqNq8oPT
NedqypSF8BWu660LyzqGp8oUnK4ow6J+pZSsJtRtFZtah8q1VW3C9EUH62wBPavW
6clM7rPXQscqQ1LfdrPY2du5PGIJDiswRxELmxodkXg8Go+7TNJo0bcWzfk/F4/u
7jEiLWiniFqhbhVJi271H2MGIIe4T6PxKgwtzmF0BVPd+p3CDggHSY3/v6/TSYlE
GXfgPAVFbuC/yfmbGl5hBFK21idRUgT0E7bFZEGQZPV4bG15v2ZIe8krqHoJWpSu
0H8apNaeOZRu7A3haitACtPdic1aX3xuBHDotCZVkMGsb5Ey7XGLTltcOPRtur7q
IgDWBCsyRggxLRz+r8zQNObbs8jEIs8oOeVwkepl42YMVgD2qp0xXjDWclVA0cQp
Odn0hinq/dhjcTBCuSPthBE/8HxYOGko551UfPbOlPVx0qKwe/Aq5xCNHfaXnPhH
nXz+FpEzuhbM3Fx/Rig0THFMKll2NnY1WZpndO9mSKUDfXMUl8CD427O+Pe7Y8ew
Qzkd/gnIEMdpzEvm5gtbBoTu6MfnUlA635dBpVCqOJumUbrNMAXuC98tBYcGt9fL
6I2WjjNKFLNdEUozvL4z6XBzYl7ro1a9OnpOR84wOt7ub1bAFrjYRb1CStDzAOeM
4Ev0ycz0ql5GxlvkiNxbUiKy4mR6hRuBNjKUCmVpj4nbNsNLjhVsm+ZkPnwSfMC5
5p0PON+aWRkxNLIG4E4xcU3MG8zwf1zK0+PdIf5jsriIUA5p6A+R/yPFlJNOi4cR
y6TxME8EthNceANJX9lsZzRtMlPUEKnCq135wsBIZpTeT88n5Rf5SGCPQyl1td/U
XT0YyQSEIgj9nrkLvi8krOMS7JzZHDLIi80toPBRYuVSQ0RBKcHKtydjN7ewj233
46gNH5ojYl0qL28eB3jQoVeKqscCBM71hV++KpqjBZOGiqqF2sOxUhP8mYu9n4G6
uHCtTAUGpS3LXce2kR7tvreWTOdaMw19YipgzUwZgty8NrhFc9AYoURagd5VRYnS
G7uQQrW295pOMClvPr1IBwzr8xcyVvLAdOIAClCsSKPoOcC3VGgOs9f2BrUBhyDO
2Q51LN2ul4zgL4hZEpwz0gI4U5YlfO9SDbQw3lBfF+DwLEbB9bFRuTcsk5xYDnn6
7De2axLyn8k5t8O8xkbYmvPkmUP8ArIHpHbuye0Nuespo1Z1AT46G0wVF5y/1vlT
eRG13ggOEXpDqBT31MI3KxcJZGTu//68yY8edAQnrU/ktb/NDS9q3d66z6lcjDec
vpnMk8rL+WLGHAlpRD8WsZ6Y8pSdMi2yCuQOlrjXmFciIrjNVaffz9Zzf8TpYHsR
QQAxd0cesHi546PpLKIz1qNXVJIBHNvvDuuoaO1TqvrcnTIx87x1+ICCI2Oik2Df
pax5vBD0WtGaawellcu3TH3V4Cu/USSi1OEIs81bDBCOrMMGOd3SmPIgwl2rf43j
Y2zfEwCb3UJlWtuNRw5s8Gv4Arwe4KWrJaufIeuFELxivB8+vUadD+EeNMZqVJS/
SZ/v/GDPK0T/wituBPm+qtl1QMCwLl2tCrWYA6I5l+e9S9ZLUF3rcyJcp/VC+tx7
pAZkt6xE6/ioi7MFovNm39cXhXa7U4AnlBYDnKe7/J1e0eZpQnogCevaQs4aH4Wa
M86lLk916nJR1W77mf+HUOGMcVrVH680HzYk29k5cLMevU+/VF3FU5sl9PsfX8zU
y22S0PspQHa/Lj1GbkZvnNHS5/YGefmd7WFLPKwzcZINU8/xLoXwXoTJdypC3yil
azQDUDfEzqe/fcoyie0ydbho7G/Wz5+Rwgf5gDKL+5zGQpH9GkcwKPzhHu3WtVp8
O3IH7SqPELKpBJAWF5LiqizMDPWeZKW2tjikXQSUd3FKW3D2VlGdRI251e5MZVXO
A88R2MSajSVdWH1Q/1z1y8X6KpEDRgolX+7fX1kR+33r5we7x+MC68uWgW2V6aPy
5b4UDG5vpuWRMzmJBE5Drn5k7FMlYI0c9m6f9TAewRo2/X9YiRVzeD+rImJ7ceZl
K4R6T27SUFK6Q/tCbfsvnARwPrfQEcP9/w43N7KeIxVRcrlMo+CVUOfQXUOiUVMd
R7PaL5VFVop9f0f2zee8zZq5hY43dTAExNhGtzlJVCX3rqL9zxR5RaQypu8UW+g3
c1cu+goZ6Df5G/XBEOGVI1c/9bxpalje7iQmoQMD9pusbfh6T8CbXEjkP8C1LZNK
fm2q3DS8F/Llyny6WRvhJK4SfHsqcXFXkDLvvX07QfvQPkEzHVAisySpQbbAijcb
62lrb/6vxbGpR8l6hW1xShJE9A+M6VvvD7G7f71F4jXDOIv1cz3iBSA2jzrF1tXk
Z4YdqvpRPjZgiP8N8WnHSdsfGJsIKzztGc3G0XEdJnblnEyjSBgqv9hqP1rJLj06
z10uX4UVHk5hHphJcKGiuVr4X9S/r3p4UdrxYmqC8O6CmLIJPw0DFkI+Tv7q+Fpj
ik7JbumTrlE8/9sF2StccxJXYwjL7I5McLa7qJmHJvYi3rfkmgNrcC7Y0r43YNAu
KFzdu5Ib0q8LwXTWFQ1amL1d9LF6M+b/5WxbrXHNsRNSB00fSNVu7NkH1U20sJrk
g4TpNjKJealpLK1iEaA4gSOewbO+RbW49swFsRmkiamUhAKP+KlxXEa0+ToLytJk
nbQL8LDINrJDEdjxki/fVOTWzvARqKGO6XclrHZBPU9BRWyCAIycynaL2nZQWZyW
65x6m6HgvwDd3cXKHGAe1v71vU2lMZD4LVAO7rEHleArsDk3GiUPh0Jxa6Uh/lP+
CtXt2iI88tT1dIBqrH8i4ObVz0n0HBXyxyWGeHCwS5CA9mmoA8OaLbCfmUZ/gDrR
SKaUxfLZel2CWdVBk32eKnv7teDs1ycW1rkIU9KEx4AeK838m61XZXhd60jxv5TW
zY+CDqYMnVngtFl1DtqsS0V66AyX+cSC+PJc/71qqk598p92qv6Tp7PmQ99wTERI
HlC6NwFICvACndPajnM3nIOPixNGtCHtuOJiF1mcpJaCjcxjbHVGeM2PuU53riho
T26yqNxKtHJ28+YCKlkndkTmmWuqsLQzsBxiif4/lgws/b29i5DZ2l8okUxLjWS6
V7VNaBXA4SnKiDqNX+VENGxGO37vaGAt/AR+qbLdjHnwKaZ1gGOv+Nwb0DXyDeQi
jfwb4stJj0sedSezQ8REC9U65jVIKQayWAM66sA96Ugv+ij6u6DdZITOfCGPhksw
KLyADEzQcP3V8ABsYSaR1SUfIgkKbh0bp6DVh/o+Opw1xjGdzOJWcP3/ud6eHOfi
CNx9quO2kAxpo9nyewnkeSkG0oeWD8QzYIqIGWnmlTRCtGgqc/isbEIIy2SG6C93
rzfonb3RvCWV3oZvfymhXzSDQJurDPznTZCngkzMfrUrRlwDgXrrO6z8ZXaBL7T4
s2PUVmrKOutrF6DgDacsjhEzqHPxnAsxc2bt3KAxTHApDCBXIw7ktt47n5Pnd/VS
ej/adtSLPc/pBPy8JMMR4oLCgH2kWByM75IcRewlsjiE73ZUPnZUoJ4KYXVXwVeo
mDWtEFGFD4QZ+Fe8JCETbkwgBTesu2PlZFmU7u72wDCGPd5Tbxf86KJvSiDd/v4+
IKRjqTp07uOkaaxOcy7GsqbehDi/nmKdXiJicGMjOzPpxrJefs6l/f9sC1mXU3bQ
leskMoIdOwptPN+GQv4CGqbT/QkvHYHtKGcpu2mYs6RKXzbobbBFLMM9SOK1Sgnl
rq8BnUoVCVaP9LjolYuCEFQ90toIfaFp/vn/gMI1xhDai+8MmHndLb+PSm10aq4N
lVgxOnEdrdtDNXVpwrx+fLWokzoRXWTtFFUefLdQOE0G2SV7+3gtp/SkNDOobNU/
rynCCSfBq1fVhmucySUBhMi5qa+Dxd8qQkinnAhJTeanV1Rh3HQ73YteexOuqBeg
gjljc2kecK4V+NmzslOgOi9emgd0Vi3OeAnUIJFIZyUYJmqXM/xmNptlrHFP/t7Y
fO0pITVmtwYU396Reho7sBNnZOsqIEmZCMBi76gTFiXvS1MJ6dnKWQidMgnHgQ4d
cAUDqIn5HAwLnqP7PrAq0fbHXrC4TicWwqoq+jvkF1JBigKL9ZbQWTONXdVYKHEO
UCFbq1HUo7bqEk3Y8NAuZ85RL3PpaNiO9+5M83E0VPil+MSLrILb/nNAXuW+X6qI
zNO6QCfwQuVBr4BrWwVR0qpUj2VNUFsPhAjJDOfUIMhMPuv87KpoaIPdo+hz+rlz
kfjcBnqIbWIVZjKHB38xI6fPjpB9cACzX0gDxGxYNqVYy31mEcBBOUhE8ivJxXvg
/kKppihKYPgQx0IVz73bcQLSRGSA2UIqt86HLQQE3CygyUajPEnvhj8+XSqgmLfL
lyu+L8aYQgk8GENru6R4jyuDHEp1cXRn67G8C9l9m5OrxRw6gw4pcOS0+rIdUreS
j0lEbZU3RqkEyW0Uje2uhxsMjsz/5WyrUBZdVt+JDysDRbzQq1arrafvltKB8jWq
z0CyvxR1IJmwBIfZt5ihFDl23Omx9PZan6sI2AhSBqLHPdpNh/2JHDdxw2ZQwmnq
cPpI11L9G35s+EOyTwhosRt+LKvD3zGK+e4T6PT7rN4G//lOAXNixPSNLU53Zoov
EudEJxxXt1BhAyKN+4zas+QkZjntVgA08EhImCdQFkMlcYm++nY41BM/eyFuqEQf
zI1n0737JnbpxFNkkuolUHKVl0QvreQPkkufKdVeJsMWpHw4DIsrbf/P3ydFSQWA
fx0jEtPvwkFVV6YuiZW5QXkZCueflaZJcxYyGJFlzq4YcmNXdgqmopC2TX4kDpf+
hySDUWMqt8ShY9w+mijgXwbNKqfrdUo2DDNU1x7eAY7X+keV3aTf8AYetvjUFTD8
rdg0frcoOjf44cKEX2wmf9BiOKtKR8+KYS2xUMljKp3xOjh1/1qz1NIxhav1qb6u
iNUZeh/4E7RGeKAznNoYpNgdgJ2AsnoeJF/l5AncreHf3Mu9uYNOfzYsuPwlbBWB
MIEPax1Y/n+ZWzeexlqtpmsXk8gOogcwzGT0RIRsOBMEFSvPueyfcQhD1gq5kcXy
u/kzn25QnaqRy8nmPg+mvwgwtc8DWtiAsxzXRwnFviAZMRy8dTeGqjMGzX4eamto
C4iEmTlsWujVnX3WL+vZZdpX5SkOx481os9eC4xDQKil6zrjx2F7F7fPDvSjIYYk
jp95H68RRuZpFlpmhmC/51TakOknyIvKou1xCZUNGAIpH+/X7ZKZ6HWtqpZOXVB+
XkxUmTdLEsddPlzIt61KGw9zdE9D+QUXhTXjTOhyExM+O2Cr2LFFZK93vYiYkcwg
FX/gn/crw7vgTDna5gF/eCyTadQHpZtZ5aIIpsNT9SNaw+KgITJfzGcJ/bnG6twg
ZmbnzTBxa4Mnzq4j1c89BuFwM1pu7ch3no7mkc6uJa7PeGjidunabU7shVKxXeH5
NUgYYveecFZDSXv5EWSA4gIrY5MG8ETGAjnUUfgDcbJUuiu9A0rUYkcViQOKqIMZ
dSPAH6agMPCbc1eeigWHFWAcEHYJ2nL2StQG/Bz02mtRfS9UG4YS5MuIJItWrIGl
h7DCZA86gWBNl6Ys+Zvomb0ZNta1EW3olgxvfe9zujaqq8msCmR9szmmh+Z+y3tG
fpUEK7h8/f6dEZNdPG/8+Xwp9kkz99EI/es1uTh2EVRE1706fGZYmWFwJfbePP7H
0/li4T4daxUcUgEjp/SQGtQ+NeKNScU2hbX8X4ijvFTDdYa4eVt5qqdr08Mwvn9t
3/HRGfE9wC8CYNcWSZ8OQlaZcKLX7jXgwL/MECtpHMkDqY53RpvghAru08IQK+Pw
xb+NptAYjvHr9EhzHv52kD0u66S16Ctqc2BlPyP1HeuX5RvVkVdeI/+2QEG6uvrw
BscW5u66C9h94mMItsYBNyGdTE8K8kxBgrxhuJhKdr4B+//XxQXEK2joqwFIEg6t
gxw2j39+wXGWSwIGmfh13RWqrYPT3+vYQ3OzTqtO2IKPt+C4tFISqqUzQUVQek77
kSXzB4rcPf3B7fUrKTciItcFCXsFBiFgv5zSYilByIKJwRCTtUUYv4kyUWqTCUpX
s7BkXnaU3I1jokLlNl2N/q8nc3eOn/IJQUWlHJrgZ7lxj8T+HjO0ohx2d7IrD2ux
LK75J8WTXea+6X3YbY0l1mr7RrCdfH48s/5hLWzaqaW9lTMpaRI2W/61fUkEUbpv
n6Sy6P+cOCRSWOJ8e8mh+/3cjEWuSekPPrYvxcVTVTG31ZG3mxtlyZZkkKargFta
bJb63wIfPPFA6Iit/KIGzcqRWhap6XKExx9N2Y+2QoVi4Y6P5kHocJMOAJ0BNokp
gfpIzgHjf3f38xSOQOYeHzxUaZPvaCIfelOl/z2waHObr7kj+/qqYouN2nAEEzcJ
rLLmZVJgG3P3EKmuHx4T8LvUbuqTZ7/IYk1pbT5xsgu0fKjUjl35rjh3np5Oqcgr
zloNTspHdDQUEJtPZVLMm5dTbvdOzpzVSfbHHuoAr3T8sUizWwaIco95XLiZyHAN
RBkwYxPJzdJP75F6U/d2jh/t/4ganj5fM1NVzLVYn+AlWInJTVuEteVvyZnKGA9f
QMtq04LR/y1L4HmPYt963voLsNOvPmUt69lFdTo+l6Kdl6vopoQI/q4V5vcBUux9
9ptJqLXuxTzZ5wuPpkbVKvz7KnsvnLpXYDKp1OXiE1N2TFOYOdQdPeSwBJlWE5w2
tRv27UHhWJdEmnvuTcUrs7MWoETbe6OzR9RKVwByGDyuZaWSUW350W1yi7kTW1zJ
AZBVY4DTjVP+RcWc4gcXCq/LkzNNRRlT2GSGTuPFE6BAQrYZ/7B96amEDHgNUKEw
hWVOpCn4/0e1Sc2Pc5qtk15ZBVd34l5ePrVYrSGOpP7GduRFq6ABVRJIiZyvzyA6
JjP7S+MO/H+xu3jELB95YOJ229ppF5Y/koSPFVuenWc65JrPB1uM0hQvG31PpQd3
yD0bQWr21/s0PW8cWGc4vilffCjk51vK4DQ6zKtRqrn3aKi7I7eYm5hq8GbUJSVD
iMz1Ayx/XHn8RjM5EzztWkRB11tN2NzQl1t9fmFwWWr/DgrVbbylnzpRguTACBGe
5/W9bqFxwIAFRcUWGXaT9zorjxlAhVmv3aIkk+h8ED55T2rOoQTocvT5wWI3Ix5Q
XciRVyCEAXu40BSpwGDsC9M0l/lVSOmMcNxBjxrNOdXD3TlNbKfjAsVDCiz69fgk
P0qQsLLfJysxfxhPaDpvgrgIAMRN1owdL60rwIkaO/cho2rRFN/n7CX7nPTdWs99
iOVwew4u1Kao0AITvIDJq9TCCtRdnuiRBMyptyq9yttDL3oyJntTOuV/96gFd0mx
TwC1ewW9oa/seEQQXzV5VJZrakp48NgiqYmnZhEk53N40b5bhRCmVU4tsJCSnahR
28BRJEBD3S7Qi4tIhnOka+OrCjTnnYmvTvLD+4ZDZPY1O70u+UrmSlYdX8b/NO0h
izNBUYlbyUcRv8VIAO48kaOPpnm2QgeTkBciJEJy8iCVrWepR9oXyYf8nXHDKGTr
CVf+3qLB2Zs8r70zgUpdkbDD01x0NhSglLlIDrmZyT27HUKf3l0aeCz5Qs8cRd94
xA6mwi9CzTJlPxP9Z5J3QKLCfzZ5bIkuHV8uNHoD4IMiL1fbGdEwInp/TLwwEMhX
AGqz9pb3CDfdawtcZmux9m5Dt5i2nczvDvtNpFVelTFq0c+0EJifECrNeTRZop4c
vkCiEGOKvkylOGg7MA+1hsjciA26Jcn1zkpmVL9qZoaFwAKdWvYD5GaIksbrE9G/
QYgwPlxTAWokj2D31V502kotOy5/Wiinpt36/ya57vsUmJFTfa6Ttv3C+tLb9ALV
+8EWylx5EbW661T30VnrefK4zXiyHTXXw5giTCeh/Y5stl7WVg37agUDjfW6dZce
LT/cpSQpslzMMhWtzNPF21xLtLQx+WZahOei6H39135wLg8QDXyjnSWWPmmeIAzM
KlT49+SXkx/vaMC/oLKkVJSK+dHe75KtRPJ+4KaRth6/pOPfJRpgqYsYCVAHmHBb
08LfxQo+PHRUFk5eUaxRt6mbsiUapfTRhZU2ooK7NDOPUMPZ4dmj2exTdWv4RqSF
uipuYgTWXyd+gHBlYmWe1Qk5t6IdXoqUIcLtUzAm3S+sjVAzoJFAOS742kVhfTmx
adrNBUa3UGFxibuFYiNRG+MH6APJ/g+Tn622kVhIt5j/xYiG316XnTarA0K5wW3+
4sJO1VNA0VtHRF1oh7uZiGWaTEPBFTPSG5edosBAfgAsLeTRl0L/PhoNqIuHVBkY
EvFnq1lRwBAAxN1inGbQ65hlTYzbu0MmR7LZyl1qKJIw9tzhAATLgJDulLqeRZck
aC9/McoTMRUdf6FPZUbCV/JBo7UEQweTfCn168AVnzUEc7/gV4u0zYytffADRdcy
+uV4rMnzYnhdUSaK6x9Q8IC1Y8oRq9UGlM13SLqkKROn4XrxzsDnqHq+xeSGiGaV
OkjG0uX/VHpopgnTVbcjmPwROmLu/TXdSOyJa5unnZWMvXwKj4iohxNOjOOxXCE5
N16nuB+c/hiqJW2uQ0ea6j9BzXEXomdLPMTi1SoJEkFAIOn4BWugx2knAsQCOCy+
9gRnhBUTg9fG8UmWLc+Qo/tX2f7uCQwfw2okSDAc3qdf813xdGbW7BDMKHHQxuco
r/Sswgas37PQjUaHrsUxh0bd5SNVQQ8xVFQpe5JpSfYAGj/B6l6ZGW2PssObKJRN
Lnhk0be+OkqTSApwCmTMEtB+PRmklBW2KpC5fIDavO5wXQkG7zKsArjYUSboU1jy
rhwj0xYd3GkD7z4SXPIZQcRuSqxZ3a5E4ylZVkxCvCPcvsLKx4I79LgFTk6GWHTR
PL14qr9DJwg/2+dXmi9rZSC6J7lJSlZbN2tPGhCSAja+WZnNq9jsRJ6asDv5NJrD
oHbq/IhFPJLV8dEKIOdoTawLw3l4LH51pLYisXugzKShErLAGW5KWe3h9gB3byqo
tcLpfVTC90hehViMQrve+X7S1KuCtcP1Phvccdepj/BuxSUlK1jZ7giVUdMlmjCk
tsiyKMSmeAeSugEy9BsP3bT0/9BEVmbDNIIIXSXdRXlSRn8J1MuA3qx3zP2tPi/O
eTfwFbltkn2xrHY9l6uSYNyts7rY4f40itaTbw3CNshOTGYTMZhYCg9pEt+ma8pJ
aV0MN2odT1HijWefyBfwFG7v1I8XGpYIbSIykhHPVTMJRbgXnM3rdtsP/gF/wptF
oDGRbNJWMiBKSbCbaXftvIgaN7YBS10Ov+Ws64JTEVSn5gSEfrcrl6J93DpHcfYO
LjEVq/ifP3noZLtFGNE1SFAwtH9ZWRmFghgqJYVYms/NghoqdAqYguYsy5B6PYfg
BBdnm08t/21qVPzxtLGivXP118cOkWDa/FJO+J6Op0yHU0jNFXRZGV2Xcox3Q92s
TvsncXEXPTyNN5KJY7Pz6tbGUvAY5NtFcSkqcQX4FIDg4VUGX2lynoJUCLBIJ/Ih
b3LwZj88R+DvPwc+sqfP6dwase0rSZQQHhBlzGoy7MIrWTyv6vV1tT9RcJKaLT5H
5C7+KYP9OCuRQv4HIym6dtdIohzRK0XtaUGMhJc2zTMxlAbN7aWlIdrwsV+JoFWu
RB89oPCrP63D2bsO82GHSlhLbpSxu7b8NRjKSJbp7yrA+xJteTzeUAxlLFIXf3Kd
i+kZe0XnCBOZ27/dwrbutCzzJ++6csIaQvXcBNDewPcKUSxhJa5TZQSbBJRhggoP
iTHHv+UCgBsRPNu70hCpHsIewCS6jN4wKvaYVifEqiZCd4xPpovt4oBkrPzImZgA
/QgcS0zKacSnPlIFw5v5fmKXtMFwdkYQZTsfEMiO+cZ3rzpYZIPdbu/DUeM+ngAk
NweXeH2Bsl+76c3BYNO2OZhimrN+B06vrjAEY661mPAWURvWUJc1oH0eUj4eCyZR
ukMG5R/81MgZznmQOCfMj/7+wgJSHNtzDDgDOGX+UmQXRqnOu+gnABJ/gdjs8xWg
XDanTE6/grGS1XMLE6XnC3UTyXIic8gPWeAioYZNJusK0/yzKT26WgjskvUorsWL
WHHM4Duig3xGt3xgutMnNmijCmqFp6e8eEu1a48Tme8VdKWI0ySGdzp19DJYoR/I
px3gVGLS4oOIbCTfwI9UbTZ+FEHUHHH/eNI6e3ltV0Og+rWXvKxLLmU4meWUVhy0
aqRNWfChybpowlla//yH704THG2mH3AFtoUqHv1QDYC6xOA5/Xui7oyoOFaiGhKO
lKi2/oXK0ML/kWYhXEU5sqJ7jXNOW2sDi54hvCpx+3qRL7r60BsY0+fsZ9c0Gzbx
ZjCEUp/4hgZ9xpsEVXh+CsJQ75IAV9x8aLCcM/TxPr69Gr/iB8oTG1+lSIBCZw4f
DlPO3R4NH4/X/7144dNQZhKiDPNsUOs2K3SrMx1Ju10oxvPfMTcrLQsb33gr5yWo
wrU3RpeFQwKOWCbyCu6nOQHuX3Lh5h/i5dBoPLE+0/D7/eDmxbFSfSX7F1hMb1Id
qJy4jChaGbWoBnGCAq20ttOQ4TxFg303el55DNyoW5QBHLuF/HeOTUXsjo+C8VdO
qFns0K9+qZ4TOofdHn3arlxT2C5w5AZIeWh4Q9Ju+LiHhxTatFkjvFZZWNcJbEYd
i2l2GRAAYcNM+70PjDTITNOaVxXgo0077ekofAzDXAp0qegcJq6pS8ANs9Rb2XPb
OWh+L8lO2jZKuDqEkz/YFhXvPePWlZ1ZCTzYFqMbQhbtZlV9Xyao4JD0GYk8pecE
OQxPlT81n3gsznJDRWqVSGvdCfDpzGEg5fwT5hMKax0xVwBK+cGukQAhiA2SuUmu
geltL9OEztlIU5TUXZWWZltYEvL10Dm+2ZzTFAMAfYh+pHXbMrruOwXfOEEsClBS
fu8BEWiGft67cGOqyRiswk2RrhKBSNhX8BavDVwmJhXKzE7+8NoycxsNKJmSK/Ca
wkc9WfTX14WzpaBOg71x230z1e5xFy8szIdPYW7S9FQP9kx8sjy9ZYPsiQMSY71/
NldE8G9R6P7cLO1/lwAI1zRfVRrIIQ2/eve2U0DM1yivJcegpyBvM2pTqwoZK8lK
RQOj0gXz4ImzP5OYI71sfyoWr5+0e/XMI/A/RS9bmd7L3oggnAyqzItui88Idht3
+x/OWb/81nE8aFBUxNVsQIIGAXKWT33Qx6MBYgaj8gBGpIPSIy+a25Nvh+T5bBcK
3kCUCHUNkCRYGycnwHfNFK/oS5coPgZyO0pfImm3bxLNpvDEqvlq/w7DEj0kMJt2
pyNtTrT+qmZZdMFHHSScNB2iQHL5uTvXVCHkExnOzC+QD2fdW7u+OIZfsv2TE7PL
ZX+Msp63l2rSSslsXmVVS05AVn6kchVMYnKxzgcsh9i6CVYW7idW9C5Vv3VxCJyN
7v/dpwzpuQkl5+ajEmY1jgw9DU6VhqqCvpzMaXnEnvM0/G2G/vzI7KYV/bG//sKw
OcUMxe2u06AjGs+EBkh6JQ++rgbudUjuc9Wrcvxd4CObU3Ew0StGBbRaafuiQuaC
d1+wmrEoYesSwHDOJWxSpzV16IMObo44Gp5atyLcJH/9DYsFvIXYHe+W7zP7vEpz
0pzuciKbLq1zQ2Pg2yHH+IO0Eu89vMbUXqerHCGKsaEfCG2gSooS+qrUQ4rAsM/D
Dyv2zT6btbzGoadXa/DxVFFreBkWiiicwZqriO8wLq3xS5D6Wb0O8ZgiXpYLdMd4
/09GDCFNI/mHdSgegqnVnwb1Z1crPv0lgKhM1YKXqWIYNZeNRIi6NfE6Gh6HkXVQ
2Ld1mB0Wb5Cv+Gg4i8MkmU75OqkQIrF19v/JDnRpPnSaFfMvzKFP7SSYkqLS+2gt
lxlSc+3ZjAfZ/mqolsmf95gRzIdwV6iO1wAiY+h0RhMUoWowyN8MTuTjojY089m+
iaVTrjiIjW3/zRroOyBiw78CRPaex8F//CP/DLZjc3i26RzGFZE6A+o0q+Dg6OKt
PKgQbkvMPNY5JEz3/KJuYBpqhc6vUUvL6ayfYXh9l0oleL36Sbh+ZEmubi+N806r
8KVNBT3N0Y8/+VOCuL8MtUA9vlgN120d0vb6gTB4fpgFDea9dR5/4ueLQhk93BM5
l5BrKLrKk07RdyDHaX9SjVo2/jBT9eVXQw58L9iaBawGUZhS8cR7bRmzGxVgC7GH
cdPPbEITeWUOnUZOUxxmavbfNPmkn7uaesSZM/30hBvnA60iaV2AL11UHG5J9FNi
xbi/7X26L1lnhYTqauy7ypoOuZV6J4rEEEh1vt8kakzWi9OV+C6hO53rAkqEjCg7
KmRZK2fBuvj5sWvqCk9YzxxfqKUjt/+pSCfr0xqIl9QKYoh48PdZYRCjeuV2rF9M
f4YQt7im2/Bxk62YQ0CH7NmaSFsft3d/fcDRVlMi6PAui8OepdQ9Mx8n32Wai1M/
ZZ4h9c+S9Yln/brjI0heLSkJncpC+HnXzg94ZAD0mXf5BMjbWYFbJctepAhsss+b
h91FrX3SfsVyEyUl/mfho5SuwyeFIFwje4SCOc3OgNB9SRXeGLzyFPoLiMb+2ocW
o1B58xW6MgbBUJs13jZeXtWHxz3Itqw4/AQzBtFQ+HLzK5JnyINpc+AlRzn6yVBK
9yznhgiEsAlx66128Xnj58j2rVht2NRtIRI78JMXNAk/fezXrWbh4Wo/26qMFXyH
EYbPcKef+aVI06SG1o5O8hzjA20ot3+XMReoYAhv/R9hzKfLFwKKkW24nkrWtGK4
pMsXn5Oc9VoDjCoFMitXFDS9JELFs4koul2bwQzRDggTyoH/i8R3yU7/w5r7652q
REUQcXYJBspRjw8oOvw1p4cJ3Twizmlfdc0o72uufP9nA4mveNcaiZ4wh4K/yHZV
xw4undFLMY5TZ8xO3uRDrFILg/02Z+OuXEkAo9kpEx6yEAT8fLdmkzKR3MdPGw56
aBh0pdgZbNzhsxtUyPfNtQcyJVjeF5uuNCgnlWITEefNphEOk3Vnh2okxwCEfeUD
/eOQw+dx/R4nZjSVCOOvFm5vRcYkTtRaO1bpC7S2ZNFEcTbx6VWLOmppvzMhuVT7
JuOwJ9cvLxBkQRX4bNJ8JWc5+ZZGPWfwNTkTH8Wxi6BmhkMs4ek7zBsk7//O7sJT
TKetRinycgX3T8MjXZDB2sY62TeAVq0q2rc9vYjkp+xeBXXQ4n9gU/g/Z3dDLSua
UfVaCI5a59YFs3PFzRWMkTeAqZ6R4ibuUVpQHWUp/P7uhatzUg6yYJWEXeHK+bL5
0+m6uLCg8ugFu41xCFXixSuATY+XsP5gClqC8gJgOzuo7NZMZicn9UZF9eB7Br6h
WVgE5x8MOZkFOxvoG0sSrdzvZ6uqd0dPi5RfiRT28BbQVfZD4qEfcnIluOEBVcI1
4l9xtN90uMvfEbyCbjZ+Lrpj0mntK47NVVuUEvXj+KtdOHMi1sv7LY8ORTktI+dV
gg7bb8SoRt0+QKrQnko+rIiodYnrJkL1H9L5rqctEWLknMGvCTLVS8qKzRmZuH/I
RdLWutK0YWpAezLApNjoSMpaVbkn4CHjZMtYQ1aHZCnqN30kEBh0Ct+THOOswODD
6Q6cWcYMkmsLvRwcVx2MXmIUnh2McMm35Ch/n5qLFE7pBGzQvoatwHX/hkYRKk+P
S7zsZzXiiqCtVn14SuFANcUMsfBrClNfnrtqzwSV+UaoadsZwkC5CIEgfHgcOAZk
GdC7754t1DId/F6lYxrzHd+X3JMSaIJCZ6Ex9I6dyu/q6YwPbjqMpeAn6v+0zyfw
bVFTWML6Atusi4ECZw3vuI9m9h8hUG4hxtJMwaEka0PL7dYduUjD7tT752IzEZUu
7TQKoZSB/TlyRlOQiCOVaXBZh/ukFb8H7og/VAVSp+EtDXBbBP43LZo9Be/jM/hq
Yv3J7SWHUFKuuetbbsPjVYMjzVnOtzDGh2KrGr0aflbC4sCXXaFPfZ4TTWrZLUlR
QFAnV0UExtWvsjCX3O9py2Q0Ud+O4bynPin97rqbdTEzAU6t4XwB+YqkXrU6ORgl
W1P49VN93tW75lbJCw6SH0lADfqQe4diAeVO2Tal1iqJDO1MG7N4FkXb9AHGkLCY
Hb15CSJmhoBlSVOKsnbHJ7UwlciaGYvDXw1ufxjvkzKV7vRYIoDe4F/IvwotguHg
iWd8Bch5hmr7YDM4l2UoCrZ2iYBSo0jCBi2vItwmATo4EUnOfNtv6qJU3BfgOMNc
k/nZtKetf/wy7usryPGbXTaWmvOhsx2Et+BC2ThMZNb3rvOhBUoT28XckpYA6mQ7
ZN287PBx2Y9G/npYC5O8wIllIrgYEo8FP2/it81YhaGBj3hH+oT1XdpeFDrfZ1B9
oZl5gIOZOgriQM1WLzceYZg2oF1gbtHQqqRAsOSddvPQcL7KOJWNEgCqVphUYzL5
87tgObprmXdvjvvqjUeB1xMitjOuKspqt7GLEjk0c7GfU3aOrHlo3sJZ23W0OwrR
XVpWE0iuhcyorihrtTPDzxKWJpj9RfC4bB8BWxnbjQU81ceVWNDcl8Qq20UH2HBr
gXzgJLGzMGE7HKxNI4n8iZ22eWEsbhG6QOJEg+br6bFEiHzp4EKvDHYiHsZRseQ7
lE0Ql3MY7MeP6f7PKRey+0RxyI4xEy/gV893GM61z4HI7/LaLsC5BvUrxZqcfAXx
YV4bLdfVlRLDQRBQKLSFwuQluiN65CeUwG04JZlul6hwIyLhzXGhhVezEOlWVWbt
RgMlGL7LHv3h9tXu3/Mzbab9/a3SzeN+k1u66yXrgwnHJJRUwtQAbt1aBuyUh1pA
/Hov4oTnEydY3hJJLzpeUfxkcIEp8j59b76WUw5LKGevwe1rymUjJy/N/Mg3mgRO
gwaDInvicg+aKLZTHGu3CN5VZ/cvyNW/2jtJiOkPjbREWoOar4+hZvkR7a8IHOgP
KhZNJ5BQ+LsmtAZVwQFEG81SNSIv+AOrwOiWt+zK3ip/AIdg5L06JdswklQmWuEO
YspSgVBoWnOiPghvjIQp8wsTlF8uaJnlR9cyIHjqvMk0/R2kOjNm9Hlc9YRPAy5f
WQ5NIvH5CZrA97EDBw1SiZFnoXYNZyil7GCZ+gaukxv15E5uuCz9BRxeg8cQcarA
RdKgTu6VLwQ4T5iAdLly8b/aW34leU8Y3Ep+ChuVwqpDU0Y/fkjJCznp+xIO4bbE
OWmHkI5SEp3L90EDrH/UqXLExuAd2cfTO2e1cll9Pl4hvf3Kk7B4fwLVaumwUQsl
OmRHfqiPV3ZdSjvEJm6bd22tCXnrElud6DJRQK/ayWw89wxxliXt5BRiwWbvXV8c
426I7Q3APaMC6s35CfSt+81IGvT3kwkT/H9pNUgnVb6b17Zr5rQfuBI1jV9jKCuf
vCgrxURHoFkwmgd1IZHn1r2ezKAD/++fS5O+yVwg1ttjfd4Sr2pjB4lFA8mFZv61
T59hUOggcwehAqOexx/Yl+FbSt6yU+yYGdGt3OiF9zfdvZApyJfSuA4nZ2R95Zns
aMLChM7960llRPGNFDqmDKEem4FVNk1q3DrBRZ0BwDnpunTn/6XAEuE2r8KGQX+8
S8UtTYeKLFjVSQjOvpdn9w6R8xWVz+cbMb6lDS7Pd1rBdR/GxFAB7wCzQfJYCCW8
+T+9JrQT57lL2pToUqQphZcXEbQukxs6Xw8ZICb9a2yavVEurzMIBOw6UpJWFAuR
nk0UoE5d+tfZwN661ejXCy0lWcr/PRbaZNkaKGMh3m9J7zOnPfqo5mu6sAtzvT3e
MMZPSOzDdZRKGzEK4Af3dxqxP7KHk78gc6eX6HGCFe+sLKmTcp2I8g+D0ycWtr/g
MvjaasC1kGQEKQEnnYZtqMWsrR+ORtGrKYbXSFQDpy0OYDEs4a9o0BkXb0j4gliJ
523S8s2sVGQCPZNMi3k04kQFxZrcG2eVcPFyWjIccyql4d6uCUSnJIRU8GtVvWQ4
fOSL+34o7MLu+3KUH9K0eXwFdNnLhvpQ0McROPK4WXaa5baTQ5ATNTK0PMD3+WLd
LIN6p1wM0eTbGkIYPq9rY0kPjIDSpfOuMbCJujEwo3XwhJ5pcv3DcoR6KPgUM+RK
zSmeuUZaIolUR+jUYmlKR1zRPRsWaNYXLaZAWAILxZhmdQEw9azTpxtPMzlFq7sQ
mx+GIYY9yvbCoaFLs+pmXylyYsXQH7W9Ac2sBN+thLelAhwwMk+tmiRpYK3LJRq8
adqQ9c0z0QaRsj1M46EpzqJ9IB43Iw3SBTc0jO8PkThmNDfeeJ3AEhRJDnfCClS7
Y+HSDctwgh/iwu9z8KaWm3P+ntTwkZ/Z1gMhHjfNF73SvJs+lmFAIEwSMFDHAsM8
/I2tq5YZmEgUd++oe2NZ/HYitLVWMe6AR2urKqsizMKPEYSG0+SUAitGtj6OA1M4
OtM76yTmJwMe1eiMxrVuTIdNcIGfulMkiid+/HrkTsoUvC0kELLE8jK3vzYtaUou
cWoXmqRwWIa1XMb+oVtOu2UNF9tQiHeD/0v6jQC9mMXdMQj+zYgLarmyeC0tfk0l
Sm+nU6srjB5HFh8BcoO11+4uYIS7iRM8DSsOAjulMvaFh1HKgmYaHXHpXyIPB5Nc
os99yad091TByI6D9TMfivjStyCNUGpnj1d6CQFQUAqA9r2URDAFguwiyXU82uPw
jMNszj+A6t3Y0VY265iU+aEKss4G0I2NDQYLNclxIA8+KTgJJ2ckRXFD9HbS1mpb
y8VtYuzkR386SKT9pDPTjGLlr0s67OYcdvTGcQ7VOi+Tcaz5iRits4Yc8v07NApY
K7ZSKlh8hXROknXnrKUA29jYHUm2xWIJbsZuqcKcIQXYIVNEqIB3oJd9lJi8poB2
OqjA/srVRTeS5rKc3o+FN8CFGbe7zwCChSzyQSgLxGYbtSCXaEVuXo3Jsm3cdcjl
CV9NBb/OOVpC8PMO5MLjtPAlPLNpjlhbQNTbu2IE4LuoBf7gF/ImveNau0QykdhI
00I+7272unSFP36/G3ilJmKZJjHtPxhDFxXuc1hf5S5A2HNp8ppZmn/0lH0s9FEq
QqnBewl4by1Vs13eesEZ9eGS+9RMY83HlzryNSm8+pvwXHAV4S2OJ8xT6xFHXo6L
GnVxC2mho+37jSuLmqGj2HVVG/rpZrENk9itogQGI9l5N7nbtD2mvu5ivmdWs1C4
t+SRBy075Vca4ldNo3nplImi/ZiJp9DIuasIa+CUwzw8nTvQQYp0xopI5z0NxsnZ
twPq1TiUtdBnlsyJnnTQlQbOHIsMeFDTbsfQ/9K68qIoH4j3Pg8/42PcX+y1KVt+
0P2ZaextnXZxhHsYs2syCn9dg6Iyaq6zh1NzQSX6APdCQKfSf+SGNAXz2CbAYVoz
kiXFQMOeqDspcXogeKy+9tgVamtyjy0UzIeVWRstQ9b30zHboyJVvTvnoSgoGdlt
wqqCQd16/DfvXcFmGltqQUFvCrY9sUi7yglvic450bOzWU6Xw0vGFwO+6nN7Gldl
QU9XXOuzlTWdB14TBpGSDMiCLfwk8tNDz9a7X9gNcnyHXVLDwp1skyOfP8RtY91m
Ds5t7iK+YP0uabl+2gIZZSGXkGkKegYQ9Ot0diqPBJTHiUfAYx43iZwdODGyKUC1
pv9hBcpfTHNwztGSCG1MIGUA2hrErWqro3fPXxTrYSBscbxUHpBatOh/3f1yYeBm
T0BFhlc9vq7O5v6YFyAghKJP4D5Qa8Dj4MrPBCwBimQeeeNNIJU2dpO40u/SDQLv
Tytt4chXveBgzvH3Y2OOBjb/ylN14tPSy0ZEwhyytHqJ3WwlNHe8qM4DooEpaCI4
1ijGDhEoA+4Ciqk0u8FC7IBW5Vtb8VmhMcz6dqpKmNW+ZpyKamzwbAUKCdVbZCne
YfTC0suKS0DJZVo1O1OPwZPyWiXCHcrrh0/B+kBeQJT9g9OBAfc6SvI9SHVcD6TI
E5eL1a93JoAizHG6Xj5XuIqDQM/EFHJ60KtBCXS5+cy756Mapd8KexwQva1w7Lbw
Rx1fi/HSAMmzE9ITwOJruaWwywl2o6rTREpH8vziDMR7I5k12UuVHPkdNsGPx35z
gSRd7C+GljRqiMa64QGi3uH0Vyf0VheP6tEZ5NyvZRsBPyc8cEli374uCsuVfD3m
4gtECqQSIP7OLuqwBK4K8YJ7O+DP+JHasNPDDkUlLZ+C61ZvZwBVd8CdUylPiofb
XGo0yqZoh7qbvdmHgXR9uPne4yCbOHJbKTKjrVYxXCtQ40ZTRsFFs/tWclVwm/32
pKvt4Hcf+SbZsjNl5tZmy7rw+LAo8VP+Zj+PBkXRa5/yizoiTCW5HtLfNnqYoHJu
RwYyDeRUYVoaGjDid/f0fHDbip9Iv/orijwjeZmuV2dSNFl3rCR/EFlf2eIgpYaY
6Okww4W7MjW5KBEVVT9nMNAIHwNRZPviiCape6l0FB0jeT7RKte4HwudN82KG1im
SIByejaHRW0jMu3y5ZWnWRBBqitT5wQ0AO3zV6vt29XTbNFZmkhf2DQk5V2/MVs7
lRBRr0Rjbez8EigXZORe1znlsJz3dRRyVkRDW3hf7LKPFXs2PPPAyvygq+n7f9bq
O6kkttMCon8gV4/YljG7JJmJVY0/I/ZI5sE+7OfhaFET7tDrQTgVxYVk2p2Bpfun
teXlePe1HIfMAiINezRPvsfU9KgXDAO6FaVwy6wPCDIBuW7tuoGXoBYRAWaZw8Pu
P2efHAO2sFU7IkxHoWp2cVyOjwk3/x4oAlY17y3xeG0qotG5nFF1mYrswvtxyQMQ
l/DpkXWM7jsznlzV3qYfGs0YcRmoE/NaYm7/RWm4m9OuaD3SSZ5/I8HUP9CEtY/O
L1079cH6+EdMa6GVs+crP7n2HTp51dxtfPnVjv5xNtkkFq1Z1DfaGUeuH1ppf03T
dp90Wq8eSUnjp73vl5F4BD5dMHgtgXLqkss/DrXyPyua0iFnO/4wla5jqdoKbz+z
LFrR16oL4UQG4ZPn28pq3t57dgTotL359GtOSlW2jCo27clStoo/0cMYyHkzydUo
Je4nzz+o2iIl6Ug8kboWCywPySI17+YnsTV2fKuDmEMXROv0VLBfwh3GD6m0Orxo
X/Kpst8AOZhDOiwcbrcgsNueouHcw7w5ZUmvDJ1y3loFYGoP2HLSVe0iaZ+x+dBs
bnQsPFF1DTTrYzkE6kN6H1sb2lOK5/upA/aeUwtK0QF2EVvBdPTXpp6PFIFUgxiZ
M9CW2wN6bwe8vYIitY6WDM61oQi9R6u2OGwqzBf0dNo4C3i5F4vWTQX66Fy39TI6
n0bjmjXP8leLKB+JtHAzEF8BHsWfO+0FBnxtDPvwEbP6+K59lSdbe0dXDx/bshss
lZnWBNhtIz3N3fM4ffGXwUbPyWNhADbPpRAwEIVcoBlhWQPuHUJmYXgHBEgo3u5v
OuMhawpo+3LbrdB1ByP0QGysW1MpMST/nzbxxgiDQlQOxDmqX7I+XJtnwLTc6pCU
T/Vd5D4vQZjZ2/t8X4woT8kCQjmlwpYnvsGnFo8UBi9atA4ERbECQr5PvGQi/MPm
CyWNS77k1JNpTZuRGBaCmSwva2kmpjRAgRMRxZjag1r3ySha+aCvS4G2MoRrXyGT
Zt/Qcd+ZMSdGuUr/c0QQBUY+X1ub46MNtTRFtbjJig+3kzw22LUoYZRRuZcRFGGz
T7vK+L8j8hBW+iwzf54Lad/HMhaZ8A+r5J1gQ9eR964nZUhlki5rhKX7Q+doYoyx
mJXsYqLBI9oMITimEi7COR7zomE/GpHB5ISabOU6RSRUiYNQTVlOitjwlZNe4VG/
p+vsE2+ybAXakzXUcmgdTOgOUKelLDXUKYixGx9VRyG86qtqUvkz3er0tgSa10+o
iInDaKFs/UL3LWn/qXHqpL6nZNyJD+zR0bU3v38/HZ/M7G3W5mH0vzmUJ1QWOtX5
OspEpS51hp61L6tdKeqrdamvV1W31zsyzJpm8ICP9d+gTJa/UrmJCMwhnZ3s0ECD
0EojMiSU6wx7U6JEKlO0XFSP3ov9sA48ngR0LXi8j+Y1WQcsaKCei8JogiTYmn2I
xtGaWbxeKselY3vV+uMflabePEsqvfmdBfGLWexWjvRO/Md5bcuOqKX+Wa8ENpJX
TOPxSRvYhPhoW34Z2CnaBzHulq/+bgQHmMwqJ1EnAdQG7SkGgKmojhzlU3EI5U2m
DnwSszwSZCqKHi7uaU8I5oxR15nGW/me822nrZoT9YeOIcEfyoG1vI8LZhMzVmlN
dlskmeTH6tNyANxPw225CGXlVqDTA9HD0d4Kk739Mh40NInnpGNJbDLgwC0UdhAq
tVDRMtyRxoLF8dOgo43PiWGlFvlVoUPX1SzSIvtNdzk5RVfEcH9QRZl4i7jsOysZ
4igcog7A7SdwzWtuoGZmCv140Df6H8CTN75CgbSsYTl6lI6wqRmTmU842KQcM5UL
bQtk8kU5pxV+rgxYnVPKwtmTBzHYZ2rPRy0Hxu+mFQnAKwled7JTmyUZZpRL12jI
vxApMxYJxtZsG7gd2AyvmH+jNgPfxyUS63eSrCPF8vh9NZN9oP426TmtwaJzJO8U
JDkagQio3nKeUfcbzW9TNdY0SsQPiINKqOZK/enJWZB4gZ+hJF1AIkquBv/YdXm1
IAdMhk/UAnKwhLQHbXD9wSufiV5cg17/DGC3MBThT/1nWmbPlkDMF0VU1Wer8XX/
8jhIhkVPQhfHaZehvQIiNA51gWWjMD1eEz4aprG2Rzmq/0qLRiPGqPnWXQx3IpnT
KYu7QXOf43knWfBTPFd7eGSN0puGp6bMwnJDycpwxORD9Pq3koMEbEa9dOf/z1ix
ir6bD2/vxuysFWVfJPxRsiP5Gg8KMRZlJF5CSjvFldlaS+fMB/6QnUpkKPTghVra
Q7XChK6yAl1EMfRxpM+l37CWnvjIzga9hQ37yR3lnqd/ISQaKE9cMMJsy5YwAb4z
0Ad8Gskex2UhjWF4044Ha2bbSeZDumYcA4ZhMKUuwF+1DNG0zL8rAARuKop9vukm
fu+sU3vXJtrQ+YMuDt2/SclXHRVOAGJFo5GNOUAAXgmM6i69X2OdraUp58/O+exp
M7b3HnyBWkXz3m8hWWDxo3xoH9BoCg2/g5w5C/XY4KEaNYuczeqP10q0sHq3dVFQ
ZFgGQmCDdxGFmc5kDP1fB8leCBYQ7JVxgB5lWe4hkNX6Ze4Yo/QcxdZId1/zHzZT
X1mylBYmRSFO3JrstVo++2wqliYVe9CjJRGPmUUSOIG2qnaEnG0ALCn+b8J0hjwi
dr8sSpQV2GRnkPNrEmVbAH0/l5lcHAA1C4cOpOefI588n3WCE2ST//d4b6CKLovK
IhuKNTB1mMg4wye8vhu4g0PQN1hODCCwY3J8Z67q6IAOs5ZKr/P5a50hW+dxsEDX
Tw6pQWyasVZHC/V0sZYGYiKLCtQ/9ZElhyaJE1PHwhJyBPDB/BoTio6Or+7w8xnW
c34BcEzhFBcP0LSTDPiA22THC33+kQ41+NuregregFKWd2/FL0nkKrp1uEFLFb/q
RB98aFBdrb8VSKzHHFZT5dpEzKDf1zqeIOmpvfjvIVEQz8e0Le7bv85ikFWSmdOE
paOXFOuG5IxQFzXljEcG9dYeLJKffdigk1Z8HSvZy4TEreQaxPSN+Ll3ZLesgG8J
a+WPrWhZzFFsCFjQfTlYLLdX8ynt20ADhnJWYvyltqVOHqtrzarJqbgZnzkrZbYh
+Xnj/zK3A+m2rnuPMnlvArgdCy31qGw6l0a7uEqBY7T1NAz7hrwtY/7RlsJFCmYa
Uqe6W0CPTg3Vd5y9icPHzMFbNQYWnu1BjnlgDd928uQnJs0UoR+4/YBZpO2aZtVL
IgdsTpguy7Re/oQd+8HyvOwjxGW1v5doAA4jemS/wx++hf+8NJ1Lc8QECT1FkoLr
KwyE2DVkUAEaWP/dflyJrYFvdTn8INTQ3kxP8WHGPaK0ahOIaIOb9qiupCJXbGSo
0zx5HdwdiJwbcEHL/ODJP9G899OAb99XZgQVAZlt3/UJYcZPXxRnOBRSFNiaLrhr
OvcxlOjlg1tYSuTg+eyECssYAD0RCtAfz8p+5/QnBtBnokkhhxE1tsHk4kzMkPmy
OPcwgUpCT5SIrxG9W2fl7TfLYQIRjmhTEydVrEPi8xUDEy0R0W0PN0gSusifx9r1
eln8UJig0aLYcwymQcZKgVLq9xIEBQZN7m0w9OVfnTCEQ275J3GIIcvm8c3B3ywK
EVfSEplH3qqngFj/coOWWwix8AvHtRHBH7N1KFgR2DddRzgPEWF4SVBhsV04qQ6X
yd3NjaA8ACtxEnfn5CPHChvQ1RCgejzLA0TeEqGXLXpo0PGfkv3qVXgdefhTBoWX
kCtkSJqUtPQ6gSXaEFjS7/1F8+5FvzMgUCAK6quX4igBS5k/V4ytr65tRjlMyIs0
+J8UwZrZscTuA6RJvWZzdETpDZLqOfE35kX3Iak+wxsBt7MCxi6bs1VVvdbYyw05
0Go2NN7ix0R04FQKSbYa7kcnGdOoNJFPyUwGR+h4MV87Oe42amXgAaUQ+/3z6qhW
JR15SbFkzT6P9n1AmUi0FsAbK2B+FdPfLxmnUq2j8SiyH5v7w4i007rARK7AieQJ
LjLOU8u5TGpK6bLo64iWmI5GErW+8WgbbkLTGU3cTJXr59pci7KZALtwDHnA6oUo
V2gsghwife0rE0D4/d2emRw8MOMQRRSuS/DSWqHqjA+b6OCGUu21I5hNfX9mBjlQ
kHgIcP871j8/UcdCPPX6SQED+EFW7lQDd8S0MsSgStKo91Le+aVRjKNs/MtJNlKY
JwQ/sgH/5+g3RgjNWa/VZJjrX0cP8Ew/DbQqYQPyyE6Si4F6YkU/+pTAVanzz2to
eqfQlyBT+5OwfhGsm3BhDbmyEqPGxV9/tLqZN4yefepOY9YiTIyf8R92UzjXZeLb
C8IyF1syRfuNGtpoZtergiltfDybMH13ymwTZyaPUFYS1ZFMiK2qfvhooVnerstX
+E2QW7jc3vtTW93xwZbFUhv2HczwLOJY8WrliFuNgGii8Wky1CaH5gpLRseN01ew
acLy5bONULBgMR6Bxwm5wFcSv5CMwgrzucfEsisi/XPbN0A+MDVR7F+fNC/W+fVj
7Pdp4zh54N3LFHsDr45hDrsM3cOLqIg5+Hy731pblVq79xvWwn+LVi7uBzI5SHdK
rPlOOp8Bt2ze5yrO6W04Jk/XgluD9itiT/CBvlABRlJpc9KRh9lEaFCpdEcpVFZd
5ZztBAzoUqLVHcNmrLL84JrrMZXfu0cvVTbmRhCMnaR2tQyv1r7fRaub1boq2za9
IgccsaWp3GcyIsEUSWuu1Pl803EbwEJeN+3uBB3bQDJpRVYQD3JgZg4Y0rJamhWr
C4As6lkIh7WBBZFbAtyEkhGny7juC32eUgJgdsa10hz7Ln0aAmRX82gqN3H1a4Ng
YWQjEpwRHKwmFCOSkGB9Rg+8yLSScXJfAkz8zuC8FCrejR7HjXjYYuwsYCWCo+Oj
qKwj3vyB4FPcViAHqfgV9ngUaIB75JluUe8VpyWx2ITOmwczg2Mv8RaoMsUUTZ1g
AMPgRvQ+Ueehh8298uvOGmsZHeAjwdSYSijm+U2M6SvAqkrIv5UtufSuWU4lYjp0
soa0iUIkaiwPnA4deLmcQDvBjX83+oP1zS5Q7pWA2kjbL23Kt/6HsMs9/w+rBQHq
sN6lRAwFHY2gL5UHW3bSkxMkHcUYm28Cqd6NnZJeqVBnRWZ6macuaqh+J992Uk0y
gqkwTXb2sA1c29UW2Mdp6DSY9hqVJf9Y1c+UItlY7XFn/eQ5iDGDtJQAt12yAqv2
zI28DPqh5bxyZdThysh9Q/Rq13x+uVv+LessIJP2Od2An6V5y8JcZJt+xcIHAbeN
U2tBnMsncmFtPtanOfju27bzWZTeD94E0fsZiy6873SkB76ZU0xzvaiudxCqHYZT
NNK1h8P3yU05cIcn6D9Fd0GawO31I3HJdNrJQa7gLK1ga3YqPG9ty5YO68cnGJXd
X1Xq6w//48s6Dqhz/2EXlJ8XDgYl7OQxbhhnW6bz5YJ97/FSXhb+UTjREU7UtpE4
VWL5lpwipAi8O1WhTe6Py1jEYGnnKhl98yHhI0AMKhF/zrFSXopr7bXArKY3iXEX
NwpfOjBn1K9alKvzQWbxOAKLsmUQmZK/UYapSedxiQEPACemUWwy8XArr+OYFbY3
s5HWG6hCA0ucpMc3EDYnXK8RXy4JTeSR8yuQz95PWvAbkDXnszYRetviN7fvpIdd
Dfj/0d/Xa59DnNw+fWnCYDrIeNlirFEJLcY6e/tByKBL6w03NP0jViuP9e3oebk7
FjU24HaYvsx/BC4c408EhcW6R0q2tsZ1cWGV+CB6rVenbIDgyF4EEH2koxhbwFOI
H1wP1jU0k6ZrvtiJwM8gzOufF0/xgT1FlH24DT17wfIJnpTsLPRZA4WCJlWIfHma
T8lTCKCjB9+YatG1aqNtwrS5UeDgTaJTioBNFbxuwPqmeS+Zw+vzrqYZ8zVZ4v5u
1mP/3wKsvQbNQGv+gQZySdcpNYfY0zxpkRo+tcGuhGg3UnHxJZdautJDT5YB+xH4
FOGelptCAqFNyJoCUiN/jXuUhW+vvgrxZH6iTNbKxZqHDduazAree9Em98BdJisV
eyEDyAB83yqKCeqSBIiXi+ey1KloKYFGTdR9pi6vLipDBh+bm3X7vAhsHO4ggeuB
6c5CKwwXYC2cduX/vinHBKFyMNTOy3Zyta3d1py022GTWtpyqLHEG6CzNOU6rRmz
a5UqAyzBj9KPdtWaX5cHXg7gTW+uwUTMovB5bHc2e+uTBK7B2u5P8ngW+caOHkiY
PBgKsQR7HQ+3yqUMVFkfDo5LIiRHpjkWyQjqMPFFMbIxw+9HNkTv5lhIbZq6kHbX
HI0QcobVzUvsrHshyS3ICXQdHTztf3FlGQ37+CcbFAXAth3zITxc313eZ7LXnRR5
JAc1CCdQ7H+flRlmnAGVgAVO86jKSSXs52oSlWR6YTFYeQ6aiObW38w3LwGpQbIP
TjeTo/QSoS8MgWsAfYrrLtxJgP1aeuwEObezK2ldMdM1KIoSi1s2r42Lx41fxMkS
ul61GJv62A1RF9YqLmVCE5ZIx8XgnzO+/8Ak3wFXgV7lItkE6Nm32YcOKFuER0Jv
ZQLY2hhcTM65MBNpbnU/RU1tF1uWC5tOgil5KlfvcFKAgXDrn+MudBLjkaScXlKJ
kSg/XKtF9HuxACTrs0KH+CKQ7c1UEQc3T/90xTExqKbOXlR9M/Lu4AWA7Z1sPPiU
3S5WJ38gKgugVF8zeQm3EXWwXrdhvvtBDeBGydZM9kSO7UwUekmTJ/MKkmFhlm89
P+N2XqHUS6z41M2HV7+X85+rnO2S9iGhhgmQRc6MBspFFCQqujUjroqY0c3JxlnS
ErX8MsLPIKpl7BgckGJzAfCCDBBCQXaVDgNsS4LcAkA/fb/pJRxjd+mfhedzXslT
sjoWfAdmwyo+yRsko+j9epnj15Sp+y/nAZ8h5MWpCAYvDZmu/hWNwv+HPxQgcAOY
HgIvqBxxGW40cvbUC05aneRjW7lPJzVfDsqyQJ3c2T8T3XNfnQt8fNvWdiMcLmO9
tv5dz3KlPEjhNL+Xied6lA6FyJVerNcaTuJyduk1LPYhPJ0Q+cPH4VuDmVRicW3/
iyelGnW+H0eIdadLQhEsPzKwLnrCXyBM4NGSMDPeLDXk8TCeS4/ZOdRX78/k5C4B
EKqSvu+NyYQHtNB5qK6P0UnmgAdeh+dt7pgJkGTsUaDawQgd1FGteDr45Iig7w9R
ugPwxlisQlW9ZzdzihC5RHDhRovnj7erHFf8ewTXmh5Ue8JSTg2tywjU7hx6xYjf
pQ2h8jtQP2HbiCW8RV7Ql6T/cJtOshTOYVx88Iu2b5VPrNzunpCCO9QtUlmlG3YA
jTrEg+G8i2hHRrqVDg3rYptNVNn7nqOJ1Wk7lhsSGq+mp+N+GuqC7q5/67UBJ1IJ
856OJEJiu9xjOH8FaWrJoz0/y5Z8I6BWke6Gqs+JPTPrQ7imbIXKtepgxhZdAUu2
1zm+cVUCK724sJW9zYMxUNhAMxhUqR2gb7yRKAsPoj38/8fDAPmdzYJEIt9NLIu6
BarP15pZlZGElIUqU5wWuUDHlpGQ2gV6Jp9sZbjbmIG6cdb1/3BAPSdxjhHA1os3
cORA4jn5g5fL7cBZaIH8SQV2deR01fymCRn9pDipf8K0z43B4Scj+IcZpg64p8q6
1v+yY2nCnLN7xBJ4/Wj/xMoXiRO7VpD4bjDiaFWkkLSskWRpTgUp38gRbxmm+Wit
RoQHpQO4Vpffjoqz9tMYPMe4US5d8hU5LixwJ603pc16YZZNdSAFgUXlIJ4YwdOa
CUjLgf3JRcpfpkGyY7DgOYRGjft+WGBrHh+yMI7vtG6Imz3b+0trnKTgTcxN/SZs
5JKYFF+uAoHjJlaond26hE9uv9lMQu/+Cb7LIGTTXd7bAzq2dHG3mlIzB+O9dfDo
NxbCbPMEQgmQYmuKCCeP/tW84TbW8BgZN0S+488+Bqjw1MaN+7JLbDoF4L7KuSP8
iF46/+7rU1wGPACN/D03fBDLdFu7UXlNUVkPQt6xKUHqPoWcEF5YGvXBIQDSbafU
h8YwCVeb/aYgXX2BMp6fdY7AntACwdFZLc64jKAFQn8BTiydUrdML2AgIp4QjWgZ
RzMj4TZ8xcvDuQgUKjsj5zYuoUSDm1PDgSCQskKqXEfIPBv0+mewQsQiJf01thjH
nejhjEvNauZ9N0FFL6WNR+PjGFg40nL5YbEg2jSX6vE9QD+07J4HFn+0oPUwzq6V
0iZNPyqs79ABJdOvmUM/QkVqObYlDTo8l1tklFDlobyKSnlprLHBHKYrE0yftSbR
EkUgDLrMq7xWpuh/mQCVutgq6xIfcQxepg9AX/Sgmx+gR6b07/TJqpa5a8ThUYXz
Ku0rf/dH7uXL4Rwr8UPqep0cy7wr/8kyCnZkzUFthCgeOXhyMeU6vDxc1ypnpe+w
eceOcTxPFTefMcFiaPlm9m2J9ETYpr5pLxQQ3cX2gTFkxksudGOYWXgSWbfYr+38
BJb+OqkEriwgG+h/lOUkgiaLlqLKPMGgtLrEfZnRni1FIMfbUcNX0D2UX5vi3/ih
ZiA30uan8MhuWKKZggzQgI/EEXJzKwumrqgA/LKYBAtq7qUnpvGujp1Ve2kGpxnA
VNeSf+3BH1/2pQ7LVl2uxJCjnTtNW6+9eAc5PKxuAcxfP8a2Wn6L97crOE88u2xl
RzFlMZzFeCeg0MhNioGspOkSuf1FS9EGn6rtO8cRni0s6wIIi9iYpE13x1+1PMgJ
QZyMB3JHwZ4NhP0EkxH/HEIeuIOot16VkRb3VucTfOsjpFehZY4vJzPnrBlI9lPh
1QhXfg/wU1XBnX3qYvLGCB8do7NORKFTLxPBxfMrbeOR3jcxM1q+3Z9dQMAUFEsO
r2UoBBFVJxgtbthyKIhRaZEQ1dN1cDNDgmd13a7LQj9gYdRgnEtpIkkWf1ePei8a
dZ/FLCjYWHzUbUOvS47buAuD+W1zbGfnuoMNjPWfbJn2Ke8LREK81k2qv5ni8lF9
NS1RSJTGNPU4sappSPYU9t1z8858uF/xV79GhZZH6Q95m6ZUag2ast/G0g6GHPYg
Ab9NOQsUSTdC2MX7BThMtEvuNbLb4LP8Ajx2viXtGxeecbmvlhb1zKHGXcQjthoP
Znl4QcZSg2pFkDdyWrG0ni9e5jM1F0kKvqf5RfeirL+VGuINY7wASQc1f5VpuQmz
D8WoOFU8eQCpnA+D3NP0j26pNNAiHPMf4jll2cnOBfaNeClkWclssZHl+02EEgfS
YCMTSqPxOhtaWxbdMQUp2c4Q+mLhy5Z4oT6PWPNYwZ4JtgWmQ42qwQAzB/6bcG0A
gWSmB9FCHVCV2Qg5o9n1ti0xy9f+QxK3gQgfessscTZmASaEAN6/wJRQ7ohHgtKJ
MyB3Sb8BTvml6MTe+0G5XJ+zecZVX1zOw57cGOmRBeqz30Yq/sSyMwEr8lY3mDfB
uezitbgsxZ+u+bwAv+e+aYpQ2mUzbsG+yeApprM/JH89mfYxUWuqYBuPUjex7kZv
GHfKJG3YaK628qCiFVtcrtAMxAhdyELvpNPwZPzyeYzis0kQqcAemkgauy7+AHzP
tpSrfo5JCjC8zOZURpucpPco/FKfEAkfsbMnkHfQ4gzfwOj8xlcCnG5lAtk1lfgO
dZApPvpcumZyAUSYjqjwllX64dXgd6QYgzP5ufdfUCi9VXAAiWpez8PApUGfE7o9
qS9vHrjMuzx0gqDR+65APXykB5GwOHZ9Pir01ghAAMrlkdjZhGZS6mHh4/rKXQf+
H7K317TNz7qcpUWZgIjLvyxiZaWqSpGzbD32XeXqiMO7lJdJdaJ5H4LwKnIYFb6u
IPAtmUZzQHLaqRAwuKBBmQPrKdAjA+G3XlQ3czg3sjkUYrOAbgMiViapyDNNnKGx
wWEjHwuQ/nDhEYAOS3aLlfrENKgAN8ObRhdpnt6MmCXNgonAPCPCFymbT315yt22
3q32f0KOrhr4OeX+KoIwD68MSYu8eAPIuYn5Rz2PmYx5y9wpyCw7tciHI4bwMjva
B631xpGSQ7HMCsBuwuFEjYDTmgw8v6rsZyMcfgGGwbN7qcN2jXGlK067aqLpDJpR
G7A/l5B9nU2PtA2i//9FwMyk0Xen4BAuNDo2BBOmbPx1XoKf8d2XdMpL6rN68pBu
/T60kskbGqK12Nl46bOLczmS07CsPc//XeijkOX/AHgN+sOdK5rYnO7BiWPeghUB
4aHqopn+ETsUjBmTdCCXq44Ilk+0eOw8bp+WRqZePI0/GzLfkRsWZxzQzxYhlfjN
FJRQQoi5w7ISL4be1PIlwlQNiLmF+oEsqdYyrkUpDNCNpGRmszVYRy44Fof58eOh
0M8Jb2TZQuA4HQNhKpnUFJYTgz3hOHwHP1+gh8AI3uPCfvcCZYxscjlFtZ0JKnrd
ZI464DeoGnZYKI+HIlLX2UhMoPrhd/p9O5MNPrPnH8c3icNOZ20f7o+b7K+SMprv
zB2KBOoqyD0zApPhUxRP6JAMHs6BVW+ka9x+WHbN1H6XVqrAf0SIx32/JeyQN7JG
pr5NQduNWS0dcedTO4GHd6lZfi9svmtM5XU4KuMwBjiMpKSrjh4R2m1LsjdNxO2C
yBad3en+2fUcSzeR57hAcdp2br9hKToPiUDfk65cn2hTnv5A+umKauhlXG8iqZPx
AetXpIrjY9NmxrXyJS5i4DvwhxCGP3L5Y4CVVrYj+SsCUdOoAGxy0NHprQO94IdO
jo7zKkgUMfDmXVztCt69ehjy07EW83a/2ofvzaC/YRjpiiH/rUJcv0iBEwQo1Pkg
CWyetsfTkgHybNC8pDBl7rov+RxQEh38oJV3ussNCnBXTobZxsTfWhkMjtsVTE0A
r8hz+4LwQqs7O3BLPNIi9Qoo6xcNItHWVxdBszvdOHOWF0Virwe3V1tY3hahyqmR
ODpSSN1lg/vVue1AqontsjdP/3kApF+hOQSqGj4GybL7LaCPystmAs4XajCAGlNo
Opc4du4xmI3QZVkR2fUeBJIbnZ9FwYp1ZgRzqBBdoHF4mi0kTFiEoNWutW/jIsgm
W35fNIjgTFiIy88TatyQvcb2mnNCV2HwjNXWLMyvGK3CeCw0YP3yOC8RZFvCMxlW
0ptMrVz3BRvQ8Mtg/XXXbtOwCa7o9/RlCwTIEMWVw9L6emJbvsVmPJxjLuu007Ee
5q28/4he1EDelswCnBDsBMcWpq9F3boWEJ0t42Ysk21X67k0C29lg5dcyMiQXM9C
PxF3jx/VlFbqmwZIR17lzx71rOU4GhAiPkQjNHshb6KJ9uOWD63VpqsxY/hyrpfI
1qXeG2Ti0STtexUsIjan57//TI8y7kgToZPiSG5m3ikkZ1NRIuEjMEch3RDlSKbZ
gqYl3LX2+eDr4OamYNQDHi4ozRQ+3Wu4IEaEUwMZ3GZ/LIjPX6adkYP4I/OqfXFQ
YohJvKTTrBr8QhY6ozQrxt9aKHbxJ21wy0JKOYeauEOJHzBmtzZQ7yOl/0TcJJAR
6y0byMDOza/WfneYUCfT98PQllOaqDSlLzTunvCV/I3jJfWWrZJwzJaqAoOPQPPi
7ZsR86ezSnYoNO3u7lFdEL7NFeHAWES1rD2Bq8ps6NwCwJxWjKF+mC/aqewoCVSA
PwC1tEa7LHvgeX0hK+OEXpZPIuFMW+At/oM2PeNqEJL7DjDsBpo0c6P+Y16zxYLR
KQLiDsmbAB4NsHhwG27GectpLNgSDvpwVlrCLJwpQk3Yc4xFTpYCORkwkTYVmbdj
Ht1OBmerTaWKmDRBicRahT2eM1X3fGskBzEXTd2MrJOTZsh60SJzjDIfdAX9SqJ9
IV0+MdeujfkN3HJBsKTCLNSY4hEMNYk98Zl7SyPPpMJk7tlklLANEXN9leq9xAOg
UZd65QLsCYQW9H1wAZeD/9BI8AKvgfAy7i+2NlARQD0i2AQSPxSyzEYN4ve2Zh06
4IpfGhMG7lS126GTaZXRrajFwwqDxvLMqcR1A7saCnfsDdA6MgzkF0bzVQSse3O7
PlHYvjxIHMGqJn7X4vLI0CEHlfz68MNpBSF1DPz5uGn4yTqdX1uXcLQp/6G24Otm
dd093fKSJcA6Wy4DeZ2To/ZIS1IGLTVIdLvxSdLQiWbvtrpsrs8D+qBfz2Pr/w0c
tl3mAqWO6QF+0WwSst0OTO1abPbfE5FW50sJndsN3+4XytlATulIIPFHv8sFP4yO
Ai3NWRJmu/yeNldzUuDcMX4HrhhGwOwdJPVp35ac+q5vHZ9VukZUFXQijNMQE20n
geiFHBRzkLoOpI5E6vim8BUUQiGD7TAk8oFN1ZJHsjcFwNdqaATESbTYp3vOSSTh
zd/XR6dBp0+D342OeZXQvQpdcqWK6QzRI7tirFWZggAcjCCHH5HXSax/XdjwjVYP
Fny55jOmtb2zyTE8g0eabGKvtZ8y6sYGZ6o0EscNTyutrv2ckuJ8qewfhkethe+/
g19SVbbYFnm0xxDJmbSXdQzGmtpqxXP65HxvfRixR9otsUmK7EscJLdMk3E4tXkv
sKxtN1MoSFMuopVH4DjD92H74ES5yu2ZdsD14MYPnrPRJ2VvC4f8PbiRVgstS+VB
LI3GZnWmZnz2dSvAWNmi1G8KFgN39FGr1HnencfId9fqOeX21mxPFM6zdG5HODUc
kmwtx1Pdb9eCXsUBsZWypE5PqBPvzb/Pu+M8n6/6r1evD1UQJgHxMe8JHhEPdUWE
M/qIfwo6/adGwukBEL4WjqIH0qEi+sKy2KkTYEWvJA10cc0JIAI7BZ7XRnEP6YRr
59+jGMeHrakkeyA7XLUXLiwfPctA2n4oxjUPVOPoXgaStJ4m0gRvwM1WVwQFkvwu
NUKZRz+NPHCz2bZOTylLTsSejjf9evZ/a5rYsAKxzjQJLcwoKqPHZzW3S/2BV/aA
tp2ia1BtJUUzMIjMn2WlXvDP+mRTDZzV4uJGlwfG/9pXTRogqLxWFKjmohKWttrF
UpNbybohUop4G/559AVnq+aVnPNeBppsESnGdX7ocyDHIfQvJMulfm+1Y9GJT9xz
Qray89Ijx5MjUFgNkspAoeXqPqMLmgTFRkyJfal+PQxO03XkBMKkSZvAxyojFFBu
KioUBaw3cPTaLewzuDW79mNEI3B9A12xK8BWFzVopOqiyVQHYBIJrHwFY0RmNEQR
i22I765OCgr9/jX5RTGuOlaDhOBd0s+FScwuqUdC+mokyUHme2i6sp6y8jrDiSSc
9VnC+eb/v4dDCX/NPot5RPxQXCn57wg14xJEEqE4uxP19e0mqQzlHMAU/vpmpC4W
c/lT5wqZ05XzEdW9QLijeG211wLZVhRBGYmv3ysksBqyGKtVyYIe1P8Pgk46LazY
mc05dI96Y0PHV2Sy3VylHCNuswtpvIP0laeWN6MViV8aAxACpnWWQ3TCd1+16T0I
W8svrWhTggj4AFWuWu77d3d40hPX7kEPfk2a6kzxfTFyAVYg3jrivw0gHn2OCc92
xAk6Fb8BcB0vkNAJaNtJdqp2Kz69mHmwIJ7wIakHUFYVmFPUmvO6qn8gsiVUwAfG
iTufYzWouCHXwP3vVMaUrzovyN8tG25RRbAz8pN0P0DWpaBk9AK/TdU8tJq33X1k
OYLL/W6FFBAB7fASH3Wfy2C0ZeTat23lvMVklqrqZdDDfgVlb6Q/ccHhy2OSAYv8
nzWn5gNDFTGyh+akrMbQvYqvqV+8YGcGQPAhJC24FSA072X/nJAuncI8zrZ8pE34
BHx5fMVnWNTzOPNPst6iRBym7YUCxkn52qZkIFALsgGcmCvRxTPSSIuHwI2wWKSs
43PNBErqSti5xNFT3t1STED47IpI7dubONEIOY2HsgwHeEaTxzTQY4usR2NxjAdL
MjRs15nd5q72dpIfTNRbTAgy3OkY6a79g2ERM46N1PiGE2/MuKNrb5bWEQ6uu1I0
xkpQV6XxCKYW2BSfJj7JTUXL9CxcrdbcKrtdFbGC33MnXGulnig56HfP/HsXOeqy
K69ExVIZCITviNeXwCbO7bgPc8XRIUg0jsInhN15T4m4iJq1suKfYnx1T9qFUYuK
5qWwZa3Tl44GlaYFrykeAVyT1pfsrO2vQVqbHb/rVqmIkKhU6Q0MiHOl5sHIzyVp
iFbDdxSxnjl74Pl8MyIWhTVwOAxG4NdaaZ9rQVtzq4DquwGCv70/rVeRqwmUdNuR
si/e05RloETeSxnzBZpDs0HqUVVENH7wRl2lUPoq4g0L9+k//WQK4Ss/KMS5M45b
uhenMNevDtcXF0bSvrXMoZqRLHkoEed8KHVzDYt7ViAlY9MSPbo7YDkIqAoVIuHc
SkYY8y1xWqXJLHNauLkUJLGbHVhBul05bwiaPeHA33HOCQFOhPjlXX5uwznszoMl
mAZJ9L40/JLYNYn6Hcvm98FYgpzyRko2rU3olLiksnEzfhazZblyMOMRSr3XqO6V
P0j/pL96I5c5rw2WxRg1XuGpqOQqBhLfX4gaV5flo+2ZTjIWPy5QwmMHm6oCca7Q
V1RHw+9jVxssc7jcc5Gv3HUjdrAyCIz2jkGEQycFkRrHApNWam9WG3++AomxJiE0
to+4M3u1au5bwG5sNAUZrU8ibt0CBryY8NPVMhsh+jzLvB45pjWHP5+PUs0YYdo+
vqQKUzmQs4+oJ1exzgXXDJ6OPFlGuUJLs1nn9HMWGaofoZUiSK1zK8UGH4alz3r/
KVVkaT3pSuugaa3sQovlLPkULILuyZP8Sw+g6FGm2Pl7B0IDY5bcLKycHVScQ7Bv
ZM3hxPUr75KCpdcGct6w7kT/Tt8dSWKpqJobmiTicnl5winuQVEaCkHGvVh7Ofzr
uA6A8Hff1nUf56mkrrho5Yj6K/3njxy4SCDlIDgCFz8gse/Ekx+5wqnH2ib4DcVw
q1Yzt5HL1ROUylLp4toVc4NPO+5uvkHHP0Im6Az/pHr1RSS89StB2XtNPfTuAX8C
Ijl+lpmW+UsMlgkXoaRWE6pbLpX4PJKYxOjG2Vr6GBMnS0eS1CqyiIAbjY4HTQBx
dEU0PZ27FKnS+wRCszh2RRDxPZL8Few3PSMWlcjhYeaba1SCvp/D1X/sN/sdLPVA
0ws/Gg2FuC5P6C/MaBYh0QA88JDDci9V9PcOPpg9DTc1ifaPyTpYjEVXtR/hbjHy
Kat4wBQAsU/0MFOgRgswQnzpnFmgLMr8m5UzDfXGqZmZdu+MeqZibLyRzw4X5eOe
wzaeyap34UytNYHRpJB3UdufWwT95cZ4bMOkBYwquEgofrRE8cUOwC/QyxDLeE5H
2XwTljg2HsLpkqATDm6reUDXBtO/WjnjQMOgaVmcGboQF16xvMlE3ReLsTKoFVt0
lB3zIHdB5sMtezCmYUP19jVrYseJ2/l5KvWPuGSHyz368jOJstu66Vp0HCJMRAZM
/BaCb7xGtoYZw4m5QqlSUMkUl/yXytnRtyiNJSTXgkq7VYvERVgss4IFiEMMmAdZ
6OLFId1MLU1lGO4Zpc0/4XUvt9h7S4IELE/LvNAgUze0gTBfMikP0DSjH3sDm4QG
wjViFLFmPyRJ6YXP+1nPmpCiHxVHebjDOOzx5onINy8zYyHYeGyZSRTqqxnhvWhK
pNmQ5iqW0woBSH/zkDulRFdYdDhU+HKUeqmMc4JY/4sVfalVquAPZfU9mM08fta9
96SxReEC++PVnNA1EnW1+iCoi9AAbHl8JcaEEUHGENtEo1VjGD/8fUVene9u0P/8
B1Aw0AXxi8D9DaTX4lkGWWHpmL2z+u0uiElLPcVN0F0toDfK5TP1R9+mOZT8Ar1n
o6xudt1R8MqOkmbnSRTTAuLx7UtdIGZ8UA/+YF61YBocmusBUFqXQJnTJ2RHDWMP
RsQ6FVNRFB8/i1FgTWwH88Jy+JhSTi3Xx2Efu0YHNp8hm0yJS3lyNAyAP5578ycS
AxeX1QPzzQIBOtVJEIZZ8dHbH0LrA5vhj1oWGkH8Pd4wjB0D9GAKT6XEbkKutigf
c/Ql1w7fF1kkYWK73Bop4bIGfrSssuDLhGQveSuJAus8qItqFM7tkAEQJdO7YIB4
YuSCg9WXex2CGmaLkKZZNJ2S3NbjX8oXX9coSMuy+2U5acjiV6QOVAwa1WSR2CBM
1D6wVYSVD1/K/UjYcN6B36eatAVGxs44LZMt7kOMdaKCLtTMUfzkockkOgdXHWfW
cKa1mDzTh057bnQcKZKv453bkwIR35Rbx+hl0USsO7wwl8e4CwPC9NBv0Y/z+rHZ
MVvfU5ZZ29RFzpSxWBTydastIqbwxIvv/3h6pYQN1TKwvb1iU2NybsMHe3zZ1BDj
hLZSg9NfyS6bb/0W9VRs87HBCYgOAY/q0IgMFYMYJKMUU0WB72WFFahQFe4zISY3
51nvl/giYtrjuUs/mFUaspcHc9BqOgawOqIZVvadi0KRZkwdP5bKepbcNhbB0IAW
n3iRzgTSAtMgg+4ySjp0ekNs8SSH2rikWLIqxG0MQ9aoNVcUINcLmIB/4B2UJsVg
Hal42FPqH1NPEa572MsrF51JFyDXmCHjB3FlE8CUAixXkP5946zG6iOJZPbf+rUA
ArvBUGwFzV6dNoMlOp+5DBfn/fo41JkhfkMss0CYyPYjjj/KQByWwQ/ZAKT0NhtF
18cAKh9XuSCGBO3mEKqpvwGMTUbSyihbCmgRTBXgCBAg7HbZbdPk5AGnKVo40IHr
WnFnD6eJ5iRXCJdp/dauDj4y3ONl7E0JQFRZ30Boy3BHU+sbpQlNTEG/lxCXfa+j
kmURCSd2QYFrjatGKp0TcFlkfU+rzebbGce8Md+Xr4uc6Hw1egKkFk29wbnJAXEV
1V0AJ5UO6ddulBQmECCNIhWkHkMmeHOPYFq0p4k342H/jbhtDRht862Q+4yzLhf5
G+deOtFFQdBAagN5CdNq3LWQ3wH+6ARqGPWs7Kja0AigvcX8nxGlu27Sritk9h1v
VF3M6D66+Ezjm76K6gpGMn9LCMYCPWOnmSNDfLiSo5HxhhgsB6yCd74H09Eendtr
/IBYgW/aVFliupopP9zK+W9tG5YpewxOqFNKTbV8sLaacyF239D070vO6/55kDVH
ZjuDvdiasrBlgnxkQ5NVSrR6zgjKqzf4HvCRcU/0yPtmkMRx4wJAVI5Ydy+0WTg9
OO7+41O+luvfqGZE2vye/KpQnLBodPylPQPCTuEouaTFOzPvBXPg0etMpcv4Sj1+
N58dgolaYthieU2LmvBDSO1ESfoCeADH+Im2A30GcxS+gwDF8guWVXRGxy6W8EaB
oQjKpIMeVgWSWmJwVKvC+x9cufAXV2L7YjQiW8ZI5AOabW6KZSZOI3SLg7/pFpSl
Ap9Sb2LuV2kM4OGt8HEDqyyxkEvGXHnvJXizXDaIOUDAXzKDGPUTo1BN6QWRy7sB
OuWOOzv7d/FdAmfxj1lemL2FckcY+XAUia9Rlnfi6TMaMazJFXGue2TtxHbOig3+
ud5dPfc96L0zIQsvZx6yQ3QWuSFKqdJirmm9ZAcKsNrQLmifsHEurN7OthqjM5GY
ckjiTLw0XFt9/lUUL5bAhvIax8/MakIB3hI9lAIqxrMXcnQN5w3PcREv6l5/1mT2
/0nChSoWyzcVoRhfPzdaLvSIhAsRNh/P7+28QMPcfzTM6mruB85/QjMVOWkhgTFR
qXCHJeV2tdIYZ5tkb6unzNctGI+kgu1qUXzmT3tKb6SNRASjxd7evkugmGRraRc2
Op/lMBLLc3O1hzr8XdDEkmTsUuJ2zkGx/MgRmHFAxY5UJW6b1Iw5xnJW3uOxgMIM
q9NtrjL9Nf+mIBZmjKTLX38nCaHJg7dY5U2c4MsCqtraBaVdquXrtXU9o/fD+wHj
kB0t/fQYyYE3SLfVpuWSb3afNIEdH9uh9h33u6M9mOiVxGvrLVayaPm7a9SY82ZQ
uqb1z9UTNKDEqoyyP41pdhFXHDpTB6dYIuoUc8sfLPp/wqmzOnilNiDoV16lFL3A
kQbkggoWWaj6yE/pOh3fvMm5VQ2GNz9EpQpdl7Vn0/CgJsURIonJ82PbdMwd1j1I
LC8xEvWkFcg4lXAIrvrqBdoOUOjEFaDocBN7r8zAOhBgcboUNXhuTGl3gGn8fA6f
fxsKtQlqPUqK4qyxSznNNyujbuYtmXxpN44dHIP4P2dnbbCJpYRozshqeH3G4Dew
RUKRhlM+L0dPZ7INuFKkOSsl+htuLInpv5OP74VsfHo+cgXwRnXjWb9Q4vp/NH3T
TW4OYaNzNRdSz0Cg4oguTrbk6ZAFq63PUNmbSwlmuGLuEMcwx4vO/rvUP2EkMJs0
cRPZZTFasIFFLBcELEoYdYIeqmbqBgxQvAi8Lk2GKPLEnQ49/jhY7tEgLvLRyA+P
n59p/m0lj/mUyMkI5oCbaYVUS8o1WepSSMrMP2IyrhjUncvtdphWGVovkMQf11P3
eDk+NomsARB+k5R15WxnyUQ9+CZW92piKVs2LLUIKQVDkum+9QaeUOm/hathSaDd
4UHzLNGgxRpDLvDw/d3vQAHnC5/RMZNmWApPsA1Ya7FK292C8wRUbjhYA8Tshwk+
14MpfRghihTXAU4Z4EKJGRKsgazLMVnYXz5MpivLrBrAjE10gLuo42IwUxY9h10I
JYqlJFeTjmbJJrx2ig8vjxvU5eXxpv8tX8V4O5XlfNuJxfwxvDZ0DdY+6FogFMYm
ojaXAxq5Fjl98V2KYvJBo4i0Whe21itHWkxzfxTBdJve+vO3yWs6GjE8yp3XZJGF
wonRIWyRAKXymM8pwcEeQ5oYYWcDxZW/Mz22F3RbWWb+67QofvFDCcE/wjtU2Bz0
VlHADjkuPldJKrEAdFUck3CsZX1AvzV7Rplyp97SkTL4/hKqerglKgRvHfnbv7Yq
BZ8+BcgRsskhWTafZPMfv5FmynfWeonySrpQbEIg/x2lsQkASuzGkjTeAPa8KE81
ej5e9KT2DpkdGzKCg6hbYe37TXk7FNQbyrCno8QyyTNGgJ2w3+fexdK18lBRPDgs
f5qOzaTvqRH1mpCEqqycof8kFnAv21s3xc+lTQsE8uTmbiDPFAKwphuKlKkDarap
pxWKJAVu0mgz0OZgD6TQxvsru7pCNvM80llsrw5MNhPIY458lEAmVjYDnLUTb+aw
i9T29wMhF8h89TmzraK+Ry6amfVOtUwbzvjDePS141scA0VFm64hLuADaVifPJWH
BHwOt9ydoNwoxTh2sQnEFs1WfEPeuAQIFgdSSXRKM4d44vaTpEYMf5tpscZ5kTMN
4wTJy4pYWBwwy3eh9h1djd0afIbv6J8UM/lY5OCTJCk8MBnAdDhIHqVv7PzHS0aH
daZTs7wK+RBgYg/J0SkWi/0izgIT+pVnz9itZcdnbJV6MrgykBBLEAD8u+kvtkKi
VgnB63lhNpt0TDK+zR/RiZp69oaM3LgKpob0ZuEp/a/KyscvpgByUNP/gj0DDDP2
HHdtacAmeKkcnutMM38zZdrvc8aTAN5PPv2KG6BXwfmp2WL48O0NRn/BHCbzvgVd
Q3AO8vHWvGY4WXBq9drh8NPvoecPbths77lxN/NLaUcsV/NYl8j3WfjdRSRDCXoE
RZxX8QgGTw1UrMauFsrwlh7AeQ+0bDBy+reu0joWn3cbzq5wPm+AOmVkopRvYggo
oWGggCF5vRlNlEGnHqXZW/LtNTp9dwM7ouEM3k1WMQLDsRNbRlqJuPMIDpszmOHD
Om+VP4NHTCbM2JDe+izhoKwUZ17W8OZddZZUx2QnoVzu0182Q86pevAy+W9/Io4W
hZ4MGMNxT8J7ESsNCYBgIX50VvABB+jbBfdBnq4ZAokk/GOW43RobiOdvjZ+w4Dz
RtM+x6v168ntmai2hC4VQ1pXlUoiQ0q76kvzT9efj6ZtXqvHSipnMG0jsBukWWmG
mxRdfE35LvJrMD8HuXKiVCDdI0o+vOyaIcv8yA6SXDUU7PBHkm/oTgn65lTYM+Gu
rYKwE3l9/v/fQ3ExBfFPpLNF8uz3pbcJHdy8DU02Dsxt3kYS+C6K1xUiL8yU+ROF
8+1+kGIYY9gbuoFij3eLmBonbPN6YA4fEFGve0Y9xpoa/YrGqyVO2ZD2xmVTxDun
0uI9BnwBDRhFrKGM86s8n1GPH89K3W7yGJMAei8du7tJ+WXLkhU0pukVmNEN62km
xlpxBKD903SR/gi6TgMqpmOxANbLOA9MnFyiorjz+SWkZSLfuQmdXizd4kcUi6Ub
WlWFl1I4oCQBlVQlp0dNtoJRxz+I6K0Uql2Xy9Zk5KL4cf9hLxBl2mVtPtoItcBl
XGCv2Qn7BmejY97oVivIpRNwBeKDPkerj9OZxt+M7Ab0WZuuzKmJK5hPiCwQvhP5
KhljKrOMplPU0sNRV+r+11KdHaEPbf6IqjxPnbTNLkD6rzrutqnC2luatJRPTuoX
RQraUEV/KK5A2cc74v8UhnF+aqc6XHq6fXLeDs7+4XiNwk2+7R8C1fdEWYWK9T1Y
W81fAVENKDsvYmc1lDTRaobyNcRWPtlQR/oZJzFrW4ST+3fQzH5Q0i2h6sAo1qiG
7bm7IEwe3AZR/BoK6hjXDr5ylcLWDC0w6bAc0SnBqpt1XE9gitGzbuR9uf2so8p0
suWCvrq5O2g/BSNANsD9c3+sU3he56gSKOduXel9HIJOSp5n/VU1I/KZlRIjjTb1
8nF5AS0w6ODL7KcReng+6y7Gv5PDaloS2If0cSkqRcz4NZ6UZdlvwBxRL32NwPqE
tjx4mxZTjnjuqXDTvoHX87TS51eaPQvrYbxotks9SPC23BOSbNz1n2x4ISJlLHjv
MgY4SA6d+WSiqz9gfvH6bXnYNFcZf37CeaktbPqXA/N8Bb34v0GIXuE7ivbrtwdg
YMOlnOYbY6aR27cVsRQ4eD+FAkzZERWHbsb9yIIbiOm+ocPpzh6pkCbXCvFKxHKE
j+iagTu/n8bpGQv2DjH4YWpPOuB3DV5j0jTa0IKjkGN4IMWGDIdtKcdKSCM42+K1
CaA8aqnXmqGw9x4VgcMzqSbuTwZEz7phsFtddwh+XnfrVVZe/D67b0HnIp/zUdPn
Kl7gbaKt2q+wR94vpQGn4IWYH3bfvIRT+vRxgVvusHKBiu+a8VOZrZXdFy2q9H7z
96RpfZAdX34iD6v076M67xJaM7CxxddK7P9UGOkbhIQDgXCQSrGd3hMqu7TQeVE3
a+3T+Lz6QtcSn8m1K0776iG5C5Vrtk38Fde634C2BweTRX+CJfDL99h1iVAcA3uN
ZcuuREZA+ysqaZBv5STal2OqMOGYrO+HH1Ea1tF3D0qv/hRJ8V2C3hiD0ntjFt1f
Ai/AQoCpjBBMYgptqL1hjSDG6rzMXyCxJAhfy4pE8VK8v2vxIAPTIVUX1//9wXPp
we98r36Iw8YH/WhN3tgaVatBAOZFjTWyB0BKrnfFHed3TvjwH3B9lqevbeG5i+dC
IZjAg+yiyPjwvLJ/cOxy9gPD0kIFRGpMxsh9l8t+OCSB/vzA4V5uufDNVd5t8I7s
DAFX+mguYBQHm//mP7hNCApg9qPKUSg+0JVgZPBvyNeOD797GhF8v1kBXOm+fifQ
IUbdKZ0JwiYsHtOZbAjGcQHqcRdzrlZVsSpVfkG0+EJP4bweK8lklUZuhm9QVmlW
noJ1vQipyTKRSOXRRxhVPkh2dJW9RbAsiKUZJ0g1/HbqqV32jxoNIbeT5gyJlb6G
cu8eIKZFAesSs3eA86SSnOLVkgr2UBq1mUN4IAOAyHvEYhuk1hVFTGEyt5H4/UQY
nalK7VsQSjzSnk+DKzBECOtprF5z6PE3NQaFUtZg8DLD4DeTyYlY9YeyctMsZwQu
o33SJ7TSVCqQC83x1CnSb83CxkgcTKToTTAWh31xoCP4BiO3dVmtUstmkvVPOBN8
B5B2l7LQxfZynfo6J4QFdvgNiY0REbEsBHKKEoZ4yCgIqNF2FmCLev5TJWPd1cXc
mdpU08NY9+kq1tI4nY1czbMBUWikF4dtXb7sSFyR5NlhuvTY+1+iib0rLcZc8zTe
wiE2lLYAudvDXiSehiDuJ8hV9r+iiJpnLz9Xd9KOqOrD2zgWgEF4ZG+1xhHT5/K1
/KO2tNQsmucLAAivxxZzvMYU/jH33OXHwaCAhclg3KUgKQ/tmBjSPoj0xqlCA0mG
xzaNOAIkuKEjlrXxhzn+HsI8PPoShKqzAfYFvyCN7zEoeiDwTVv8s++kXIk4nzWt
1hawCd/hWa7Uy/MxWcAwUFP1libUex//aT98jGa0Zwy5GZqALnfJ57A3MTj4dYuL
P9UKEZDGmxV7jwKp3BjcXssETqIIgjLZT7Jf4dImaomDXXqDkM0PpbQahDDJMyW6
e8j/4sfYYYxjG9jaSKDqJqA9SzEIdtSI+LGUfChGGRA+aTE+9Nk7JNTwPc4bA0Ux
XyIQWUTH9KRl5v08wndhYo2RqLMb3p1XYLdhDG8A/xXtrK7IrTpnD5mgqFvuI1yZ
GWaxTuF1Pd+QX5gGUcIXLs+fVUNRD8CSWCW/+8r8/cXRQ9tOy5WJFNNWwePI0gK4
RCxQ6bjUzNMVForwvJkDBJvqzIT/HDufgl5IffANt91Xjg6xKN1UjGdSdVJt8sO1
jU+6MDpHSwTztNwKW8vT8gxhIVUlAtwkEDRu5E3MaKeIvMKtVaiB1hU9DNjIOopZ
ty3veFx2abRuwm5gIod9uPgmVGZ92ERIzADYRgZ0xL1nIS1YNtwpkqod9zEA57xC
4CFIKFF/D293Ege1wtDIIpmvXfHC42b8kojnFAFil2jcrsApBUDlaAEpV2Ps+JmQ
VQYUh/fvr3pAhnnL/9R/DmDJ3CAV+Ei2WlNaONWY4RjQkPyliYKvwXoYZ14XoY6K
qx3WMdWRuXfg0vr5OxUpHDfiguWRnu1BKpgXhtIQ7dGKzPNd2+Io0WP8tPM/j1pl
J9VqxaHP1YaMbiguEocevcDD/d+5XAgIqhZYonbLVmv3yszxAXTaL6wCvnwF2s/1
P0y2lk73IlLA8Ap61gYm+6l2VfDjw6G7r6K5pf8LhuzUdb7V/uD0l016wyXhoG6D
6Y/GZsiH6aZA+ZTMu0A5TNM/vFEeBMH7jYEj5IrvGGgTicqiLHSQZVLsG9cyRK2j
D6bvGR2LZMLInD8/QZyImZIsTwhK43Oi0q7DF5Cdbul3/9Ff4PG5h9Coc/ISXO51
RteCDeB/K6ZOrkoUfhMHcjfYqMP8Gjug8xfmH6DZVE0vn4/ffeenqHtmqykXlaWk
83xB0kPXrC9q8NC5mePbOgd7dzi6LB3dMbWwpb78/FTMc5TR6YU5g4XlI+YwUlkO
20Djm0xB5w7ko9Ser6IkvYBv4Ik8KLJ3enGS0COyW85l+Kgy4kj88e3x17uwJBx/
fw1p1IDKIoE7CsvhNGvkS6tTHu7voWNXiToIe8wKiJ9gBu3VlZUjQp/ZBVZ2TQyr
DmOuaBgFP2ZIjcWWGjSjfd1ip1vOVYSXxLIlkp/ldA4yj6N1BykYTh675P7olgvT
jqJkYpI5HD22HppxHFHEC/dUJ2YFjDStMMPgCKPmTWDIIssEgn+M1gpeeeo53HNc
BSH4ei0p9fT9qzIjrFKJ6V8fZKk0B83MBJ7TtK11DRoqYq/gmiXos9biHJI01Zq+
aTRLQB8yV4glLZHE5PETqcMqdW4kV8KeQJez3SFQnuzzoe876lktaBW95ZAtLJrm
6HskeXZP1Y8h4JCRIZEUAyOKIL01QwyTcvS34ai1vxSxgqmjshj07+aAo54eocQt
c8/Ep6XFOD1fv/DndOgbLVYCpq/IKs8HG3xg5IsRfaZdNwaaL8d3raydYzBlURh6
Ja00usC/fzJNwajgWJR5juyHtKgvaqKdDuUhgraBg4ZpJ+TVXa/Pgv8EbTEzUJbm
OUdEBD5mhSkghI7HXAcsBWOyNX4zVw1rlpUEYYkir+jYJIYhpA7rV5fMElLfmVBo
J0Bm4t8golEWINtuCsxcmW83tpNsoGJhH6OVjM8OTncmJGKGeD/P+3H2ZHuG7L6w
HRCByRXIc6wNhOWJwffadY01LpxC3UfGd+4+WaojmsfvFdjhm89vN6o9FM3Meivj
1D18cyzAwvWVE+8zM49vBz9wBVDLLwX0ugZJt/uHE/rkJMJS4M3UuviyTyMGbaNo
PgcymgTFqiCyXBBrgGdtWt/Auxug1irZLhiQ0Ha9OhDdB9GFFa2isgiPhDOgpKRX
RyRP4P/5nCOzCsPijsIT3b1zLzhMkOMrzl+5enHQPXfoPHEbofKhHG2Ky90cSb28
qYWig3yUkoskK3hiZZZM+1a0/85M4RrABwZSD/GvLBsu8SI22We6WbvzSC+elwOd
OjxuBS9q1o8BlqhwEri2xvO989MfMQvoJbTxVqqdLDpR0hH0giSsLp4xS2j79PdC
8yM36/UFPdlwMzvOhUGrx5ZwkBoH1P7RqOvzUSWooFx7pi1yPAlXkkp/XPiLy2be
3Y4PZ0L8saNnQi/ALGtEB1zagJvQP/fqGmE1oo/WskSNWGIY1x3NOcPelgIfEvZa
RmHpofNtFN3Iro8TwDvFF7zaZy2EWE4QofasFnYbEux0pdngp+6IEakB6CZhtkFF
n8GSUl6wttQGlhr+l19HVE1jj/KTutU8XI624IHumYaOAeohgVUhyCuLlRZHkma1
EukMMCTm2mRk1kkfhyTxWxbUIh/JSdaIYTNBk11tBNfyG05g8ZaIUdfG+m25a/o+
WvZkafkSWXD2IfqEKOMHloC0pDJVnouBZHhSfbkIFDPsS5Vryhzj6U4VCm9/2W9z
PfVRopOQhi9t/C/vzJ/cCvB0hLCbucF45XLz6zxdYnpIORlrx+eAQ5Uarb/n7NVh
N9ZNnVlQGul816ZIQfZ7b0R/R+jpDIu6oa424u0zyd/8b/u4OxwvHlr6/e0o8fa3
BSyneBdqpPKMMGjzKCBruHdMvMypO6yv+2V5uUoHERsmYsQKoghnVetJoV4OD855
Z+hCWcISAumIdyZlxAFfL9O7yi/u1rrUQuevDRkaDcxdft5nkr5t3EnhmGwq9DGm
xb9FEW516fMC1cowa9Jf/Y/wwOHOJR6ezENR8sDC1Z6h8GVTBI83XBasHCZ9rTg8
aY8j67WMK0bFwJvroLF013rJCrnKjd6mUYz+yAc+pJW/a0LZrrFVF0SIG+C6LT1Z
wbG5q8D9TU9WomDif9tNGvU7amAd6+w+qSThgJeZkSZiM3vvHIObkjST4P0pHcPq
5YCIAzECm8thVvK3czKCydyse8rjaxzQUpEgtI8vQTEpF0T2+XcYyKoyfaWnBglY
1ou24meo1VSX5C5CX0ncJx1QIdr0UGJwEllpiSYg3XfPJwKmVjhCdKFdsgMut7ko
pWIZjrrmNkouhBWaMmOV96RMvfQBBX50n8Z9cN/L6Syf9zCWWjrUZu6yqHKe2682
kZNxQKJLfJpOPR/9KijlreRMxL66b43S8sZSF8j065Lze7DuuKWtU1kj4ozgSLJp
LCsmmLH9J3hHT5US9XAw2u48oO64WRO8lD/6fnjV4JJWGdSV9aAedPWgTievXLUs
7UnYetL2rLyFqME2aygZHBIGE39Gpxlji91A6VIsRF02NL7WDftDcBeekofJRxIy
x1cSantg/+3H5+9pnwtbaO9PRB6/X7q7l4E12YYjKtgY3tp8RbRFidsj1wQqp+Dm
AOJmi1W6Ge46mV3iCN3cZ56ZsEfDgkJwNO5nblxXnZebTcPwKT0rpbqaQC8gbRo0
mxksUGju36YEFvAzk6AMGyN59dF8KGuUiZmMzHYDnGQQqDcUlnL59n8vK4cghKNB
Mv3+x1GbsZSucS4yR41MB+6wzBjVRlFdqV/vEz2BB5GeEpeuO1oo7rruWC1wGF+l
Qy+Jqsy+qpFWyNCOmcl67PPyHswyDkzLNF/cIH5chCuAJXhWoO0dsmVgBOb+Cg28
xOSu7KWDHTytL/TSzWMQ3j0xC404gYQqOCY7B2l4pfas3ZKCQzmlbxL7xbGj/Z+X
4siwTNSX5gwHzIsgFaNA6Q4MWasiliUP9+CQY7hAjB5EhaBWLoRZQswr67EkDTTU
OvlRzgMHTTBljVTKGYYhIB5I0vwGQgmexbi9PWmtb3dJKa8nzvB0hdMUZgYdct+s
iLe1xhDprnueAxaUM90wiJ1nyS7nMxRu0eDR24g3OIkTlyV5XwwXSrYPQRJhWRwN
FRN0U5S+vRSqFonNBiaXbOxJ3eEMny25SvC8PgBFIc8K8SdTUkMq9RmBaI4EKJMY
htaAeqUqAYKXvU1HEn5LXSamkk44rrG/xZHsN3rTNEK1Dy6HN6N3SWaDBg4FAYjO
ghSmyxjYH2FoezLCR/rWi8ujQkRH/P6la2oh3B5Zx/ewe1HanHA0OrNw5W47APUi
lXjcMJkXncE0PL3EKZwK4gN3wd4o9Ka0m2H1npiSAUYSNAyVcj6Hyc/CLCDyNf2o
HI5wNodNZJGde3Rls1quqP2EpX26nRCy7IYW/pgB47sZ7TK+v+mz0oCZ5dMCW0Ht
IQCNl52Y439ij0EoQeXGSgXpRGFAGGKrUrzJPPsKEmBC/SDh4S9HrvKO/52nPcVt
MAZXgh5TuU6c9Nj15ft3ljqWnuZpWA58Z+3+iaEldMaLgn1g+A3FOR9cn7y/rCHC
XjN7b7RcK4dagJsj7alHuEQZ8qPrt8tZjao+SFsj4UTTS73ebXwE1h71iLbhrM5s
uhtPtIwPBGpo/UeiuTuxjL99UxsG2pX0/w3qYBZL1RGy95y7JoquDUoLULjT8hbM
GIYmuyz5C4WU0SGDDWfzdP9brtpf4oRMAAlu5VmAgKI1kE+lbUs9NPbxOdI1T8dg
JgS2sJnhfTsLCeTlusseuZ3CStvPm9LLCcl8cv+W1nStwt/z0PJwA81Y7v6g0P0b
AEuqkKrTrqIodjpp/KNPzmOyOltfzWz0H/cRZz3PHThaHe0rB9+ToXgTjNxOIwTv
bPiw54cNs3GXN7uXAjjbKy3Vg4Qwi+TnIJkkijvRZfDY585X+3k/72VT6yEyuPXi
`protect END_PROTECTED
