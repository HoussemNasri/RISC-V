`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jsyQnZvj+bWeH3Bamf0ZkjOmNzimBKhPNLtFZBfeCYmpWdeoF4BVEVoR1Inej9AL
28Z4BQX+vZP7/e2VFV1C6UuQOvr0PSFutYnzth7diz34GTkZpq7vxJHjgi+6xaa7
qnbnFmY9GZVyMAeWsslCoWNWt3Ssnr1sP03rbUtVY4QIcC/6Q2PI+iAjl5rQgL5P
lVJweUukX6itASaJzRU6qtQHWbZ3uormHICBaG8XmtgersrnVh73ShZ2ek3bgrFj
cygPeoJjzJMHCwdhm7xdTP20CyHUa9S/S2igC/U/06XHs5/+FYbE72VST8ae/KMN
3Eedr/rh/jZunqm56jJ1dHDW6tR/ox2xU2x7KEycTBs+LUs221cF4XAfKGjaOhgd
4qQsUaW7FotJlFWS5d/5ZsXCSnG+ljOG11K2/X0WidKJSJ8RRlf1AQxRyapDmRrp
hhBshee0Fe7Vc71Yxa7MAsmnGd3bZI5V73tyL9PSW4cdz81yePyWK2U/0tKRqQDQ
DcX2ara8mAXxgq6MlPbdA+Ak7grZwRik9V1YDQAwSO9zglL4VZksm3iFzDZviUkX
8989q8vqEOqJV/jog1H5s0FvG0Bs2YIh3lSR/9BikdEEGaEMsic/stOMIaDu+BgW
XAMMWEyqueQNFBdDgXm+2VpAGeGaYDfRxqk6fZO3nrm0/irQVCJe4lpRivuks8gz
Q+GTc/qaGCYvngZ0D6Jgg35BiWNycrQIqiITSa5kS/6XLpHFQcIzZljCKDsPotbE
sogFWD1O0G2MKLhBEYjKnfbuu9A7OV/bSbd8HIseRHUUyo6Ua2MSkcgmqt0o0blf
Zl2b/HG+vJbHW8uK2096HHzFdqIUE4T/NRsr+741OlmFpXqvhNFkWJ97LJuMg6Zu
ZUF2PExTzOBlrgqDJTyhz9ETb6oedYxE4nfh1feYxmEAePLBD1wnFccuR8qgep50
HEw2WvOI40I8p8Yh/epycZfJiM61RSqoD868uFOVI/N65syTh4qJ+LdPvUEHmpGV
BiGG9yIT3p7+CXV3FcCNmRm9LDnr9DJrCq9XN30c98qs9DpvMxk4P0miT8YGnjZH
Q15rjMyRlR0awc8CeM8zztgzDt/dCsfe07oH3JL9SXaeEWKKjvcs0RHDQ/+ZZKZq
H/sWWivvPxq7ZZZu+T81K0zOCW1bbcnJX+PH669prvEPwrspfs6LszYHFfz9Un9Y
guuuvznC0nI9ngrYxswF00o/tXOM0NIojK/9JreW/UwDxS1A/WJa730qxl5ILESY
SJ4LIRD9IR+e7xUz40K7f6fXvR+uaLAglYCbrm78phvTDtYKVUbzQ3vYbDtwshYj
8vA6PjAtA6WfQqunt8AW8yomxgNMTuOwpv3vqZ+17kV9imcAz+G7ogXSqeoqV6r/
e8SEelxxroJmtCVLl8803M4XJCYxxkbsXbC2RenIC12wAiwSK/LGkb/n4OmtnvTH
HpqcmrGWWHzsa4iEga1f12L3JAvwIjRkDKou74/O6+oAIa80w5RGYIwrPa56JWZp
/hS+8ZvJ9edAr2BvQRSrUPU4qUTBs/Zq1Gj1AdKMyTm86+fn6y8hItJ2C6N3/ISP
rBIvkrxhWZoVekEbFWj4I6g/HbLmbOwGkVkceIyVqmGO82sPyq6IjOtRE331fv8b
bwheoLkY9DoNPibus7aGTnT4giEOeZtdSvdo8dWDd8o223MHRHlTBEsAmokHKyK3
jnkNhsczB8+uOs33GHt0hr9bF0ApL/4uWwqAZksFjAyznry7gqs48ekSpq3ds2tI
l0Wss6JylWO6MM72V4JCleeKOttlN3knebiABYHhQf3Tcci0IwsnYk2rcrMx4gtV
G6R/4Fwwl/Mf1rLsQ/AZmkJDQUIa6HuFS5YQRVMU1KoTzRiBbVR/f2NnNmzQpoyV
MtkMDATL8XJEcqDH+pd4IRLgvPDM7HhnasCVgsdh3NG5ssODamiuKll5BSnMUlTZ
jrL/VhHaH+akB2uYtGxh57se27SK7r4uIkJX5WlDdcBg+1Lmfg8MZp9o2bd1Y2rD
4ISaqTrjg/HU4TVp3ahArh9EBUgn9jPZyv/4AeRrcSd//MFl/cwAustiPVXX90MP
bHUBgnU8LvWuyJA3SM5jhchh9aNpYCVxp6S3+DSSBY24lbKSngGmsXhZn1ZhOEtu
YFmPMFUu7acY2LCxe8YWMWrzokyLe8Xp7kqFWfYCbbg=
`protect END_PROTECTED
