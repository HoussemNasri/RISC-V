`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SR/GbYBlyqb4B8+tK9NvNRaSNqIN6a5p5OtITRjJhsiqmHzlsXLHZexGTu08cTlV
22upwKlNSwpy9yCZO3NkeI9rVdd3vsD5d6Nvx6rKhL0nBvVcZkyreJQ85vqDZrTm
3u6EMCnrck9jJIiynRRKFpsI0vHHkS8XSa8FBPv6RQr3pqYntuEbVsXph2Kek71r
4Z7Abn02wxCX5EaixMf/dv8bxVy9nNEjGUbWjUO2z3oPHwMAd88rqENvm/DseOqh
oxqbTH/Oet4vMzOAhTmC3Y3wV/MXk1dojatf3Y269yvs1cYYdlC5yOZP3nJmLq/d
nrlJxIJFQfAfmwEuZGLFefccpEmy8lztKVAf96kM1Jd5zaWmueHJ6ZiUYaUGerRN
BWhZqz2Nsupub1CWbgpId4GTasQ0jHfzo6tB6ArDnuIPMQVXEcgTFrbNL2tQ29uN
w2n58UfLLdZMgZHbu4XbTWNPGgdn2ce5EGPUsyN489BMYAT6fjBZfqhl0VA5B6og
+CjEcHrSYGY9IuuGQwinvAuoOtNdfmdyzKJRDjcijbiAfys7tJwnny2/cyUh5hgP
/Q977omUoZ80zKreSCh97bxfp2jWhO8sgIykbkO/8X0S+EtHrUVxAdqd+MjtUy+d
8MpWWEEwMIxZVFOCjJoOIL2KSbKuLOZlJCerFoIp6FMTJzBQG9m+rf5VNq2k2l0V
3h2l81H3LRBZI8OOTCUmRTQ2hnJ4RALGXD91rjt7Cvc=
`protect END_PROTECTED
