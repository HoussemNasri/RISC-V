`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3AH/+ZZS9a6UUQ0nUKWKLMy6TOWJUBBj/rJl76UxVqSH/KTKhBRtUTADcBv/B84v
QC85Url0yxgxVEU/5o2cKTcM7jGvnKao/B+iAhQ/IFfePMeiHOjYgrrDG+qE3+1r
RUsdXjgNdSQw8+lSJ5W1i0m2RGWCeGi3vpcYq2eY1rNWjYLs/reM+h0BaPV6Wqlt
yZhVcygZdMHWJ6WRNngWQyywfNZQx6NC2o3HZ7rLFdCl5XUhMHThefy2UvK0TMmF
SsWWg5jcHadWqsgzPOYrfixDhojkFB100Zw6JWROvhoM2L/PVe5GAMVEHwcePdsH
g7tAkdXdajQcMps6ax07b9yDBfSHQgWZlkFg9UUxSAcdknkiPZxzmqp+YoiH8HGN
BaAfaXg5gO0m3hzLGUcKjGPM3Bl0ix62C8q8c4SaNvkUSoX+Uh6C93hn+0pWqRJt
UOzbL6Qxu3ccSua1JxpC6cJNarAgKSUoNbwaJJPIk2thRJgOlxk8fDoMUnTjlwuk
iNSbAFnKgQPZbDxSViisNp8faAv71yJqiZv5J+XRsGQLp0roE5W62XUot4wcgST9
PX4taklt/2ri0yBglzxYrKjCNGkcpgrvH6cNzIDNOhuWRjZ483I+g4PG++7KYVNL
7IUK3KERBMgGlhUau2F6ZASlnp9gdF4PU3eOlKRsCfUFyfm7mk1IXr8soi0cor+y
Bj8EBn4oL2RX+UKW7KH9I6qwyFEqt/Z5N0pbuWej5hh1Y0Tyybthlvk9OvfdCr7t
rwZgIaK9ICY8CFJEP8OrWvcDwhmuVj5moF3Lej503HtsK/TwW/OfSMb7LrN9ro1G
ziD99pBkEvGotQdwZecvfzNEGuykifbwhfrMTxwQESvmKUdD4P4n6heALkT3yowB
19kY5GPg7DooUPg3iREjt3nEktHstRUNeuSlp6G2yhDcBGguu+MwFJEOdyYDw/X9
XPBydJLO81hwQ7p0Cc+GqfKgwXHQVHBXOsHfGeZ9LdPQCxDbYGaN+K2Nqt8NxYMJ
+8ZqoCucLctwkpSpmD5gzQWdgytGR4fACbBeW532SUFHaisgI3O6Zw13FUCXXvxX
Imo+qe/zZA6WEs7lhB/uflS4KR1QEITSGQPqA613mPxKRSYKoMgOSgGWgiPHwpT8
Rpuq1kf62iiZZi3aEqdeDpdYsjJKPYkMp0lh9aZNl4K1Cea9roJQA/p3o/Uwu19O
iGGtOp3IW2ZRuh6oEbkpxg9xO83Gnaygsoj0f3L6f+13eBxt4yzDuas9tlmFQl+a
p5WKFW8JqaNUFN+NETtkiqvPHlSMiGFU291pXcvkO++g62C7YKO6YJHfJq9v48eb
muAOiPIN6OqyOTEPYZqDRJEYw4szpS1Jq1BT9H4dZPU4QiPXE1CIRQrsNamSPZzp
zLs53RqhNFwkNpb3DYtS3LHxMGqDQYH6HblYbinHv2HKb4jF4zgREvh8q2jWLNWY
NXf5h6SyrvQ86mPNQlAY+4a68UcsAt+9OXQ5X9hWOeWS0lzFk8Ykp1d7j6bLJAGY
kiCpsD9v8QtaVTS9a+As96shdZm2l+oX3PXxVUhKRwimVWV1j91RkcAj+80KnVXz
FlyEm9PB6CqoDgYQiOBBKwXt+fKkgKRT49ISCoQyRvruYRE8JeMZtsF/qppW/aWE
5P5meaWwIWHle+axRfMKvnFZ6PoRBREc7kP/09Kk6kGU+Z0Fng9NfLAIbmBJw0mp
KJkVwy+GsioskGYuojYTxXy/MQvPKBgq9BLK9REjmEtQOcmafg8zvuQiloIj8bAP
sEVJncYI822ESNoSbHIQuKrTVBVOkbLk7qVMFt80xtdZt8LpWidsmHK/plc4AyKk
4yR3WxK8yA627VdndGrMw2001AGFN6SrSf116gwiYQLRx0hVT17CqaONp2tqi2DK
8EGlkIDROH857zuU5GmR8f7jMxnFwHcd13/+SYDmfVDSk5+XU2xGuvW0EDDGefsv
3iqOtgvuH+2jHFv9fHfLb4v+qC04UqGgnJPzJZf1GO29q2BZ5giaOSnp0+w0n2kJ
Wl9PD0RiX1rHOWXs5+a5PJLrcvP0Em8WQQ8LLmnUSPj7KVaDygzDbjd+kN1hXOWh
m6dL5P1TLx43o+b6bOgc6uav5RaUm943gr8jMoS3J7V3icA9usrB742jtFwmJuMx
nbXvApkmdpHNHhB2epmdaq6tmWR3Ao5ZDIAWqzqxlmln9oG8VDtRE7Ori93JPViJ
D+cyvrLvGj/FuILIH6WmUhyIfuhmTYqE50ug4pvjLL5HknBZ8hRSiUdez8IY5pF6
lvgR3cZqxR8f0e67/GTXx0cCUvtsZTO9DO2h7ja0Rem1Safl6hQb7cRcuN3BRe+O
jxbV7+SKU653QsCLPNjRiNIWQxdUyMn6OWZdES76DXcX+Pp9miY3H+TFe4l6LL2K
9gT9DLGKCnaE6XaK0Dfh8pX9zu7aZKl9RnzwkNoVrw7UqUqtN6w6bpmipvRfzOUM
cvblcmmodz3Xozj7OT32i3lH4yeQcplaYrxvgwsswlAGaDX7M3Cc/Ke+geR4uhGU
C/94/N9j0PEJAPJZawYQUBEjRqxXiDs5/k+PMSyvUu5lvhO53fxxiBpQ3WMvvBHS
nbXGBbFQeYer/6dZU3Ii4kvFFeNEgcaiGDS5ksusV60i342mitrlOi2ArOWAYAqr
MFV/PAtRlXzn0uQhuVaXro2LixFGgXg77CIwQCE1a9YatoA/DaeYmq3z/b1QDbem
wp9frIL6q20KtdaXlg/X+bzmpTW1/87ACL7NT5L+NaxD0msCbvzg8vZuFWARMobF
6vZGzQUyPQ7ohlFsUzSywcP/Oa+QyWmZpb2yM06GUQiNuUI3x1Y2hJpqVZ1g+vEG
EvYG4PObSizoNaIlibZQ4eTgZkW6UjKIl/vUi/2lgyBxEaeyIU1GcOOY27qXGPKz
FfXnoX68vlYAP/3i3TpDIlCzbWg9rhYP56FvCg6fVFFdN5LmmXtwChf0pCj0VJpX
RtKDTPJ/tiNsykAA7aIOsjiZGpuQxUySto1WSaNNttWtHck01ShT9OKYio0E8rXY
6Xi5fxwodXGohikp6/6tKD6iD5ZebM1rvFTZgl+cKKgXDIq1lq9MPQVsXm6LCvdZ
xx7OJ7HB+3f2EYxqTxHGc0dphqNogxzC4CyAq5My7NLV33jp3Xc/cFsVSydRQsUZ
CapPLRJONU/4oaHN6bHr3dEu3mX2I5cOAwk+LGlMoPXuVOlgm0Lnbagaj1jT+nS1
FZHO0NWTV6bwXmXnjM/UFSf07vedR+yarEAjpF3dDUlEli8Dz9JNOBRcefxK0uky
r4XsxlAqI+MYdt9M0Swf/DzrUjgh2SkAfIjwTZa5xZlPqvktuDdR8md2UMcDRuCJ
YUdh1BwwgwMsK/IvgCCCkcA3Z1Bdph7875KYB3Cnb6QWvfIxmWjhcDSZ7DnRDxMJ
4VzqVaWQo/+4ppZpO1WsRpQ9M2+9Or/RwamIfpPxO9jsKihVwqbjoO/43nnK+ki2
+BiHxJ0v32h9Ch+G+XQ6zXZQ1DMG9KpVnJhnOqOCOi42HEgf3OJ0LskF6tkcACoy
QNby/D0Xj8Rqve5yPQD9HcvOoxuFUsSxEdB5s0YSlmaVDw57a0i0vSl69KAALDGL
3PhUkGhxTK+8+TinwDWB6+OKO644BEKLd2tTyu0oDfqkEIHJfW+WshuDmeyAiZEE
aoGX+1blwxTZ1sQfH0fiww==
`protect END_PROTECTED
