`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJsr3mL7lDRxdKQUDpmt1OoAqCrpsYkAUh+mInRJmbhFYshkQlBI1tI2hQFgnV1o
K3/IktcZAV8u2uFY29b3pkl5ZqNsw++hKgrMQYkiMEZtuIiW8tmgf6AaygRQbCHt
jaiIkcD1o+KsDsfZUmYREHlyh/gJB28k+vSKsEZiH8Y7n5zYNABl+66HAPcB+wU2
TWH82zfLSHG2O7kRvNiSw8QXDccMAu4wvWFCEzHeDBDObmf3NF9iUJvcijA6eEja
6R4qTeBYQl+7LFlAk/tjNoQVfnBMXk4Qh0CmERR2Qc8+Huy6R3982Uup6mIfojHA
oxOv9U1MlaHIsQHFSCmsuaqAd3/bj7DeZeNrJ3h9W+0xiYTz7gf8SHHrJ/dM069G
E+z3eQCG2EpfJkMzKwRVPwcnqOqym4z21Oava2I77lmvqaDBm4ScHjNulclIgA6m
FfecGJx26k7svos61SQOgNUkir0bml01E1KI6iszT65AeR1L1w49i2wKTfpvYrV4
QyhVD0PRndcVInLRcaaZeYXZ5Qh0knGT5mg2BjziUumzdIqVf9U4WFugDOe9VI6A
sE3uVrujSgqv9WiGnDXTYSagcx3PHY4hH1CuVIQ+P7iSV1kxTlBkMc1kwJmi7Jfj
2f/pAnPqf/4Kras2wpo/KQTrrBvMDiZ6/YwQkdQ9W6Fldzf0kusre33jF3w/gFan
04N7iGuds8Q/hBCXpHnNW6RpC80jPTKC646miPvsH0JeTA0rEat+VS9B8UcPYfZ/
WyFl2B56oXsvZp6ckyDGkGqqI5g9xYKM/sDY9Serc7wRHPYwnjhqzCaMmwOzX4eU
+IJ3xjsss4Pagsv+Zq4FDiCYE8DLBfw+rfYnrC20A/l7rj6RH+WtGcJXDgErp4U5
BL9PR1YIlvXArN/1JKSw3Dt7oqz/pIIinjAxg5yqlXoX/jWgswUTfy2OrDnK3BEr
0Xv8jeFmYSeD+ChU6EAbj+lEh9H/U3micbBT1Y/tpSLZbxIf/712RKTVMQll6YoO
yfhAl44Bl5sf/bOfKNhNM3SktLoTpEfcEEcZn+tWkAbVXVYSgR08WwzqaXEClXO0
DkSqIknASgimIZo/c63XloRoCzxwK8175Ma7NgfPuHb0DWdq+OHfJgumOajw9oqF
ZQtk0cifFfsXXizpXJ7poDRqJXSlk1ZkMDn0zVq9LxG1gLT3KB8zg7muNypEpZIV
TsQMlcbCZ+uwTXsC2UgO+U5qQ70Vf8B5YL1cOvbFdZlsQ6zCNU9UAYGLnemznTBU
aLaVn/SGfki0lTh1etQmO6jBcM4xa/p83CUy3SnMOKM+mVV+VhfycMyOpm1d5CP1
CZZnI0lV7EeVTDs3nsUCBOoY4OFhlVcWwGz6F/q8DG5/V0EdlpSY3nvQ+HVBPKh6
LnO2d5sxGuyceiOTTUbwL+4EX37oiNmlVUqUlsVNnHn/xf6vmyTtuwSK3pZMyxDy
X7HL+G2peIYANnigXgFSe0R8gI57LUAQtoanzDSWX+kQ1n1fQZYIb4P6PtnkeUL0
nB3sSUkUxO3QuCy7M/P0xcFk78akZW5YeYeFuWwKebMoEaz9rP3lUF8pdzLiJv1J
81utUMrfQ5UVt5kcQEO/gmxS0uxlfxJryZRy5kiSvyUgeL03fNU1v9D/4ee5L1D4
QVelWef4SG1F8ZztlOIxsnQxtnAjY9u3jlJv9GDlLdMnR/mYtjAcI3+mZMZdKIeq
WM9440hD3a4as+kYNWf/96tZ0hJQpM1UmQMwdXSAaa5UOVRtgh9yRwu1imWQz14r
3Xmpj7rd8l80Tm5EmQohIyfahaAmkoTdd2ox6OXfv2959hkS8U7/Fx8HWUmoAxc4
jsph/DKb2TlMXx90PrbePO9pDv7At/fmDyaZiVavVUdMrvluv4J8qapd9QdGe/Ho
ZMmE5L5zmhCos46Bn3lpAKl+KpBhYVm9xxnFfQrwgt0mMnf620Dg5EKh1egswD5c
Xcp1gP+zjai47DeGNbvlAGP5DCEaC8MSGHo1BVz69JHnsvUV0vztmpKj9nwM0FEv
yfNuFvbp8W7XeOb1FIXGItWHix9RUM/ZX8m4ryPkAKe5q2NnV7hFnc0FhkBLkHik
vxi49kS6FvRmyKRJNlE4XySafFkZiu496sGCm/1vSjIZ0ikf1BsO4A7h/MVU/3j8
+5heWDqa9i+CULuptIaekihoUxB6zlxHEJ1jZdIesWkWluJFB+H2Yn15YvPodmWl
Mfrj6ZlpvqqCP2KcGni99sOlWUUlQDWDFI4Yyrf9K+P5G7bUEU0Xos7Pi6BBolyQ
5R/3vDqIjK8AY6cdY16mim216THISpFMM/rbqgK5xf2cIgLY6ItMDynEOikjKc1+
eNcnj1y7/L3w0fsdeqGc4H0AMIIeYrQuPxWXOXp0ZaOIpJ9JmfAr8+JdAont/vYR
eHNY7Cb2Q4zJ8Z2S6rsMCD8iossd8Iw1IkWyClSAPdvnRxYV2IHSrwLMn+td9ioS
LxNfJdkMnovG8obGTY+MOse85XRADJcJ1HK7TBc4mfkxxHByHzMbRAVwydtizeuJ
C1MSOg8vkDXvi5cIO+zcYzjEiHy3/3PWGQUeMjnePk4SNsxZT6fPZ5/abX5D8+wr
hhU6s9RBXcWg/bB0aLEUmrsOT+JfDPHL2WooNKzgzXqzqyADZ19TpJ8FAvTbu4rv
eJvMXoOCjSmNxw9er1wN7b20GEu0uUryValbdiNr2uzhSi8wUJxPwoI2lkCNWQoi
4VhwpBTWSK3ic4mk1N7Cc23iTLwA2tJvZtF/K+FUpQA8bBg1kUBh7GkfFkR8NE0M
VfqXaedo7CHnNL6DkyN1q4H1axBchtJCSlmwEpXliqydiWkl1mxPDiOWfxVam0CZ
FaqRsSwHoVsCRooar7W8UxOVt1Iq5TK06354rkuUw3hA1OAhkqwXHh/uqYsBj3ZC
kz+FbcojtixJPHkRGwShIP9sJ/EaQYXeVCW0dpqYH3s6On5kENYjrQdVOAiNpkTy
FVzHVfU6nidnxIYU1Td9dWHn609dxLC3VPCJIdy25/iZ1sT1wjUniaVpIlmfEQM2
2Q8XtZ/AjUEWRAtPhrfe6gojq8fNQ60jif5d0Io7DdxavLiMew0K49Uz3LSzHFpZ
yw8DZ4LOb18Nap7g8VySj2dzk26p5izGWGrvDmHx83h/UN6u5VE7KHPfq+noI85L
XCVWsAlCxfEe7v1Qu6+HxIIZVJQXBBozdlqtIMTnlPh1mPznzCnjap0eppCJoFcT
T8QGZE/PO3tSOLil36D7rTJJ6+qKOS9qqmc5og9P39fd0GI9iYJLrSu8iiZSXdMM
FzeKRxNu+/twz5lkuLX7EPO5r9UuHeITlCXLwmeMKxCQ/xLwZwCQjjvVNPQHIuJR
OZjpjJAAxMBOiN5X4MKsU56Vp/p7+OGBvAw+PBoKUj8tt+PmpgyymuhhnS7ynbN5
/mturxmOV2DBoEDkrQQnSCr2GtwobUMKqumeKcdK87HnFTlquV1WKINPUGMeEwih
euDUG9lLL2lGxN7dkDqpVUnKVeP9Mn1PeyZnQeaoBN2iKausoCJWbytY5pGRd2Qn
Flj4mtvV3W2PGG24EOA4dpe7ncNfqCp0Zh+9vBhQ36Pe/3YTrRPHyW3iLHdsE3Fj
ZLUTotMYmf9jPf3eLx3WUVW3bT351UCwEk85+ixYY1ZVQmaNqhV5qGZ322ApKHKv
Iq1WCK3yRwZ2bLJZFiAcs3P+GkTBRkd1+AmJcLJ/nIujTfz9QxIBpHbCqdLUtY8B
QSbLbfC+XOWH7luiDu2iZrJ19K+7hjMOFTAAccGNUbjS+aTroGLOFQM/yAMtUYev
/RyGOU2RvIExjfRzxIRqhSv+uTiwDmJq5/8A3fOLCVS2JXEce9c4n+nTWH12kDhW
WGwV4sndYvwB6WwgPNf6ZsKWLqS0yImZt7QjUAUIuGiygH8XGqy5kzxUkp4cRtTr
OhmNWc+TF1WzS1grTnNXAkT15eff2idUOKiT+NF4i+jA23iQYh3NaXwi4RIULVbp
+m1p5E2daFHvPnRyYtGn8aB97EO+qQUDwrVy+BQNVPtNb/Y2vexeYXJhR9++631K
p+SzMTlxDviaDb1/D07eBTBqAZJ8Bj7GAKjaCUc3rWpuQPL26ZpSFRClhXCnhd3o
Al4EyERu+Z5dj9Q27Fvvt+wQds4XuIzw7y+0Sy2xZRVLvfVCQDHOFQlqX6O2yHDH
20qfjsV+1QUf7k3ccxZnSvykrLbQMp0xKvQGtx9dBVYQbtGmzDLCznVAWXYKPJt6
KCNlhsp/sdFa00Bz36EPBlULsZVFQziYhjIOCav94KF+WGpmZjWqPzVOCqB04Oww
4gmTGws5rTs5M3b8gYI4OoJLsK+TrXtWASxEObEfjaekd+jGs0w01UyBUD2g+u9F
c7s5l9pvp951PafEUfvXfdBsaatGuEvwf4hFawgYcYvuwWu2/s+EHhwjrls9rxtg
ZcV28MsB6mA0YwDIRVehkKQHJTKMOFzN9mSiXJVR6BOWf6O629CJ+d8+I2U3qRBy
MSs2LR5hEM8RyBuzx6t4yH20bdSTIT11/dtKP7GsmSEZbPRdBerjMO6QZWaOCd31
QEFzJ44YkLtxiKvKWL6yl/EDo3gH3u0QiyJOC+h2B3xwMHp/qlhRSmXxOoFiVBvm
nMCzGapxgXErpfP4l6r+Jeep7dYJW0Bb2LzBU+e093dXXAyTr0+mvpRk1HsgL4XC
cHszbzQQtCOPMCeuUGYvhF8gUn12ryNIMYHuGoi4TWVM3/HmjSdZIKsnKDljnxsV
V1FDJLemiI3RDm/5i5jmXXao+oD7EjHZ6GAUO9gOW1mSUuViDufwWgfwLfFLzr73
xak09OvTFNDnAG5hEd7EcbAC0PXkkJonEdoyP6sOQrTe6mwPydEIo5IYWJxZX6yu
86fg159ONyNXeel6V9CQ8WuAL5cv46QGFKR2oDTyEOuEUGX5W6XVBJGWtjXNqWO8
GePVWQ3ZHugkDIsMDwM6Icaz7h5CP4lLsnNsNaagoy0aqXxjkHtywQy5MqX2nqb8
nJj0dLtE76as9axTGq8NLh3+UCZmHGSrbpj1Ds5PGpUetgSBopobxjg3PDCOUQcp
KMmcTXL4TICs/wt22X6TPlDj7nDFYFcRQo4CfbB6WSzH0hbZT1rp4w/eOcVkobu4
KyqjVaNOX2ItBt54ylbrc4sXzvWb3WANyBde6NmPHOXZx9L8sS3sB3v1b4kq152R
nJko21WPdQtT1PE+9NGAisRjBUVEtKLrlNoJMAbrMhUF894ooOLMZMpSKh0x2qOY
HAk3dtzSbcxMgKWi8nUZW6+pNQTzupsEMsLoIq6h6CK/5hjbi/OBU5XPPgsdn88w
AOiRMlEN/0q0JEwaS7S+fnwiJPh4Sfthg6WTjpBj1kA5rn4SSdxDD2/9j9UqzXm+
D3C6t5mgyqm5yEVfQjjPxW6KQtx5x0CFxsobKLvFOMQZ8QcASDgTS7atUoTz6yWU
4xSi1Y/EJ5Ie4o9cvNMJCtycLCYbtUmM9jGqLfYI6XD/OgYuvsGzD7YlVcce25cb
81SYroU1dIY4nfhWpcBW9p/RW2pm22Ai3yrZe45Vm7tA6mYeaaxK/joNl0kwppWK
99yg/B8bUOgyG0k8qwxBXhmChoka12iohq1kvQi2itaTmjxAH6S5OTUd2gwV+XdR
n9ErHacaANpeJaVwtr/xXDTWSKyjhlEFXp/FL92n+3XvOGmLZ99UgeWx4TE50jJZ
YXyj33YLhtXo6SXDPeS8+mhaUXHV9x3xLFrlhxArXjwtcNDyroqPBGX3dItqDK9j
sPDIYnHj/B6gBdYkmoakprN0B9KWLL5cbIve9R63ccntRk0vCH8zSStalRXMMTxQ
beuiceaEgUYR6ERz/U+mVzxURhgcXW2RrrCcbCe46mRvF6DRWhAUHCKBP5PdMP8P
ywjzHWNClA/uo8+5SuTeFFThhJIDoEdVk16UZ2rSFUggLHOoGBHe4hRhyorFt2wP
PgYgwAi88MdM3+nY/8IQhXQ/fag0YXPtQSs41Hlme5wmt96YUevTptfBbjtd4Byk
sEGvmI8B+bqYGyw2ym3ZPXzLM6uitUcHGUjNTcATNGgCtAheN+1a+xHAbE5pMOnl
CwhNu78oGbmWB7s2vli77GciPhJW8QVACrt+HNRAnXsA9oJBVMdwFqF8oWEauKk4
pS1PJr61HwjRnwpfX+5wC86Qf3+UnOzCJ4TRg8vEsad3vfaANJMocJW1O3LVeAg3
bTl/lKqcuCcPDpTyNM3g4KLtbIWITsFGlWp/fI5lgjM2IhbAVS1fLslJP4fHwOcS
w7lSSEQaTIVwZihYADkGE7d6Rh47h+7ECHw6dvIsdoWtnbVGBDieHdiyGDOrVYJ5
x22TBte4ljuubtyxUDU1/XNlfxJSDDE6sIJWg+KnS9LnAKZhothHREwuF+hAVS8w
BpiYjatTsLVFqR64yZ47cmXXH40NrJArzfdzdMIHbPWg/d12yPpqEA1p8oXsy60K
J4j6IGBEip4YJYWMgIFUZX8u5+WVAIzQyC33DomXKtn14fqXxqpcBRZ5eAm2fGKP
O6Cw4w4dKr4asiUNU123b4kxO+ucK352D4Ei3EkcixfQVW177rnAIBJxw+J+P4vS
wLggjfu2VC0Z0USoPhPVDlSk36O8HsyUXz+PkutwtiCHFau5i7MIAtMh/FMpol1e
BHFqCyjbWnFFTD2ebS5Yd4N5cLl+ETpmQup6hl2vEXdNQkrVG1ciux3TB4wvzYrl
fZ5BEzGbfuPTUnreh5Dz57ObQKeod6H9CuzNNQZiynIAvNBfSvcJda/dCqUz/sXh
NKklTgTqbPTLY8XOW5nhcLZAao7XlZP/1WkykM+qhWuvZa2rUMdZ3satmvCEuyBs
eaxmN1TATNK/yRdbTSTdjlLjw1kSuAQvrOekz4bfC46cN3XL1H3SXJXLxHXvcS8J
W+CbKDts/g8u/HbcyD76PkXvvlUl+bH5+w6/JHiniVL7tjZOugx9l8m/gf5HjWEy
IXN4Chhv8teYdZeTNwygrQhiry2Denwrtp80BbD9uiYZ3jE1Tvg4Xpnj5l7GYdDV
zRPzi9b16KIxsTA4blZjmK9Vzlv5o1wxe8uNcLX/hqU9ecfnfUt+lijitYNJPFjJ
++TX8t49xLw0bvXCbf1Je8r5EEz1M+hfAwFX+MNIOiL/4c09fAGZ5mHvBtAOSrUJ
vMzw/admuwaWob+KQyKzz5L3yjvh3CVQD2C2SKgagUMf3rmwI1vwPeQgcwtGjxg+
CmmjiamaRGsn/+IZTOC45TPgRumCh0rtp5vabihrad3USc66WlBFuQiapDxZAcJT
8giD+RLTjaY9un45ELmK0q0W1qWoruf5btf5P1XyEI4CbBw04tc9ZRCeibfvsuxr
mWb5tgQE4WxlmfxarTzEA1Dfn9n93m7gW8W3nG3wEfM5vybCFW4aLv6HPlwvV6qg
1rp6WiNwG2OT3+yR1aVO0MHPq55hJFX+gZML6aOKy/CYgEsCoOStXJJHfJU1q5kJ
UiCR81EAorxxSFFsyjmHkzy6yobzs0nT32+Q9nNN5CxEFNQKFi2F45hC0sZbulYF
nabaNBard6Q527zMBYhcFuCYZDVNwJpwg5x84e23Vbaf4KHKzFIVdUXerAtDfz1A
VZsOlP5Flh3KsQsYHCQdCNrgCgEkXaELpEf6w+baMWjsfOsIyb2tZ9sDLqD1+0sg
+pnGQiXHEROss9fACG+RL5XY8w09GSTDOCoY1O7YeTHL+HgfK4oQQeeqV87h17tp
SZSyLlohO21rYldQ8q+y9hkZWOu/koMvhxLqvHtQO7cMnoMiNmHygYAPPkC6x+DA
9LDVg1O44kZSK+wb97RjY2rQ3GzKCq1EKqL+YydDPRVKz16U9iOfIG65NOyN6mkk
dzCselTCAOYEuOrQCENQELDMS2dGPqZVopyRgyHRAN6I7pI0+TCqJcHsCZvypbQy
vZHfOvkOexFPUtscW5Cay+dHqXZwfirGJuEsI+2J8AseZIxZkhLAKOS2L7uizGCR
xkPHJQOKI559caRPxIBG7cFfg7o5B0DPujW5UheX7nNUlK+U8tdfXsq690ntVoK/
MAGuByqBhh7oBj8gkgZYBffCqRMW6qp2tlCRn4NmxJo9RUFKWvzIVxbJysapAz6S
3UqOrpGCRx2Nl1LzahLeEt8sT+YxbYUfkHULf3h92Vhk5oG1/bHtZi5kBIGquVZq
plcQ11f3E4Kr2Yud663tQmCK9Wq0ZzoO0++35yqWiv2Yep1LUfPlqWnqtiKY65u2
w02uH6eiwAS9rIu3p2p9MYDb/Otmm3QhGGrwkBCV4Vp5vrMVGwMQx6Sw/+znO6Td
5a6VLRLOl29N+qQZIGyoFc36qlQFn0j2i7NwV7waKQoQiiHK+P2oBqwWfS+r6lJ5
E51oJXtfFE9USgafnHzXiYYpeJaqSl0rvw0zfEl83Tvx2Op2o6cv+1H7qWXDYrWu
bWascZSHOw0EVY1pvB1sJe7BbVL9WMAHS3kFE0WvcftlFC/e39TUo5ePEjBJ2FDK
czW+wkDAfCppt4N1C6YsEm10KeK+AcYHTTZfN1Z71g9NQ58lG9Z2mwu6McJz1Plm
91qwWT1kvWtThb+tIOp/0ssM+mTrUPvn7UDKr01lMx9ytU6aw74kTLJrDFC3QHTa
GRebrNxCHtg2iWTk5yNvQ6Oqn+G8iHVrZF/yDO3N3nL+bPjjUZw5oz6z9xQg9lRl
JX6Bm1zmb1Z+iZj0529X9Bfbn/Nj+cN9TrGQp4S/9elKcGjxKX7tRej+7fQ1c54S
eKDmlAPytpnju3GZpssRveQZT42kdy6JTev0gzj+AG36VoWoNTDMN6HvRds/qDgM
GCyfJUgLT+mgyMYf3Fz0I4IkesTdVlG/T5G2wJnl+xOZ6hs+tfBnnB2Msv481YQg
Ax1nJ2BmBGGchIh1VHip3tvBTHkUGJIYMWBT7I5LGpYvP7vGH6dn1AD7Ly3LhcUM
dS8DDEOSk7vIcZnkXjQ4JClo53okZMOEoh2xgVN3ys1DF/tP15vLMa59Z34sSM8W
YKNhxgyMLm+oMZ/spGfLkdB8AkWXZ2CpFlDDAUhWN2nJbi5JOI/O1QAztRTA7qkD
w0fu/WkXrGzCYagVApcoLulxERsBur8C9Y2MubVxGkrCCIKbmNhM6YqN2gpFQaBX
0WO32xdjCtCFFKIe+dxvWlU+963PBjrYw6/X8iLGz9hZLNt29Gw+NzDU+/qXugo6
bFmtNBM3HyLhbKGXC+yPYIuuW35IjOxpcqlEs802Il7MeAuyL5nmt8P2ftP8Uw9q
Qn2AfEjK94kyvht4i+1MNQsTABw63SsVUkkMl1rnKM0yCVFM4ZRQ5c2mALi2CjG3
ghL2i63n4WcVEAqEDemH8PFe+E0nPl0+8mVZKev9sgcODCHbDR0dyM3yHEwnoi5d
cn1SoPcF+wu9kqXyt9O52GkznW6cDCkP/r2CTXu26EuVs7ONzGsDc6/CChZEAJ22
cWNBspEEcXdWtttpB+g+oVziPUpSm+7E08JLw3H3+pffi5cBd/o99B2SKMi5jlZF
j3TkPv2h4fTpQYn0gkC/OVD6shOCGjiM7NXkOuT6kv4TGXbr86XgXjgTwOhMbuqm
fl+aGUoYbnbNS2bSnZkJx5DY4/XZEboO9jVhYPN4Q8PvDrRYv4bf8nGT02sNvorm
DlvtWvbGiNHFL/KtVtqopey7ZvqaLlefA5RwqmuQ9zauf8Wx7Mryf7GPLkOHAYpG
XwS7/Zs6X2xBvZAb1+9mXSc+NpqdPl3yveMrPGTOeVFT04miv4MJxwvPRI9UtBQI
t4TMzudMFIKlkV5LNg792/myR0XNuLdc3ExE/VxZegpVXFt6jIesLQBbtuGGh7RW
Ee7+hhTGKTKuyC9yt/TjkCpbYCy8/tHBMTHD2fGbqS4ooKV1OSODXwTNMAq8vot4
mw3L2iy6BtTw7OHc1Xl7KTc3+IgKxsjWVMuhBGOv+Bqvbfwf6or34dBGy+v6gpwc
HzF9XkXLZexNeqgXdTV7p3NyHPRWjl6Pv9bL/k+Gx3gVB422iEhedrcItz+WHujR
/vuGAwK8Gr/jVSPGW/DgzVcLF4N2bQGEeaI0KB4lqQHBUEMST6RmUSD0ncz5Feqf
LqDudcUZssCtgrsXtjsS/dphR/SKRZhE+lU967LqppuSq3fadyeHhmEbbWdgN0XW
Roxxd6ER8InBI6LgX2PDRQT/krXp2QA2KK8VWJoRwa/ft0MRw1vHhUSUD7f90YZl
uE+0EZUohkUlKBir6q6isjWAhD1qs6eAbY2xUMq83VLiKKAbBMXHUiLG37wfD0iu
J4vTL73wuoy+m8+VHM5aiqJkLx+7USGdeQaUK2w5GqTOJCyakgjubkC6EBI4GlLV
sv9LLsCQr83sFIiC9xH8haIEFXM81jhOiqPruoVNu+UxCdFJRsgrYNpie19yZJf0
c3cmAzIFt/BzN9AVxb4rygLG+yNfJSWsx4ycwv4/OD9j4Gb2NSztsG7oL6m+tWFP
xKQM9iQTdWb+WeT/mrkVavmRxZOu6Ni6e+sWZoipp0ZxESGRm2VUyyMpfIh9isRk
n+Df70hV3h8H1sizmyvd7X2rl5Oq4Yd/TMmmtmkTEXOr8Z7B5mGBdd1h9DPhh2Lf
vGSgeMcZ8ZxGs1xkAHDxvoPaQOahXsoJNG+fAi8pJsLZRQ6NHeIOuGtzc03hDRnt
Cqs2kMvi6T+mD2f6skGsZPOf1IdF8XIHAndIQbElLRCJ+kGEJcO8AsgTLLJvXrFq
z1fH8CMk9uyioS917esQ8DJbzWgg7bLhH28dX3hEUJcgetEY5/AGJ7SCxuWBGTOZ
KMVplCGLP+XHAMFip4zRS07lx7u595sdtpKxlmvSlgbDz3G9r2RzlVBR3R/30/ON
ugA7Ov8NpF1/bQsReCG4juokioqQc4iezn+ivFFVTa8yVfrUgVJjloNGeK3rgTw1
8XbIVwp/7DwA5gk0iVu+BoJMEogkRgtO9B2QO6+F89za8Yrlaf1S4u3dOw7iNPVA
q93KPmIPN7guyrISaJFkz58hXmqUbZeU9xLKd8+txSrXgpf2oMP9JxxmLDK6WXYl
4sLExpJJfgv57oXvvc1OVQE0KIa7gKjvQbW0A4zDFscoJgA7wPar3Z5wWoc5BqDe
yFMjlQ8LSH19EUitkQjuk2q7gpjtW/S2xMSrR4umi52ZGpVno/q/OiqdFyoJlZHa
py2VocS7JS9/QEmW1X3Qm0bbPMFCdIxe/KFoALT9b14+bp94Nrws+29J1znm2r+Z
+pEhNGAuPXCUGCBlaXDj08rumJ1s2sWp9SiQd1vOT73Rcg6oESOmAxwbbreCKZOl
0blxkOcLuwBAnVambpQLoTv7uRoicmWsb+iE5ec9KNuVB0wPx7R/BznoaIcVBxwK
lBfVm/AoW91UpO0cf52wA8QC6Kb3ydEO1dYUKMaaxZP+TH2xpofUY/0Qp5kDgIKA
nDh/ox1oULBc+rjtiH2X9zS4PWNpfhtbCLfEvpS+ECa9Nf41RglapdYT7QvZMDpk
L4v8VgBDGrdoE5jF9AnFP6dn/Hscb/XTbiNyVumVBTXKuMXlwB9C7smzwjcc9WA5
6QDZoNEdP3e6+/7H1oEwGGNmYOV4dwdrBjY8GTEMcqdlBD6WuIZl+x6PVwRwjRrf
IN0Wqc0sxo58rlx0Zm+B5LPzyFf1nbKveYcd/AvsL+i7x82ocu2qEiNpAZPG0sVc
0rAWIBuIn8ordfE+7hrWUnz7j37VQanUyv7ujvgQkNc1LYiCfKb/JWfMg6F+d+UX
FsMnW465tcOZ6mSF6MBWn6wbjAHp+UYREBi8+7e8fx5DBexJZ3H2sn7fO7hzoip0
CMeGHIPL+B1ICA7v4VxVfDRgR4fBzBuaLTNZo6gTzFy11NwesfgvzvLTVpTwJMGx
bITxr8tHCVtJSAWRv6DQM1QZ0fNjGihFGSXICTjdUYrLp/xjScfi4eSih7Sa0KGB
rFmyxb3QQpWVHLn80RzT5VI1IUnAy9lv9v74AIZz/77K9exMJX+x8PUuf0wYiGnW
GNAo/cv5lBCjByy8TQFX5guirUv1/RvY8V9mhtX1eWESfGC/1hTsYEYpQT1TNTb8
TEWgDro7qrS3bx6tdwtUNqE14u2IJZ2TRMqFlLcoU5NBcUFTVByQkkdw5UaXOL4a
3eU7Snk/0JJdUkbAE7sN0s6ogZnlYhTQRo5S8LY46NPJIYaRh7Fo8dg4JVSLKvGL
Z7vdwoxBOyNpCY34ljarX/ryvPb7uNJZw+Ms6mjHRQmJ+xdEo0UPYCGnserZT7ua
rEGXfySlOKtnlfxbkvD18sSPbewO6L+66bTy9RgcalO8n0b0twtvOsCbF3955zNQ
sETy+QGshkEFjberGLihSBbjOeB0ixQ+mlCttCJk0suiyE+mzSWh7WBHtHzO4Jfj
F1W6yLavnU5x1ubTrotd+2ydCshfwltkeoFWwdF7jyMEY5yCQycHmdude4YYfY/N
FJfsJMvereknOPXe+2zxt2PowPP+YR2qIqtAeIL3TUI3qnhy7jsZJi+hukx4NVJd
ZMZDDXosAiCE9/wZZga3yNpDuU9bkDcfU9W1izAOpaYAxlVpjBBENx9jGYfiFBLC
cnDR68bj8BOCnvwrTAnt1Lnloh5nbu0Y7I3kdbL0ZYQeHBd4ZkMqA2Ty9UwzasAH
Rzgmucajn4xFjLA83B2wFrImTEfzjrZ5GZwf+Nr8s7sxJPSmBwsmhbMav2EDkMVG
58vZbzlJ1MjScZHC04Ixh/5sJ/9IlsEEQgZ+zP+wpIwGHXaFVJH9alKfi1WYkdr/
B5S2EepYJRH9DPCl21fwREvgzC8kX7jzGHTM36gzRjWT8RkK2uNIhnEyCFFxwYqH
8O1SpJ4BfzQ8rW0QjWj2vhwFtEfeYarMcviq/9al3uJXdD9cJjwZQKCsYAL6D7Km
MSLlmxVJQXD+aN4KVL9Ta/oQrRHYwnjwbLr/mRMvGZ7Tut2/UNlCCtYSU1rYWy1E
QbQsT/0wslbxYu9lw2+hI0utu6gEaFXlRVGDFlHhRHvUwrnWlVdDU5BNpOma+10v
XBKGo8rBVW2irYGLakC48ZbSDERG1vpKma3rQ1zJhQy3KH/wCVeLufSkp/Wfkksc
o2tGtl8sBbYB8gX2ZTPhFkfkkgCD43iAoQ2MNOYZo/WTGEHpDifu/Vw4VB1Dwh+w
pCMKgTUWQmNwJuhSnG8IP3h2Lte1EXOx++UXxpGWnPMUVuxWaWKTdn+CYhbtT4bF
rp2nzgyeamlKmy7mgCsNEpQsg+bwztUw2z/D65p/uPAk0WDDfUp/+YZXk0RFTt+s
EKVWHr8fc2gDSXHs7QZTM6edahr5OVRsOkOWSGiBOiuMoIC+prJxlxNmc0GtKAlI
v6AIPHkq6yASwRwxbE3YFqXKGnytARdHsFHWQBvFISdg9aZV+3z7ClRc81QxhVHJ
CdSF00lodYnJT7Z+jDNHaqsnbPJJUKLduexFtY+scuaiU/kAZdeSvaTo/uvOv3Sw
iu52yE46p8iqCVDVIqvNOkRpaL42UmFaKVgeM2EQ+XDso63NhG8p1F2oRDOrBi45
UbYtDeIZv9emzC0LgX2hvMFIgo3zJolXm37vZthA3AuNpINseL0UvndCnS33ecQQ
BmDOLLHoHC/QKn9I3hQ8zlCSZsK5e5sXOprU1sYo+X3RyOLJkeCYDTB62PsjAI3a
4/iDc9/v58OKHleJqxi5we+3SAsDWuggnSnvAk7zuHMDISOods3PyyKor2jt0smi
4TLocSisanhliP4Ypt6AgNTyGketnQ7Ovd4RwgFz/j2ViX826+VKYTvEiX+k4zJA
IszJjK9C2A6K5FqwLtGt96stKibqiTk7I039vLmzB9eI2s2lT3w7nM5O4sEZFR/5
wBHzoY2Ichro4+Ci4KADg14H0ERPQxTzEp2L8v8SRfHuQSo01lcNYbXU7oCARews
r6WCcY7zqFHiURMGIv9ub5ZldtivB1MPzhk80THIGhgYCInrB77/+7GtV6Vuvs+R
6q7k8TYDXaLujdlC/DSjtSkgvUqOjRyZK8HYMiStVGPkd3/5DmI1aBVYSFm4jZ6x
1GrDMINs4X4TrgreGRfzUyHwLYpCrgAuLXKVsZOyh0fTKG+qB5g16efbnUx+pShn
SpZpiG9mLVCnqmfStJz/C++VVq31Ozxtl9XV/ctNEDb8WGyIT+kikyayZLRQPuZ0
r8NcuEPLOCOJlFfCaBAInusiYGuZ1I/IvWgWXPzX4m3su2E1rNrWFXHWdMRmkHhI
88BLnhEvNT9twBl5OSzzNzL+dXgpwbEN4vJdJn8miAb7VupDrSqBnlkuva7r9zAI
uTQAeuYU0uMv5jExhz2BbJl92ZxZzcNyaxgaBuztBoYuEOqCo3jxOlE/mAQlgbKJ
ucrjgwSZhd1TOPvKL46MMkHRsYKhJYSxhweGLBBJTMriBVybNpOrUwyL/uZANmFz
/WtbEnE0LNL6QejTfoh1V0lGSjbJ33a4jvFfQzrGMM0qWxX81MekWu4cOetdN1WG
3a7D0V+iOugq6T6kNEjzoGuprCL9ZgTk7dfL7ZJXKA1ZEgjN3Wf1Z/sjT30YMOCw
lvFe3e9dN2CtUbb7EDinhYFoPjyCofk/2SlMBcV9Ofg/W+aBMqN0m2AXV+fEJ0SC
sOezvAtd/Ujfg2p0Gz5AuLlLFyBOHTDmFRl8F6vEQlAI+X5pNxi+nFYRr1Q/p5NO
muRvI4UrYnMthX3v+xQo1YmcG7ArUVi95Zw1A4FojbZ+pitt/+e3MGqFk/4BzO79
I0ugwv46/lkmO0uCzudKvAAmHAFNopKgiiq5SPGM9rBBIMRdBr54oNfArNtRC5W/
8kQzRILL94KDLGqgxI9BeVRZhSMFDimEl8xS458s1m2tV79MLLb6LQg/FgkRxLLB
6pCCVvwn+sugPGA9dTY0h4pD51VMUZ3MKkCRpNpfevuEyixP5vWnci7liSoGy7D+
fsnvOnQILXaTEolzoOPGlbn+jAke3KXyxJrgTryCfdLWmdgk5R7lXGEeuJYzHyLF
srewwGrQRcQbOj1L6b/jc1OH6Ox4Yf51Xzx8an3cihTf5nljTM9sppcdupOR8t3c
VD8RSECVtjKWY0RJKq53+CIwG2RsuPV2hbBa/XRRI0sUxqx/l/cEMSvfyfce4UHt
Bt3/bLY3HV1IS2p6t1K9ytyz0LlRV2YrefbhTwPTfVF34zbpv8omq5Jh+PI5QjTg
hI0C8MIJqxbfWSVUd8g9PBsMxo89tU9RNPGxyf1jUH8rq/+KDbE7o9+dUEaw+m45
ZrPuVUR759NtitRwcdkmH3zsZDIRzaz0c2bspiKF8v+QiZ6T9HYkEoH+x/Egw1dS
qZ53b4wAw19RNHolSYiozGjx3B07RpXnsOzgBg/MqDziokYk/jDSEWZTVr7hcpPC
QzqcG1aFyNj899oQ4Du/OYpDROR4KQbFEn0JfgvgsogIe6gWpNGtgxMAS7GCZOMd
MiP0oDhJIqOL+1dxmad5UW5KGgZNp0UO7osglgAhcD4k83Jv9u2wzV1YDsCIH3Pe
3lxmPitPwnp4MfhMpcUymwYzkeZu1UXy/rHYLQ6/Bt2Jhv62cluqC8Qb8LcEzcOq
WMYT63yam0/Qi4Z4R4p1fMhjv2EQ7kxaxTuFmp9BAqzBsrIs25J5mTlBY6NFyyLY
vPssgLR6Fls+HonFUeLiXw9Wd+OBONEhP0DBkoKME60PPFd4KAwZYDlBtxL82FnZ
ajVlQAXd7AUa2O2pnvrpIXL8jxdkbJiYS43gWSpGBOtDvuwtXsy6UNY5SZrfiEVv
a/aTPUlZqfCUTjCN1KomYYRyyOgozhFFaHBLMcIlbC09lVyV5A3vbD3ZTNOHXnp+
X+9KrgTCVC9qGu8bvCheyiksT0/5xDPzoN5NYNezHV2Y4cqWRr0NCKS8vB5z8Cdo
weSL06NufsLo5wzDo4XQq7wCSvntnZoeZlLlc8Bv/Bl946wm37jmmbNAOALP3H6j
QTD/FTb+s00XJWwh5wFhNxrJ2vdcuusy0gt2iJKpgDwP/e1dU51M5X6e/H0Dfc2Q
CpA2mLPbYrTEs9A57fkJSoBQcOa/QErGKMYRSi/A4wL1Xe9aP8o9VtIBXBiDeSfN
yH/jlj1vFeS5XJKQm3jNj8iiIuFov3/mO/MjkfrRFE0UTdikTBFit1lLW5bm8bpD
B+mffYYJEPvBDL1vG9oRwKgQ3jL1opTaH3PkkZtervqUpLBayz49v9ozS4jWnhtk
wR3JYZgPoS+ov7MDC+VuO/4UYuF9m35VJBt7u73jPInnHT4WxGtuvnmLonZheqh9
YMe07gbTmWU254/Bh3qQvUYWZkMUbUF+hTfwQJe+TR1ks9c0SSrKsSi5q5SOSHr3
pclwwFTtwXJb9KawLxladIOpOmo0viSS6MNra1K60Ejz4Hcqdl3d+TFNPQEg4ALp
kFwjraagfoeuqR569xjfO2t5qy+pM4gbT0Ju6wVHHAefv1buxrVLiotdA7NBnjtu
imO/NHIRgi2wvCXFWM5D4ZOdc31K66cVLMM8YfxAjfxY0i9d5rnfR4AxKN8GYKUN
MV/pKaqx0FG0YyYj+L6azcvoiO0X8KGLatg/lIsMWV9ekQL+lPadeeX1htPeH8RO
fy37UBn/XhkNyIRpqDgDbVLdJbPi6b52CLMWu6eGtTKcwnFUgq3tcQfU1osbBEQR
rAn1jCqNaoeGlChZQolLzjG1OaZECY4Uu563+DTyCO13uBheq+QGT9dtb5PyJKt/
1j/jT4wY+3Zz5s0TenLQjlqDKkdGFy8kxcepTtBEr8KEyo/lhWkvh+V5xZjqQEkC
ELe2Noae9/EI9XdI/Tbk0Vdnru/Y3FQZP1M2FJBya3u+WHD7gbSnzXvXT1kqVfg3
qQZQytuP4BqH0y6+zrYXW00f+ix6Bn/Q2PsiZIrTh++9mRCn8XnzedMUuOjPrSw8
K/QVZRIuzpLQxqgIaYyFMN5liZRYzObhT4OM88Uw5VQ2uka1UCfynwQKfXvl4Bmt
sGkAQpf6y2q3+rmQz6UVKnRARGKe84MFoJicqZ9Lnwv5lqy9DgTAgXDlvzHmxluc
KmaJqPRnVRRO+nwy45VYxAHSi8QchalQbgpmDPGbBIhuzkaQIjVmfV5FWk7gGhDJ
qCX1tbkV5UuZ7U8Tu040LUNxq4B6rVUkLzP4zn3RwQbtvp+MpL/zpWwJVqKl2h8G
viQrj1ypPejW38bTkfKeEKeoOO/gvKR5+zy3BRDXmU/uaiCuz5kPnwO91Mkz03ES
Q6B0hp6ThAwhYpb+2Q1CUSimljyOEL2l4ntZD8g+7G0rj+KZ8g3zDc6xg56Pc5T5
YvZZotgEoUIXukykPUY5JPxJco5Vc48jrcLA5gL7uHzcoFjR5hxZBg1aVjK8BGW3
TdanTIFzD5J1gZ1G160IseRNLXruJ8lT5KNhtB7EBukzi4QWwyLANPk3yaUZzL9T
BBTaecsyxXElKBmVcAhwlIxq5cQxKiPGJsvKpG9K7spBdoO08DUgk+7aaTMneWEu
Kcr9eTO9bwsOHFqRgim+qoiTnz43OJknfZw7ZXIpMUeRjgDmxeQ1VqXzpJx8nVsf
nh+ZaRinIQVrv571M2p06xhvWxir0A/Kin9aS87QWQcq50OsJ0Y6OsN2OT/echKl
R39b8NrtL7ie9QLrNPU/2ZIBkkOcrO30IV6Xvq4EBS6OjHWqC3aSaEZY4hRU1E8a
Q4Gl4v6wpcAWqjj5nm7/ZO0wbOqA/p7k0iwcMNsKgmOw87cKSVBJ+M0Ol2lVqzEa
VzsSy/ciKJqDJ+LqLursRNT/98+tOl20SVMYloddObMYuBa9Uq7wzvSD6nFT3suc
PAsdkfC7B4LVNpqzQwCxIrSz7ld3T54VDAv0YunXWBjX/uHzF6E9qRMqJnBkPEkK
vpROsMNjMa8DXcmffSU2XrQiwqWQoL5W5gaQ9jiFl8PAYLNnnAS/m0Y8C9NBajWE
Ouu+s9uKh2Jk5lrp9HfTMLllYJ5NsJQuZPVYYn66RlxyoxdPacJR90tJDEIsE0Vk
gmE0Si5uRZQHTSfXzaxBfLdXJBQSYsAZP0iCQiiOwz+Szon1i7FCGZfBTQypvCe/
+VtBAqLoZLef3WICJ3d6wdAza34IsNfGmDcaSteXKaRx94+kcuvjUlFdly/q0C+0
JeZRMuJhVIP6VhyuZ2Wa13zVtsRfqj1z0wB6ysVddP/dKTlnMhcrLzpzsiTgEXS6
JCojXXmSBpC44GoreMpH2ulasriAPxCtYOkU17I7CBiph98IoYxsq4zXc1SZjGF5
gmmWVdVTTIgk38DcQFbUYVcDFZJCYYfR+njwIhXV0AssVQssfib7L7Mj35MoIoby
nISWwMzrLo+Tv5mSm9abCUix3Tud3ULxN/rdoqUDzL6+b+49TEEZb7D/Z/A1bTfy
+6a2i4ewP7LmtuBWHzFuE6P3waUORtczh6m04gyfoPH45TxfON2fFSfQ9R4qXc34
DjbMRXcqcLN0W4cnAhWj0DpJtAqu1VrYJMqOVHuS7U/7rCqSIcGAp0i0/nTMp6eC
OYb1LmF/rx/1+4Rwl0boBdPgxE7uesY106P6nFwfdhb8EXbj9mSQi7pdoiozHimz
Gnxuy34aIme5iINSUodnivaD2i5brTy4OLOdcziFr01/AqObX/ksL1xjK4Qt3Pfs
sNIbyqDw/pfFI9zmwp8AfTzIoNLGos4o1urCe1lJ+Jrk2KPJvn2Ru1aa4FMtPbWk
Fs99pxCGqFwVP99GkPSmWmdcnBF5oPFV034kcVe+/8nJxsOIa2ZVfcAcyFi2JZpA
g84IS8pVC5YrXtqw9l+I5SCOh7hJ8sDRRH0IUvLgeDVXvqqywrydLgjoXOl9obJl
OPuAJCBVnKxNvcf14O7Xw7/wHyCGJTYmzglVHXzDGuYqGGSrXooWDE7zRgQtKjM4
4Sbz1WnAl3Mk9CF+3s+azQakKzAr8lfSPZGbPtjWtiYNuHDl9JnhnOAZI9EMoF2K
7wRMXNWCkYvV4PcNa4MgUg2YIYEPh7yLJlbvm72e7leJ76tBnrIVOVugED7ucqc7
DMyFZMZ5lZQEoaKMJOio4ZEAQ+ABK/2FfzUhZ9yyYs+1jpasN0+czTu7PlE8ff1J
bqOhkQTtgz8KzC93tsdviU80GyLwzG4Z2V1sAH7n9NHl0A5EGe0sG5ZjhqdwXSJl
S3Lg9tvWaUYFRoYzcSkpUfJygGmIGdbrHeQAh/2hHhM1gjQCE7BU9kVfxx0X47il
XaP/fN6D9dSjn+LEM4yFVn74oUFC21JeC4LdfsQ0HPssUbhnadaRmAlcOuuf4XGi
fIiHTHRe6QfqsA/L8nqn+D6sPLULzLKrY7PS6yqhnmJMLc0PqMM+VX8evpuVV5Df
FoO5TmX6G8PKcgQVuLl9lxEYHxcOw3npFxGuTPM2Jui3kARqsVunIRM/m0JTSjy6
z1spO/vl5Wfs8dfvJgW6XW/MNaWbmc2EpJ3Z04VMSsTIYUYmU4Q8iGm+6yOHt9hf
mnnxAa2VI9sRnfkINEvBrTxXdb/dzrkI3JrmH6oN+Zne6oTXH82Pf3gV2eIkzQxC
aYUDtDq6WNGSATJDcsNDaAuzEWDwk6fFG8PR/LCeHGuODRCe3basGbKn79kWDzAW
r5EvFiJkM+DuqhaM1FJPUZxp0P96G8RryjxsvcKgIIbrtkfgaOciXZ6cWJRDxQ9C
6kFt42xNxr0BPEs2daveGIS1HHx9BTSYyAj/E4fhJqd4ftZS1Q/60gNaFsKd+7YK
YMR+5lLhb5S1ymkaaUxLWinbqEEnsuEbyJDvLNXzeZ8J5zRLZzwK3sqY3iyEh819
e6vrwW9SV5f5eDrYr8sS9wI+CEvVq1JPVJYPpXyKH0RxJXqUsvKGFB60GSeLxmMG
2g0YNPNyBflI2BG+OmdHrjlMVEAtMl9lei6z5PFGp8OxCkM/NX8zy4kE6Pmoih1A
wkUpDNp/ujCEGIj7jjRbu9r9c6CazEb60pr4kWnxxy7Dgl6ZMZn+mYKwowW1HLSS
rczWZvmkASXHw/ddXyOA8AJ4Qw5inaCg8R0mjfEs/LJ+cm3wrjnAmKTdhnVZ/UYZ
Z2xA2PqqTBTirakIFeTqsDqLkJ864FKBpJyK8dj70+sEVpm4cQFuJLY2utFjmFlk
E+TXsUr34buXfSSX+xZzvPgL34dv8ySOMXu4Zmev5b1nCXTN9p7x7Jp4g4MiIF7f
HbQFDqFolqQ7Y+twXug9KJgqIL/hOwAdgBg47OrQVFIU7VeBjJK5DTqUTD4PsI1m
lJJpw0ib5Wy/6oJCMEEvPZJu0pMLKupFh5tBId3b44k1i5IyflU+8n3f7iUK3gDP
/ZFAIvt7bAyVLJb+Ucxz7CoSHciN+PoPw1TEy3uZrZexil6ImIV3uvbbv/65sATJ
I+dmBKmsl6lPdjHpYiepvXHU/+J9UF3TtJtgqLWNwlUyKcs7CRhzFQAxnvTATIyz
MShJPA8BAhsA84jBddtiH/hkwhdJ1XZUhZotBiTs9F/EOubG8Dp3tgP9Vf55Aorf
BDebD6GIOWIkl+bZDKb1Ia7luOODEPn1vtrKw3juCatv8n7SSSsrI+BfPUN1Pbmu
M4p1XAyZZCenEbAT3/ZUYaGo09hnVSArA5X8AZHjUQt9ggHr1LzXdII717t0kK71
eP7ArH1OTh/e4ST35SdgcBTv92ZoCdiw4KmXFY5X6HpxVouvewWJyOCf4/ta1LT3
CnEm1UywAcEWvtuNlEBaNvY1db5OBL7eLb00sea7BsL18Qv9gYKPFSqHIF6SItkW
08xS9F9bAlLf8+n6RdttwVvN+f/mF7AXbjfKKMRqms2NGoX5w4g8HaqthuNfKMXf
E09yLlb8F3mCaw0gL0KFlWdrlEK8h6NcxuFROlffuiDhc080TtlkwE/GXoWu0vyF
9pc7Q3cZ6QgiIsN09xv0tbnlK1K34o174vMowRA2BziamaXUXgm2g4kNWXtr6Q84
5kY95pRlhn0S4JSTm9C2U54uhiLjC7SHZk+Q+GBTY0FB4LeysQbLbgH1usZHoBNl
8USWFObRgmqIt50EX5H/gB0Fy52CHyPjQDFUwGM16SNi7HL9mEnrSGPetq344YZ5
ptr/Acknho+fNFljC5lbgxBkecJ0AtJoHHvc1+VKLCERVHFm1+qxmPjthY2Hlt9J
eazFi+OzqDiTdbDSsji5MfZEO39r4YUNbP10nbz6bmM8epleoc/r881CNei7bMvY
FaTgXxZmH2gr2UZ7kl9w+/2CMJxY0VvHz7jaZpSxTh9MdNG+ys24LYQVSKHw+Yt2
BsYE1berNmFBQrLcZfmO5YTdNPBCZmlRM8pwILYU1KDv2kKxs1s+Q1tTIUe2bAXM
IwOvI3Fass5A0FE6uG2tZhntBIQrI9Tuwc6AZdP5P/3SFYDzG+JWB4mLMzoYuZYR
AxC8OdakQml/mP72igYXngH8JBLElTJWUwwm0gImmZY5uXPk21DmXX7abE47doIH
hj64Axg7gEDSmaZI+0LvNKzdnAma2f7kd3JGZs8OtBl8qsb5X5K86UKU+22vgoFd
BilCspmCxPzCKiKPfTHj97XY3p4uLZHBnhaLpkSpn73VxQAdeAL5LnmJSjN1Oiat
tNeaAmj7CKvEmVRwxG/AIhk9T61NOCEgq73iyDozlg4bK0Ix+4j1y6QoXmSIOQBW
ynde9n9KjSz9N8ybOkJ0jw5LHmWDxi8MVZEtWYsH7hElVqxrFgi5WAOynMDY5Tn6
PZP7mepCd8l4S8mQq0fEhX4l4wg8wsxJTHsAnnxxgYqbF9jks1xeYFzQT6ZkB0bB
NLM1YSwCBi1YvREumdnwqMP2HIEWAOxG2eo6GtRNTrCzL6wBaVvjuyzb3ll9YomY
vhWpxG5sE76e2PEocedXrzRoETk1EnIIEyOWeG2zaTsunoIvoJlFQ6Wxr+4ts0/j
THRISh1C78oYtyPqCObAH23u06xOuhsKdG26MFyfDl1mo8/8d35HViTFXU/87o8Y
irvgcfE7x8fZqU489BWYkDi6Bt2hgR3wUzdoRXp9bFy+k1y6p+pL54vutbDYzGoW
ZRnJk8JTbgOMVZn/dVJUOYMjn72Fne4N2xFFd8GiqWoRKusbC891QWygdz1VRJlz
1MkS6d1Zgky5HSAn/w2GpITUsFuZo9T2zlB85h5SPcvswyEFidjVs3hFy/acbUxo
F73LFzo1Wndxx0zkqhalNrvbraTbuOdgVjRLmwH6BJvhm37NjH8pwejqMwXgSMsO
aQsHgElTqUydlY0DgGCIiVCjbAoY6y6HC6aXg2Qp5rRvj7cIuvCsilA7d4YZkoGK
IEbJINBTMCsunNCg42KwIdND2ciGuQQ7ICnlPn0lLlXxJ1zrn4YeMqJLF/EnYVa0
LWPadJeWLkyD8mriJtP4aAp/6aR6AniDuxlX3auQhPupTe3fEsw9BnASOdDnmKX8
ndDRCGECLetoy1eNNkXi1s15j1TelD1h15RiA4q/VuHZLn+6iaK2G4dHAzjAiDg7
Ed7YKY4YPpq7fT9i8RCEi165+Q6oPd8df1FDLLYyE4Ok4UbBp+Ufb0RPJxnGNKoK
RmuHPxbE4i3WN6Z+7Xg5ZJ62oGjq0eYdhSZm8Ml8UfHwsuiPX7WN0/nBP20wuWd+
6wWkMjNfCWaUKKd3bHkAuqnUtOHlS8sJbd8TO0cx7Apm3gfZAcu/TN9ulM+8yh3m
PFezl2F2CEWizcbKjmqTXg4kWb7zZfBohRGcuzEsd6iVN8/gWoWRAX3OTTYaVu8o
cgaMTAmYjGDlyXhWCQPscNrFGNr0IfnHit0mly8ptARlWzg2kPcN6DQF637Mcqk2
5NhW/wp2XFRtzrY71MULGCPai4YD3YeSSc0xBdayAJLXzHadC0TB8eYs/cdTCGCB
DqhE/UdmooAeZupfWk+LzDLQqywFaLN9dIC6uuFD7fN4fGCaggC4fysQXy59rFxe
QJOrGH1WzjvuYlnsjNXUsTAlHoIG6DJVbFe/8DpVywSX+X+qk4qZ7MNGLlhVUXXp
bU7S1W/I12KybQg/XHJsVKVj01hTaLhHhyrxvJO5JJBreDVMSI9leTzs9dcFAzd+
+E6IAqvTs81BLnE5GrI6Sc1lL4Bqb9pNMl9qFkmlrUksaKMFuaWN1lAl5NAexU6m
5+K2UlU/fE8aGOoKXvWxK28e3Ie/qsSH8yS63u9wr3qnV22A0K4xckNt9QdvUen3
HfVDRDl3yQ3MjGX4fNwtXatbxOFj4PBJgGuX5IHUyiv6pI8+i+sPe9UKMPC/Z7Ot
JpBohtLG8lhqBCZT07UxpN6RaIVh9vo2mi8jDHCEmXb0rbRpaGWty0lotH04g1qB
/l4cLS4nDc/rnVNHXH/6ed9ue5WFIWRB+vf0HH84uoacRL8YJGY3WXC2krXThI7F
WDZ7EMgBa/Wp4pZuArmw8nAOEFfdBykn6sgGP8oJHmDefXvNNvUAgCaPb8JIH/Jv
+naK8gHenMcjYYpSBJEocrlkk31o84Fd0JlrQDOTCy00L73KWYmopwxkOZrNtCJS
5qxW+NG82hrDXTzBXdWrQ3/z7MekoF7ewduTsvjg0Me02BRrSyOmdBu91CfG7vYl
Dh3X2KwFCAY2HEGMXf0Z9gXWWRA1+BM6FFeTSWt4EPIc+bsGIdcMAYAK+k2s8jKd
U1ZoDC8zTWwqAMpYWP93aOMf/yaBc/Z4jaLoHV3gfaG2p5bVOyWStxgoPZFzD9uG
F2mYmpOER6QNtHbIgfXL+Aj1yWNG1+c6jHVWcBUkiVY0A6d0rgBAouC2VIevjkC4
hU7mMBnmFxi7o0+D+1nLshNA9mo3TFXEsQ1XHypkD6RPJYjD8n5ZxCaCcjpLK680
uDeZp7TnqeEl7th2/o64p2Cs3OtWgX0I22LnSiapwwZo+PgBhRQfUNIfDPguP1xz
EfQhWeFHp+Dt6jzC4rqKyG0zxTrlCBtPB88pKcCxgDI=
`protect END_PROTECTED
