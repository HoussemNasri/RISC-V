`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6cB0De571IVcETaoDDbNSsRb767h0geASwXWyTUnHpskYvt0apYrQa5QXN6jYbj
3uFrwPjfLEbm1o8Cd4nPIUTLmLhygkOxKllAXpBi69BuakUD0T2065IKUO4TKYoW
jR9P/8XWXWi60qy4cSKsBxz5VL4hLIKKp3SMuo4iHpXymizv92NyPcMcGRzWJjkX
BsIPUKXvWKFbgMrN7Ps+APJcSF97W7KikPoHPC+bhMa8pY0WTaJ8dlBpICJmOW9g
Ztt6Xac1ADizH+WeHFa3snfFxp8EhxBy80wR6DPgurOfXac0Mhv73ZAHbqKvp7Rr
9pVBjWbNZLyhzP9M9Ef5Kf8nhJd45cja3OqkZiqhqpzEzAhe+njt8YfU3jsKQ/tQ
rmx7/JJ3uT4pLAX3uqfvGKDOG/EMo/XUEMgnVPf6ZeKEEKStF2rMftsQWM6ma3ot
9aAuE4WdTN2X6L4UkDUaNOUqrkvzEKwwqDXvfd5j2fXvN1g4pJdlT2OtB9y9mu8D
Rkw37vPlh1dL0B/BZHNfU5npHRndaFEYbNCuBO/JhDNf6PsDPXKxbhpcKPDG7Q4d
7fWS70WwgfP15TkyZ9HSwAPdkdHZ3vGexqWdsVyjBqMDKUzWBcO01f+87SBpXIMA
aftY8yv+uUegra9xDBWYpTBGhzPZNYXTfhaMeQaiwNgwx5KvYqM08f5gRSl4N/kH
aCqamyB1vx4Yk5pgs4HdshfNTw0tqw+Sfd3XLvvLjHVaF80yTTFar+OqtIBNkA+S
7eDOfNwqpONevePs3YzgJqWYi7E5OOD9cUIzDq5QfX7W8DUgxAqbrEeCOxDrwIjb
vQARI6zPN1zAhcGa0BTQxl+eNgnx5TKCU22vNii5ZSJPLTJMCWVM92K4jbKQrONz
G+/9PsiUaXS1ybzkMeidaq7nz/4i9fDu1HTeEVNBVglLj6CLv6zLdCYaSWQlZvAo
i39iCQh1n3Mb3IL2W7z9DDeOXV/4yvjLGF/Px+oRt6dlyQ2uTR89/mh6Eebztbzp
0pQsZG7rSTjD702R4+vO49C5THiUbOw2wRPsWtnetyxUlgW8AXl5MXpHwWW+hYHQ
/EMxcNLRCrV2PeSTy/DnkA/4WelhfVuRlnsuWG/6ulthSUZcVGRD5f2SBt0UXVZq
P0BSRmj5ENcnJbTub8aDdTV330S+ulCaEK6b9WVvDudqUrp5clU9mTokYjoYQPRh
kKWYtP1iMOmdc32QHhC66EYw4lkj/pHWSpZQme6RAc7iPhQz4VByi3UBORDci0Af
2qUYSQBgL8f9n2hTCLLKpe0GJOkurL2/hQCH1mTs1qM04G4sBJdLTV+p++yLh1Q7
7QswyAzQBgslIUgMcouZQIfAKYDf7ndP+UpA66CMaUs1iqey1Iasvmn/wWBQIMJ4
x2UziDmqYJYnEHzSZuq5OuULg6dUMjh7eTt6YJ6AP7Qh4BXm+vidvSPmjQeEYv+H
ixaKSd+8MnsfdtjtZkdPpU8qXXUi3yUy464L84QsJTF3d1w3GA9mRkQwcoVZrtWu
/sbXW9tDhd3+ERliIEMOQIDQA+9813Cbj0ihsn086aCo1cbhSkLmp8eKRVUgjNLs
eC1wpv5gDg0IRLuNwsxVrP0OUYjW+6qpDBxnDCFDApzOBVe9ANCSAu/TvKJ4Pdf2
Ds5bH1ejGjqmoQCDdF2/F8RS1+9lySPiw2TXZvxbmgK/dJkN3X70YQFSXqeFcHzm
8AOYB3dnCtcRAvP/TZiFuC0lsHJROW6EuhFH1rIMK9G4PODRjfWA/ipZBaUS4fEj
`protect END_PROTECTED
