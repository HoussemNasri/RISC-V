`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N/auRas734GZ/I2JpGW4BY4B9Wvqvwo6+3CluxnuLYJsyl52uzBnYZ8g9YDTJ9W+
sy/OAu8FnxPFDQ83ze0ptlrwKw9n3123Pbp470yn0vDJtEpzSe0JqeWbsBKsD0dP
sDHSAPcS9JdHj61x2oScqkN1WAdHGTEJXcXX1xABrJKO1feBYVecsYnmtJGUpscj
6tlZIw65bHA7jATXxC74mQPdm3HXhly5j0l4azZX6qdBfsnum2k0Yxs2bGZzYxu5
3LRS8YcbucSD/gqw64pZ2NsTme+M+N+r5uOvH0F+HlHub/wOVl6zQ7wTQeZa1sQx
fQMpfPISNWUVcjZ3Z2EIJTlXbRRrXQ6qMKL7C4EJbjFSG94zG3l9YPYIscn30cju
b+BvOv3+vkoNv+38+YHmjzv0+tJioT0MAZLkcKNGpgYAbTIJgfScX4Xzr7M+STiI
YI1Ho3SBb9PVuRJx4UxfgbywFORN9rwq8CC0O+r56rhwWCOyKrts+YWp3WWVce5q
xhK0mxeiNN79lJs3XqLuYFo/DJnGFrxGK/GXdt5hu2R7uwSkHCepElr4tPdOPKHw
OpRwo345A6qyw4Rqe6i3d2ZcgFKa4QlAsd6QtPGT+Y7z+TSlNgOoOYDTcMwJqbIc
Y4yhKG1y6K6qxHLk5XXivJj3qxO8cn9d+AibKZ3osKGGBvc4O9a6457R3TFaxzCt
zm56bItBMRg4Y3NMAHvTDZCrF/RS4NgkYcaiF2+n3TfopCmKs8fUyjC8DW38ock/
ysSl2859tO6kq6oovvh/xZyjHuIryFvffaR8o6UlTwJjZbt5OxxyR1uj3h33qqhk
6ooxF9J8DyxpBJVMSacnqOHbK9baUyLFVhtnhyX5OkOF3YdwtSt5Ymj8Ez/Z5yci
Gs86fBfmK4ldKHbM8yaH+yrex76zVquY84DlqnJNjAFdYtVKFw3p+DvW1+ZjTNVD
vqgbnCb/E0GIzHIRkgWqsk7GUspjl1zC3BjZeP7y0d/NQ6PendUnmRcLnOz25dpa
vhyRCWFPWEB3kXsKVHy4I2jj6B542x0lLTIOr42cY2zral1BLFk4jDPdTy7t/CZr
8GT69QMU0y6z5z2aGGDxuCuA90DnpsxN7p39F9SoeGRd6mBoKpzCoSaMaHstQ2r6
Itx0zZOvE5cOhwsqjWlkzuidWDES26N8AZnEdTQ+4ph8UoGy1LE+qMl/8gFx9Rsq
kw1oO4aGIpRFG2hb7GOQcXKc/902gh0+WDCsRl7lShfnT8q/z6N7GHyi1OujufGD
WAqnP4H0pAY4rgt0+yV7/voQ3tP4furEcXSkyZh3IqSFdDAPVTycN3PqAzGtwEiK
W3Gcjzhtd0go48rRvYtgrZrorEchDBQGkV0Saxn5a/dNPZaA4rzAwOCN43peP/ki
cN5sYaWyjuGCaI/XD0yHXtzTvpLEjO97WvC3QNCjITLBruwuOY5ed7VkKqg/xBN1
whXe7xNsqBDqJnksiP7yE9HbXYg5rRTYnAQyhl2HPTP/zka2jAlq+kly0kCymZiw
q3YcQcDzdOmgAaZpL8vx8ER4ZrAVcKOQpBJg/Zn4VGCifpu2H2LYtX+t2Yl2sFvH
l+JVVkbV4sVbe71D+EoOvjeFjuXg9zaun/wtibo0qn114YOl2PM/6bLvYK/J529J
tbmYPgfpxM4WkATX+Woma6Hows+ixUKteDnDfkR0Mqo+K8TALSP2Y6ecqVgfgY0a
EWR5sYKuei0dfNuS9tHL/JAfDIwKLrBdslUu/allkZj0reiMVa06Un8LH7qTmYG5
oawKJBJd5CwZjOC7jNVLY22IHRogMI9qN04NJwxleovbmNvV4ufiLiZDLpvY6lNy
OwD+p7PszNOIYpZxnKsnx30b4ou0QAN4p/jTNvR8CJdQpeEzTRvkIf6grE+WS1m1
ropILmpzAUc4s9XkxBUn6xX2hH4VQq4f/IYQsPeT+6jpFrmnE5NtR5uKiEAYTCcC
KI/4BVMvTMlSZVHwPETd9MGFslSTTVwIPt7ghq7dxQbbm4/qov0rIVBKwfr4vOSl
TeTs4eeYqHtS2V/mgZ8gUYAx2PYjq7wWv/PB4k//HFUAKMVZ07+PDC6Y2B8Q2U8o
GmSIBVl9JAKwOu5AYfsziFU8Tzz7OkJrPz2M/ijPftuVgeqhwevmjqilIHFdREQi
PvG1vYYTxvbdK3fa+y599v1cjilT0NSzqXDVfzp7GLHzw3p49ZcSNM+jhErJnrX7
Xvu8cVc2pw5X2IHl5IW2XhkHLpUam4tXSGJmITYk9BKla73H+1tWEo4OtPZhGAk9
ot5GZbewRiinRfCetnoqChpAKL5VorKofGrOuYZ8vI5FfcXqFzEyJUf8aYwCfdzM
ZcHQI/cJF+p4qinF/sey2LXOdQn4smnxumJVRUuf7cN0PwoRe+BcWeYvw9y0XZqo
M6DkabwWMA69nEYARfnTjJ1fW6vU9xMAGxiNs7gis9hZB4wKDcekvIIXdxEy77ug
LJmMXuvpxYIOYPiskfSqPnw8aZSHuts08KmDZRFrxaKasbNOxIowwHzUqhedueFO
KQq8XuJwPgKIbIDeWQchS8NnJaKktGY809qktsfzkytQLUJIz6JEFOfWfE4NqmpM
RLDKSwg22wE8uUlH0X5tIu4/nsNnb+MyA1QKRXMbAV4NF+96Elr83FekatNdoXZd
sdmtX0Dh5yrsaPFv7Ov9TB4BF5ZC4g62r6N6g/3JQa7vwd8gas+NFWfrA3eISlAT
YmMX7R/sFqzXmF5y/mZn0v7WzUC+QJ3HQXNYnW8H5UM/NJ9uSEimYZUCjCHSlsjT
snyd7Cbv3K7Pn5CYwCUfFnAhRZlvBts/jS7pPpU1zaSoO28RJEwcaQCJoPjAVnJT
fGPdeB6jQEp50cJRAb44gZU3QEwTzh3Z8xxR/O2cIx5axoHf0dQhK1uoXI35ET6U
imj+Jr8S/5+/2CcSpOD986biZ8zQqpNoXXJ4OATVZ17kboAXMI98LI1VHfpo0ze3
bXZviUZM7WNzjmIcZ17DiRsb7qjUtGocdKtkbiWousLOoRyPb6aFe7IbeEjAXE7P
E3larbH2TC8Ynwu0fe0ZAx69NH9GozaHIsUIaMEcEzeS/JDAUonR90jfeBNOc+Pt
ireEBWOVVvQBsKpiseiaqUdBQ/65k6sd5/HY7YcmIUukuTltDvThriO0f0hb1yUg
L333a0FK3/Ojy1tde29NZhrp69WKwltDwprhlU2E2Nb2ZihP2o5pV0HdO84YqD4T
8qYu3jlt2nv6kjM0dCq6w6N+4PkR0X971tXSO10VDEL3dOOH8rIbq81GjMaySNbH
owKyfwLC42YAsPg7XfeFXeytdnOA9WH0AEg3jHM0DT89xBUWoc51OTgQbirC/U+R
5xS1Ua9d/utKVrVyBRI1h+tUz9EVJuERCLYOZUFfrXj+eEufZXJFvAoaRx6fh/LR
JPEoy1phGniFyDBVX55+Ot04mElOz3Vxk/8vEStpjoZ7UCo5Z7jwhRwQTa+iwmgt
fhbNsuY5FPX7P2WtcU/KSDLoVfE9HcjLmYk/fIhajvbHWOPv7QI09rxqyMSb73VG
u6cCc5ZNHtMsBh/zKjZvWTsgEVCArSF68tAStbfssif4fOb1dlRDPXpikV4QXuxn
9N/dhPoNqTsgzUpP2aiFt6312WHcMR7dixwgj9qWxxLgwjkIhBngLQ2a1FSZLTsr
63PKRpdd//ta3J62g8Y+pO1VwtKpGJ+qsspCfKdytnSV/yRN1v5ChyojG53/oc5h
enKOTwHrK5hM/dG3EqHrlY1tfYbbl27CB14P1Nx5OUkNilOmC3xnw12eJlPXRsYV
P1YvfJs8xOsZWPSaavgUqIaENU0CBU2Q+54k+OPjT/f1WLpDZJkDaHFtbbx4XAal
Snn8iqljWPBSM+lYV/JKoZJKbdmMcWaFqO0Txc0J/TVtgYnZd1tionul/o4qCTwI
Su6iIjxeNhP+jOHuN07MiBe8HgALCKqFnBIeEt1hXPzvaq4CTkOBE9U5Loxghh3U
nlJmTzYSg3QStrA99OtFyLig3A7GWvxdxLjcgfIdgLTFFR7l1+PNMUJP8F9ffnl9
TwJ7oQvKejIt/E37EAo0DV+c1csdD8IybH41nQ9535qttZFnsnUhW/xJNHFN9cw+
steVuP8oFbycWGRIRc3VOjRrAocwNpgwcgl2OpqyWTzlRidoS31l1qN82sv5g1iu
xK1Ho2h24Zv/fmizSqyGFgKISL9UtdQneQS3dGiNtt8fL1XyqtniQ1yaWA+6Ngbc
mLZQfe9k/TgdppLC50UCRBnH7xIH0PVH7FBZgqYvLRMFqsdYBM7deRg/D2Hd5g/M
+ftpjuSn/+Vzdessb2rZesyWNETv5cWXOmdnHrA5tFU+5RU7DKyRJ2i1HWoPWegP
V76BzTzVvv+OPn9sZIQFV0gOwr6mJ7kaKiodsFYN6RG5tW17DDQVQRa/IKptg//Z
j4D5KsMDPAr7cZZTiQMaWgoCcUsryzTWbD6PzNGsBAe3sPcpekgJeU+7xsV77oys
fsmzIptX79Eqjw2gmjbOpJNQp3XM5TylL1KSbA1mtYpZyPMoQPpy/k5rV1jAfeyY
XcczelK0Cr2vw9c0odq+FpkI1KGmx06r2Y6iz61kslcqMysE6v/1rvQt0M/0iX9Y
EhUAvfDS363TynJIGqOzC4bK2pdGIPgTSFror6GHEJKO3gU4pM7TywMrl7tSK7OA
vKa9WcmwNntNrIY7kyfdzzCVTNe7l00WLxU4yQaVuIBl+xvQIhP7JjdbPbdghprs
rY+x7ou/uvuBHI6iEOHzPtVmRAsA6P4+oGhY77GTNp6+oqZTVgks/0Zzw1/RORM9
VyscgwPgNdbFiIKSY0qRcDJHPXJyBVYWD8l6Ay5naNersrN06nKEY4lnqumMVv03
z5aKHZ6c9wVZbzShA8xysLRe1tnepfFjY66oBkABOIxna9psolZPU6uJrmeDrV3l
7yM7aDzdt8c6wCfFaAndeAzpvDtNSjOLqOjCujvl2zopueNfiGvtV4bU19rrlKNl
h5RPbvQFvqoRYUeJ4CXdmXoMNXI4wDq2IZ3HZFx0xrs0m0mtkwtEv05RmjAU8tNd
Tkj5BeNMfMeLVp9x1NZ3XcwW8sKfk4aw0+xtL94B8RfvJn0Li50LVBjsmGehecKs
J20o6nASBtTaIi8Yo6/WDHrQU9JQrhxc6F2ngzFTTBdHvwH/wCTjd18KGp7Tfi5H
dYCxVF1QHunnDNKA9bn3VXaWHHVcdMk4Z/vDBYGScyo6uWTuG42Z/7mZNznnIRaT
Wi/j2LD4PVF0oSXHyin+h6Gc8VKZVABOyix3ZCjYUsivJgJoxLZhpVDs7OCMlRiU
LbLudlY4TaQaD4crqqvBMMMR8RtNtu5mLmDvVjYtdLzjsfh3A1hPbgbJo/JbrDef
qGD2ldglJ6AuYXUExkw4IxAjgNfdnXitMMa2PcMEk+NK2fADcaReB1bdh/sDFwft
jkRW9WbrdTGhCQ+3cleGGG8S4VcMEBZrKUrOVoVSOh3RK8e5QbfdRqZ2HXwIP7bR
1saxUeSjgeUgYdeP2unyIGCmoD/i8B4mmgBrhZ9ow9JztzcWb/pE1UrVcdIroij0
uERzeDUy8QqIydiT9SdZAA==
`protect END_PROTECTED
