`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZpqiEv144RLKvCkvY5ofQc1fQnTanRePBlJ8/m9O8vppWTz+fCLumMvaT+pgYxLX
PZb4x1WFskel6NeEEpo0OsoUTBF513BNL2oZYLuHlBCMpKpq0LKbZLsKtqaipTXp
WQtKk+VW4vjgu2t1sDtKpwKWlDrTiFTw1c7qfpbJhHb/vIprRoBpXVScLBHsqMbR
SeFSsOh+ZJmK7Dx1bYhY/Tx9QoPWVzjDwua3JgwfsxCAfRLYjDr5ESdOgMhBSM3s
J3rwASgW7FbUIm+oE0UKWkK6kVnat+j74+fNlA2f3OH9HvZvibb6RDOE8ZMIvu2R
eNnaP8QTZ7VWfd2GG//XoHMdSH5rIldpuHLtYFDnymllbMhSkSd2npowCg9inLri
o2BOOLtL5JiMfchfR58CdSXFsPxXeC4VXFWSL/iJCRcBp/+WpJBU+0yRruDGSuMW
KSCeqVlyUU5fQVf3H55b5qPwxIgYsVz4IQI6qTef2eofrpvBurYdZ+UQ0uY3G4ql
luGVwz9Z8WpQQKQThUlPh27ftrQ2F0zn5wcCZyNalrxc38iobbMHufda1JUVc3sI
atb4PVm9oNEkaD7Sxnaer1wAOH7Wp8ol5lzAAC1Xqwwd5H2Cw1aPZSSjwwVEFm3e
VYV9g3b5aj+4yYL0oM968DScWTSymw27UHxAh5v3C6RepsRGChlRn0+D+cu37EsJ
JLHIbEfq0KIFSlQdjeSj39RXqfqMqdWPE7XFQPrqOvLCixkQ94NLEiOefW4/7qFs
4ZvBMcSAoHWzfkavzoadZOiFuppIUOAg4PyoOM7flfkXQtHpGYWSXkXy60XTHEV2
tw83cJ11UolIF42Uv3tFtkX+0Ec7kmEx8f5MmZfQHaJAXGmpOWG3K00Pgw9UrJTq
JKkUJ7wXYBYnk7eksP/el6J3v0kPGJDuZiGlqTgSBDRnK1oVj6AxI2txXF6ECqQZ
dmHFUcp3K7Ib+56tQWsifyCJWDFlDpV9oMw+2+WWtItd79oRjHGA8GQvcW7uav8v
FztNeWiWmB7SccHSgpzbA+qql550GBSkAu7vr+ilKInIlehshaQqE2bFjSpWwV+c
aotF5Ny/ONkbvr0PPRhreUvS9gaAx9mgAviybmPOgy8LQTEo471jnsQMW2JWGrpo
kdxcS3iqawXkoNY3iVbyhTqf1Wp/VtPgixFk44GGFXpo284+kkTRfveZpVs3pfNv
sCCFKfTVqqRbHUNUneV2dNv9UPyFk3L96HGNcxHSb2avuNT0P70MsoFYnWenQV7s
`protect END_PROTECTED
