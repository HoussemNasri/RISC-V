`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HPTXWY5sLhCy9Av1Oo4yHSRNQpASPNP9RCOIWpIwZ4yRCQrNcroDZXoNQb2e2F1I
KuuG+Npm8ahgUEkrKuMqa5+iMdmH780cA0hmJeh+495nWifqLhXI8EoD+dvN8GPN
yX0RqQdeOtSoM+vMaetQ/JBHoYVF87+FDpoKrIwwkTfaH5p8EhgAthHX7DFqREFQ
`protect END_PROTECTED
