`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lv2YOC2CFAVed57AQOwRtx1aROJT39Q343SB5KfrU5PbnSRqTGbamk7+i/o8eFeF
9E7MMhxXFXEtoD3GwJfIGlJBtdEdHnh77snKaQDU6c/L9zeKm4V+ewYWno8cbMfQ
2B4+V2UYa5hU4ctDThFe1LdakSJoGP0p8spvZ1CJrDSekcWnmQhjf5GNseQcioiJ
h0OdPXVft/J6seb1Rtin97G3daE0sFAm0m+OWaCVpgvLV914EOQmj5aWB+sAf3l+
wgFK7j0oGhnXVftzTIOHna12Azet+UJwJw62ytkeaPdW9aQtX2g9bdRJc7TYDhNU
OFsk4qOEDkpeUkb7kOv/qVD8IcgXqNVztpDM1rMPRFHCIE0r0HLQRhi8yLXhAP+s
gtZx/6juY6JhnJxuK+WiLNRoHbY8hnSpnVza1MTO4JgUo/RLmBotrwmUefp72sat
J/aW1jvTyaGLza3j2OjBuq1ZAWfj/2j/Lr2IuMiygeW/gr3jRcjCX5g2JJ8NAtYW
XJ78G86zLAwbcCLr17jIjbZWUFexqXLvOczWWgxwjEezpqnfopvXUD/syAtJgJti
G0fgaoB+8GBRiwI/ej/qkV9ulDAugePIxZaBjMr8vemJnhEN9FbLVcuIq+kCv7bG
CEw++etvlmMWy/xoSOD6RsHqjsd3icR5U0+HtFWy8Mi3rSS9N1T7kdwzYkjQFCRH
Mq1BZvEUUJ9JDDVr5WIeFYViP45083R40a7/SbyfahlvMv+OsVAL+JnNYjcZG3U+
qbV8FW4IUPYzdiYZWgyApNEtbkBqNpKIeJVXPRiP5c30A5IpouxrVQtqvJRaDNwn
YdFcxSUN5FGaf348FwRd+B5E8YHzNUz3sN3bcoHP36HYZ5ppY/XjwDHuouF/hjkn
0DSaS8YCed4yzV9kQN07ewpmYwRrTSVnEp16YoxoAJE1zyedBD1eKg5dzr5ZMkTw
0rdXRXe32d52EMMifOxwgNuoLAZSLu5r7vYXWERiqJmgfL14bb6ViP6LnaA0DVLg
y71gjbJ2p+0ewVT9HYhlmEGR4e1HBHAUa7sCAZQ7uWuQyO458cYR7eVSabizQu7H
PhGdjNZDb3H8psdZOv27JW70Qf+APwvPtm4lENk74xrXdD4dS8PRnQIXBkF+8a00
WSqR/2bLx5YV8rvUGPN3BSKi1QWn5fbjD4M3poFBBfw3IJtP62z3Xj51UY+HjxSS
y3LIvYCO1YwUC66sXkngEho0MGpic4yj20tw18PQQBlJy6pL2utI1frdgwAYS7kF
sLkUh1zCVNeA6xkXMc+/zvhfDiXgTfDfg1u/82vyL3EYmeIZP1HF3yjYxdJsS4kD
0pqAfp7R6lOAzGZrMfy6AOtAJAe/uqyKxIbDdIAjDt6DZAwQb6AyyFKhe1ZUxKTj
OA1a6WeMqhvevZ4QwBQGnCo6PzOHv9g71XV873R/I+OTItW6jYqIlHAFNfdGKvbf
Tz/UYo21WJ8o3hZFjMzUmsuGa7QChh0Nyl6EZZCcm+JsiX6Tfa8BTuFUoMowVn9Y
PVjEEV+Qv499ewEvvf+9GwOKJ29RiCLuYMzIPzBIK0xKPg+F5rbQ/mc83yAnSuDf
FCz7AY4qtPZawe157+pe53mbubu2IsZSKxKNFrxp1AD1snnmxQbPrFfzYT9Dhrg6
+AgUuKIQob8hvUmnGrjvDEM6g5JjngYUUBUqDSt6RFlrbodD8ChLYU6KO0Fpr52R
MlH8DdV6da+eWJMXip3TPRb+rODgRVXoCSUni/1+REfOrDP+k8FNaoU+CxT44OmG
cUOhZwaLfk0pjrn4IT3AK/oTmQbETjojd5p4SL7a0ftJHShyG09r1RyoCOdO50GT
P7xJ09VSYfWaneh/WLvnTEyoAD7NHe3Vn4LSpHHPlGwLsNbanuqGEXtcvMfQi0G0
O1lfKcCOcwcSyHUrS/2HIQ6b5gG3crPItuYIIaY1MRefVJ76DQru842/FTDzdHgU
Q6xiHCzoMfMNwhkwFQkKYObnI9SoyzdvY1ZkgjWAS3qKq9B5OnYjCsf/DS7vbneT
1jtruxLr60jjJhnz22ToJ2rqOUQ7ePlH7Q5zHjw/cp6amaUsIBxDcMHze2s2l2Yz
EF5XYIGQZINvTWyAyMFEeawwxvoJz8ErsedSuQWaEhEpWM2WrI7Pc7dc35cfr9U8
qHwsN21U6XTu70zrTkocMpCUO9tgPVfdOvst0ogE+svS0iQ8cFlBTEOUjE7JYQaI
qKbTum+BaMH3YtpH2yJkFce69WTfYE0gyqDolcUTdnSMC8gaZI9M98+/mA1EZ5Q/
/jMPHfKXSsfaZJhAKvcH3p0wy9R0ikdgfCudJltnilX42y96Ym41V5x1nRHYlyQU
TDQ3oHxTKv3zi0Kvo1Sd2+dxjbdwL3X3SWBO4tmSnYf4FnzbBbMQbpQbbav1srz0
NGrPXsVWiZQzDyQvWPPIYPJpY6ryV31mKBSwVNxxWSzajWOKzoyoxHSq4KiQZFr1
oU1wcBlQ57+TqgEfc0yAAgnFUNIkwfC7zhtQs24UHrpJfpOcuxJ1tk7w30QSj5uv
het8TH+UVrhw3SayB+uQPPd/HCKiUSVuKA7Motkkmb6coLzQoStaEd1/uljxGZUm
JBLI92kHile3piz/5V3UWIN6lFQo6A0/7wM0Zck+0rGtHPz+Iv/Ho80W5iSKfx4j
U9NQuozqVGTnKAizgd4O+Iew925uLfkj4a9v4Q1OE75gxH72abBr7+yjQXAOVIFv
Fafg1Etqa4bpkV+DM1mLz9tJlOU4ZKVOezLcdgyf+1qKpuicui1N1jAHk/MF7Rya
UbFCAfZqKYuHbANyaE+9mkKBzDzPDWxF2OI7FRzMT5a7PKTOCwNPaGqRAUC5Iwdb
boaDikYK1eseOpcjZSE/jLZJI913z1xLSlKmtby1pxE=
`protect END_PROTECTED
