`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRJJ6q94TRBzfLzTC9wZyWyToKoLFi8yDSssHOr+lRLRsmPIoROunXBTjwd1YFJy
g9Te2DQWvEJPPYRAYIAGtDq4EF+CAOSNRBuwTERYruWf77iZFrnp6tkY/mOCZKom
FFzzoMlkmRGb4VPIf8298vp4YlQXNqsJfcDGZo5wSIfT0unrYzEMIqqXG5XAXSb/
gREsVVA7531MBm8KxK0fgmYH7iORSWHf5culDr9EO7MJJc5xu5T3b73Mrxid+0/H
mFpicFq/U+DXQSG5n5E7GLVCrZT/uy2S/1OiLMWZhSP1xVxq0d4HS3+ymF/iuZPX
/lzngBFEFoCJj1X7RORv5IMHMuZHJhzcCWpAsfW2IzskSsRVvvVWdnI8A/tSByym
c8HaedT9rj1S4EmF0AeQcB8n+I+RezOw7u8AboO3/gfpTPk0vxv4MouC75JW77ru
vidP1xdJtPmuJt+H8YAgQ/LoYaq0rPTHT92BgJfWhjCRdPw1hxHIZMinc8Y26qGT
u0Z3s/ugD09guyjPuzMkz5vvwIrCSm4mwZR0a6XIgnBSmhnn1YbxFpzIGtvDkTN4
h8qLvN8OaKitNd8x5FWWR0KgShWIHm64WnUsebydND6EbtjgIIdIFu125TEl+I9Z
WM+aoQ+ZbLn2OGrHsTM1TwyESYrcyx+l7LGzeRfBPwzL4XKcbm7v24e+AX9MvRfx
SF+Ck4FsWavsBRrxVvHRYldjJ0j3rSHb723qriUhOlGmln8HQuIoSdmCTTANEzco
fq1lYBpYbADHBxpbzANv+LMZvrhjKXLafqemZpRjKjn7ssREMHEqLNN3dDu3LCO8
`protect END_PROTECTED
