`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tF0HMmA0knfUf26BmjzGwkdUM7c2hZc/GVjSxW5O+hQEHi+AVatnLrQ5VA8Wk6+
af+bkn/zkQ4m8vi7sapdE2gMkqa0CgRZCvTmiQQzZJsAnedBQPEyCqUZA0U+b8Dd
CfWgjOXPKiZziQsFnK0gMWr8V+fSKETmmrR8PwtSMm4=
`protect END_PROTECTED
