`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hzVebp6BW+BS/MmNlFxmmwLrVIpaE02usjVF0aXgubMFoMdkKVz0S+d7svpdCOf0
RsNUsBrQ2VNeTMmIV2zVATBmBROdc258fEvDf3uwM3JfmGTwiX+bA4eRwpr/ymhp
XJUGW/V0WOqfiiZHnVL7jsQNhTo+AiUfg4ed+4btCjLD7jsTmq6NuE6iaY4xC42f
Ag0lmqxXdP3DMOy2mTvhK9UL/7eEwfH5sV6UcvO7fHZMWHQkOf7okFAkctAYM7rb
0rFE5ChzLTyJdc3l6P9z9yEUUrAjIv/Pb3pPvg8cCD6YkoQ8OOgT1PacpGuBOrCv
Srf4idP80dhYN//ub7RyVXQbuPtfU1FG7b+UD85cKzISAhtLQbfJdOHxpCvOm8me
bQiXXPFHE7TjaUFkGY60TX5aq3IwGhZ9D8LWZtOL65uBT044XTOb5FRx7j0IYCCE
JTYLTGRneGBok5P2veL86DLXVJTzIUcc9lqfZcHh6Gri5vmTyhNmqag6l2fPF/h+
p3Rg7xK/2qlNP+mlh39N8gK7LqTCyjGRgwu5aKoHaTfcdAQbFUHsPxRgRj/x/bQz
wepsadFVKRsTmwP/tzTM+ABNjlNUizLn0jB9D/HZv7QCe4m5Mhk/hDwZjtsekazg
YkYuVFmPYVybQ0kqr+7VXRQLcYRebYRSmt4OUAugIm3BEwj3Rp2tYXwd/wy5h96F
sDWWjdtZtITvy3gzoReIS4b1Wf+IwAU1bM2HSyQTz5zZEIeHFAtzc53VGfg8e9o9
fsgR2w9geg7bEeFo/vNln4EJYWNAcRFThwffiAhmIZWjJKJLLQkSuevl9wbwZPZF
8/EDrVgH1HbnRHwrQsyTtSKxncd0cY6VdfLU6Zujvy98LpaTdWGIOA46FcgBvack
gGlmIWb7T1FCLFtiI+ynT4jthulw4p4Fr4hLirSsAYMgZK3/4+9Nr5Y7vfpAtOmt
oRz7LRpv1OQTUs2rqS4KXoCJllz9d/yBkqO2/FQQO8O4yKGJdFXsn+os/9E7MXdM
Q3XYct3VNBQXVo68qLE9qMOIVtPdNOnFkVg2G1Evlt5CiF5YnYFs95309qHMEfOR
J1a3Xeh72BgQ2GoPTZ11Adi38c56GiHEZAmASiUScq4cv4DgojL0GeO9LBNyZL9Z
v69M1gxMnn1/jDknFiTyQIpthubQZmbU6NKgFHgRMejjGlskdbTItUScYPg6jNLs
/Qle1sdeY84jZI/iD5OhYTH3zHbG3L6Px77DCSnCihgM0p6/8vzHa2kjkwWLPFt7
+C9SfeAFVLvDN3/NOQbVF1E4UcbuLKmcIuIztDwMhp9updMQJCOEp8pqybGodTNe
5NDjAFlvkztfF6ghoGMV1ohrHvkDxx8yZ4LaQ1rfsPO1Bdye+7qsbVDyVn1hvI3K
okC56ACOp2n8WVbcfwmlItKMOpaoz2WgX50WyAO9YKoU0XdZNN9LzMLn1145qa4X
bsOYhS7o1YtNSy6Q5K8Qjp2f8xt/bY/ig6JYQnRs48yzSXwN9NxvBb6SNofyo1jH
Tr57Uj4168r7qEpbr4yOGuNakC8EoaDdexqCY+iCZYLPigRJOZ5jfdZspEqhGqa3
dUxdTN738ILmJ+eJFkHoMntd39p2S239Igm5uamJz9k=
`protect END_PROTECTED
