library IEEE;
use IEEE.std_logic_1164.all;

-- The Control Unit
entity ControlUnit is 
	
end;

architecture Behavioural of ControlUnit is
begin
end;