`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mt69IXigaFindss6PFitidwc1WhVEaaEWjkQaH09alXE+FcfQn9/072Ci5A3iDX2
bgE8TakFk6iB18QAZNyHikcjVfaRM1c9u5naObCmNNVPobqqGpnOJ1+SGuV4dMuq
4+hs0zrCke9C4SJJ/OgIfTzaFoFr1vXQX9CGvu8mQQnbRtvNjJ9n0Z4LxMaJ6d9n
wZbYBUBYssEcPb6AGgIdjCePkhDw1g7IATFMNLzaK2aZEfnvzFWG7UaxTj1qMpM5
T9lLLMCRGYEkRi2PXO5/ZOzSyb+D9Bv1cj+hEiUpU+1iEiQUwI49+kOhS4NJKvJn
jnFjhjM8KwVUSFeLmvMppRNVs4LUAnJ7h8Z6c5gQWaZWg1QoSmCHtaTSN7SL+tGG
/AYg7vFhl8XHy+0rTh5WDePMZQPlhb8vdce0B6DUoPtr7xPJjdC7mMgQDmw908Jg
`protect END_PROTECTED
