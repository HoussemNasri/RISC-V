`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/kpEnGsM+lDV4++SJ7DtcXWBYSc1zDkCoD1lBxlAEUINZwtTU/KhCzfBeTJNt/S
ewt/k7UqbRUtZjJjIXzOrsogShcIPIvgGcTcIjsU2plSFDbtCWyeiEoM6J9iABDY
EPLPLlaQaHB71sy7JYpN25IVRlsMDUPcPyHD+odqNtak/ifn17gf5Cgumf+YNR4b
So+ndRPnbEUvzjBRe9Z24W+IwueNKkKXZy0ecuj3/IngbXJcvfLTVAxwhIFWmnzO
7qywa7rt7Zu5WTwUHe1Z6qJ2MS75YUDvEDuze3LeiCnHkDANIq3lzJUb2VZCQBSs
oQz6w8Slblj34vDEI27AICpOm1J5m3WKCOBlnrpmcR+tOiHDmZTCNGUGE7Za7NCI
FlizmrPiI7Qx5wCJ2k1a9tsSWKqtvLqy/TDZ+ncwrIy0idKV98jv21a3W0vrBX6Y
pqVN3EJg+RNWPgO7zgKy0keyIoLK8I++9UY/PRY4PgqJbB8PDMEDGQgNwWnTmOif
AXfMcE4pwEfZvtAeqT2N4M2DoCpjoc84BWF/Tldnbocw1/Ig7WkJA5ufTLnHWaYD
+a2wgCmmbwsHp5fBCQfcorYksQprzpwBu8UD76yRjQGS4KFYVMDDNL9y9kSU7gxq
z9eNVcJuwsaqLqqIc8BNHSF905E5cAFh2G5UeVCbE/+bOdHKQDsxzVxph9Tb2h9B
XnMCZAC9Gf2I5ySmSXyhOfGG8EPLn6GTcV9i8EBzWPNkV4rmpc9M6Kt7IOWuur4Q
ePtOQ+7eduy7qZvmB0pYOTEkyCRVu5LjQUWsp5sjq7ck9N/uTgmYQSK/v/bxrTG4
XN+Bt3+9tB+Roax9AxEAFudyLdw08q13RV6+/P9IZeIJHm0sPvPvRe0yP+NWIWbf
XLDz1Um717PR9g887ZtKrUh6Kgnmo3lvYFil8JEBEFBooDVhP4VrLzIdFYjYvush
/kd5yttkRSoiBSeNItXxNHv6+K841nNxG8G8KL/pXb2w9xNg9tc+ogxGCFDa3i04
PsQxoUQgdI5exdSu3xpgmKyzybdNCRw0eACnpr+i61MIfmmTftwkdkSjsvvBaK++
D8ZtW9y6DkDEwtCbfdEQwrzDfr0+3HapPGViDeM/MATuQE0xr026kZyRMnuxQpr+
K4RLTZDLoYu74+kzKm9t/fwSepFt73SVR6qtuUTAeRyEEPSsKDzUmKxGD29BpgtF
Lt2j0jyn8whOGQOEjbtqNB0edIMH2m/smIgAxGRJt2/ZOu2bM7XxBbNgw+ixvsJQ
hfQzs4tVRgolIw9Jp5nkMFqm+uU6XuHISsteXU6HS05hrPlEl1yFiLc0ln06ejHf
+ZIgIPcWX4W6B2BKwAbYQpf0AFsDVmMT9W/cBs45DWI7PRYaveOUvLpvgA+rMwp5
ezM5n6/OWqE+K3+7iifccNrvJi4UGz63pP1H40Oqew7HX3MIa6q2YqouOFPc77Ww
J72U6lib7gBKfzdzvcLFydUCe10yQBheLu+GeTk8gsGYnlw4ryt6kTUhOfD97SU+
pK+2BVEuwF+8SwyckHbaBcGRoMkmo3j+1JHfh7Rqop7llcQhMar4BaXWbvby/Hno
Iy8ENRlFXlvcw1osbtO+zb3pjz3Y1xPhpD7JXic7AMUIc5ftPqzX9BJt/1eRIyOi
kRVzWYf33B59RM21DI62HYzEg1tCUdqVno7Hw/OimZbZm/fa2vmnPjml4SJTwueV
SVAnA4CfROvNNZbDkO+TGxMshK6VykNrqC30IAHjaJu5BrIvd/YYItj70YF1bY7P
aJiYvrYcsyF7wLaxq/Bl5TylKQJS7SXSD1kUuz6OBjYoSvzJS11Tvg5rlDQ/hjpX
3XIHpGYEeae7/dC6QEMnlNl+W3Z9T2aJuz7lxlc3ym5WaYzWLYLtszeyaTjLapgw
DBSxJmdhWI24v0ox8GySZU7D3ikRr/wntcTb0v7xNsDFhfOnIjlMf4xfQrCtBqtR
mBFB3D3TQZDto50xrVjLg0v0j043LXHhRTpnwfepXKPZ/Mu4rGsWKOjssEFgWd7d
siDZQGKXmSLsAi6dXsVTaF1abTjn1RLQcftjGFv6QdM2WKFlapJXkjRiITB3XCkW
FxRGWND3Q3SNnhKrrit06LT+MHRa9ZtErZfZQxzJCmreyXUWxAvCONxCxOUcBbJ6
0fF6cMT8BhV4h31mxRCrC1JMmacPSyqEXlarbf8uoC/eJDdQhU4MpHcpXiylp6xL
IZ8U6dm+Rx+yyqcAaT2H+ENpmQ7EQEI40HlkUZT3oxTlvISDZKYCwnwKxojuH2aC
luZcNQQPWuKWc8/MzUm3TFR8Mi9zk64eDu1bIESqiImwpjiPFnq/ZOxIavwGNJoz
cdZSeVj+soojYkDs3I/L4yVFN+ei4Iry0Z0AxWdcWKnk3xh1Y4sy1bwYq3Tmbdjc
o+8D9CBlaXvbUlVb6Wtb0lJWfQXbUW/hCJrdhwzfc/Bj2Y9h3PhbaP8x0YGqB16N
S9hY/L9gc1emTHTdXGtlzJO8MH2UCJQ1ZLRfLIRBZs+RdkPr5WH1FWioqrgw4bs5
HY6NUALoAFWm0s5tEBA5CIqxyisf5wwoB3Obo/NVfixGQ1aT4YaYmVwKfGmv5Xqy
JFKFOEyuF9AF3dawtQ71jKY3ArqjFzWv8CKHw+DV/lecg4MEmUy/Ctvg4z32rRtX
lV0UiFTyzmimDUbdNmM6yHpRor5tnwP345LwFiFlFRVwScAyOJ+YdoSrgRjd9AZN
ylvwcxc36TtLs109LQi/ujQNCEwU82vx5+Yh3rvEUgvgc6rAz3OqOLRRTym60jk+
CbmIPzs/WpeNMTfCh0197pbZgCUysEicQguwZCqRZfrXIz2/1eUHMRZAulvUqYM8
Yw7k31mMoowWyT9J/ZyTF1VMH8N67Q5polqT5QM8LeV9PW2+KG7ZxObUjzYxoDxE
TPLsKq5Wko8WQdigB56DpcV8M35cKeQjF6jaUWOff4tnfMFsk/9ECpAtiZ1oM4m/
jvvgJZhg6rGiuhZjjYaE3PYl9K/OwJKNi6bJcV+FQcfy3v4hWiXRVp5xLfQSC5Yf
aBC4MDYhBD4DSHBaVSo2bGcp23nhQozMjTJCDUZiODMOU0Grgq56FV+6dkdkcEno
8DmxRjb+BaEqAo0pfBClXcZBDIX0IdWxgrj1GpNpC3VlmE9CgBCU9XvFkYHJR0U2
ObJka2g6Ju+eOTDtW+mbUNw0BS/b9Gqs0m1S+Ph3M1MwBzrq5EMEJ7Tj+mz81ECj
4J1bi3lRKpBeyLlDEaQQl0JuR7Vn/nbfDjlAeIgWVAMOyZ6ETUJb5RZQC9hbNP1v
ZKJa0C9eQh/5rcBTBYU5ccG7mcl9WLK5RyRFGBEMjObM6zzyjuYhfpaZcZkRl9RD
wtyg3TvRSiJixXqnBDuqbZy+RT69rgUyt/YYEEX/EtN7YgU1rqynMHBVnSOY8nXE
SdUpmlQ1/5gweqxHMOZSQEB+FbjbZ6e2qioYUZw7+UajWfulrWXrXz9siKkKHvba
zCYZrQpfetWZ3kBUw23pwv5IOqiussUYGPH9po/vSr6w3CZ89mGXLIumw0nxE1Rm
rGpEpXCqVzFSEKwMSp5xL/FIlFDVzl8NDfPBp0jPvvVx6zQXfiL7X9QNUcx4/aLt
jZa78B6+87XFKFXjrlRMfpx++Ql7HkWzl5M2lBnIUCJjHfBtrWPT/+0Qh2q+u4yN
ORLgRzV7cXGXfPXOrjsYi1PUjVDJdnYw9JEWZEhqTW8ZYWIcjN+7WflmXroe+Eno
vkYsTSo9XM1rZVATlMoiQHGUGqf5/z8kV0esrcTerfuiIVffJytQEvH5XV6MaoGw
/jblN1DZZTP19YNrB0NqienmKSIK9JJtR/OCkMiDXQQAb3BBnTPDfgxengR6suZu
3SVXz2ad1sGu3Bm5+HcmPY1RWP3TaCgt/fNwC338ucjAWjXR8GNk6cbK/qVMh83X
hPX8R+sPxa8Mq4itqsfMe+DQEjjwKBaerRPjNsoIxeEg70jsfBQuI20bBAYrmzjH
8xs1R/Ucqx4+SjvqjnzNyXvlxzrR0u46e4qK0XnRRLHM6GAM82w+pzG5uLiQD74M
am69diwz/n3rG+uVYZaTaFohFk2Qu0geruE528HL0w2m1dhQs/qP4WaHZwqBLCl/
cAqJ8zRJHoLUlZcr+Gt9qSeP6wh7gMOG0cpVQ9uNdAZ6XVT1QlpijAYhAxB2xUgr
F05WGXq9kz4gsZOgElm4IOAElfoh5WGdP1XesXaHoCTm0cgbZjt2JpQNODrxTTyN
S3eHH0RZaQJN9Qf6/MhYlLgPA245D+s9lR6OWKYKFpIJea0wXQQ1xUsJt9eK4Fna
RuRPWS2HPr+sv2vqEmvYr0k5Ep4gJSFJ/qDXc+MhzDNVAPLTOHB12sz/FT8G+mI3
g0OIk9zix5o/V014tJRt4igm1ohkOAxPs62fc8qRBf9iyJiw1+3GWbjRk+r5zfke
FDdX4uCYR4/P+OMGIVsue3ngnR6+6JZ53fyPlF8Q9tnFp+Y/cKiSppIip9XYpSkM
UImGIwdScTNcqZ9aoMpARAHjxEZ6+zmdKSuR/GaG9v9G4e3EgXC8CRExAlnPMDCY
rO7KXjIYHOfgOlsWAW1pa1N+v/r8CznhgVw++vb0xg4A0ZsWYSIWa7srXvuMO2/6
WKRiFdJuAj8Rc9kqPY5jZlzzlA2W7n0XOIDEMTRCR1rHfGWisUARnELEDW3KiziI
DjVdbLZtk0N+dPJ/xTjIeGzlB+6QAq4+O1fxnqeFf+MYml++kOq3sX7Sal82m4Fi
y1wA8iJLAyp38m0IcKhUi4fL0ZjB0t0ppBdnTUFtPLPxk8myb3J6FzSeg84lnJz0
qT9R1E9qxtxSzRM+08cNQ890ge6Zj7y7jPPqcwLgS7FrrlgNCDjxRUrxzGNZkJjv
GWmrrBEAjb5pHAWaKhynrNwANbda5MyuPSQjPbTg/GutfXlpBLT384gqif4toCId
Fiq5+CF64QnCGfPjF88dzX9aolLsGRPYZE9GSmIRnhMbAgKD+RvcsMiuLLnMlquD
Fslk3x0IJ74OrJSuo0fCkhlaJ+TXPYpUyuEh0cjapIC2DRy1O32E/ArjRDZ6RWQU
fd/9TNhemwZpFlMXenZV+EXrZe0i3XTPRXXD1ZSHmhZRzS+iqLFeUpUVKM5IVBlW
r5lxmJscDWOz1jQs2fgXPAm1afWJINxbYiqEze81ttwo22zG6kKSBT9CfV5B0xQe
Adec+/6WXEMbGQTDljpOoA==
`protect END_PROTECTED
